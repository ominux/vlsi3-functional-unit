
module Alu ( Z, A, B, INST, SEL );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  input SEL;
  wire   N52, N53, N54, N55, N56, N57, N124, N125, N126, N127, N128, N129,
         N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, N140,
         N141, N142, N143, N144, N145, N146, N149, N152, N154, N155, N157,
         N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N181,
         N184, N185, N186, N187, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N373, N376, N378, N379,
         \add_x_10_2/A[31] , \add_x_10_2/A[30] , \add_x_10_2/A[29] ,
         \add_x_10_2/A[25] , \add_x_10_2/A[22] , \add_x_10_2/A[21] ,
         \add_x_10_2/n113 , \add_x_10_2/n111 , \add_x_10_2/n110 ,
         \add_x_10_2/n109 , \add_x_10_2/n107 , \add_x_10_2/n106 ,
         \add_x_10_2/n104 , \add_x_10_2/n102 , \add_x_10_2/n101 ,
         \add_x_10_2/n99 , \add_x_10_2/n97 , \add_x_10_2/n95 ,
         \add_x_10_2/n94 , \add_x_10_2/n93 , \add_x_10_2/n91 ,
         \add_x_10_2/n90 , \add_x_10_2/n88 , \add_x_10_2/n87 ,
         \add_x_10_2/n86 , \add_x_10_2/n85 , \add_x_10_2/n84 ,
         \add_x_10_2/n82 , \add_x_10_2/n81 , \add_x_10_2/n79 ,
         \add_x_10_2/n78 , \add_x_10_2/n76 , \add_x_10_2/n74 ,
         \add_x_10_2/n72 , \add_x_10_2/n70 , \add_x_10_2/n68 ,
         \add_x_10_2/n67 , \add_x_10_2/n66 , \add_x_10_2/n64 ,
         \add_x_10_2/n62 , \add_x_10_2/n60 , \add_x_10_2/n59 ,
         \add_x_10_2/n57 , \add_x_10_2/n55 , \add_x_10_2/n53 ,
         \add_x_10_2/n51 , \add_x_10_2/n50 , \add_x_10_2/n49 ,
         \add_x_10_2/n48 , \add_x_10_2/n47 , \add_x_10_2/n46 ,
         \add_x_10_2/n44 , \add_x_10_2/n42 , \add_x_10_2/n40 ,
         \add_x_10_2/n39 , \add_x_10_2/n38 , \add_x_10_2/n36 ,
         \add_x_10_2/n35 , \add_x_10_2/n33 , \add_x_10_2/n32 ,
         \add_x_10_2/n31 , \add_x_10_2/n29 , \add_x_10_2/n27 ,
         \add_x_10_2/n26 , \add_x_10_2/n23 , \add_x_10_2/n22 ,
         \add_x_10_2/n20 , \add_x_10_2/n19 , \add_x_10_2/n17 ,
         \add_x_10_2/n15 , \add_x_10_2/n14 , \add_x_10_2/n12 ,
         \add_x_10_2/n10 , \add_x_10_2/n9 , \add_x_10_2/n7 , \add_x_10_2/n5 ,
         \add_x_10_2/n4 , \add_x_10_2/n1 , \sub_x_10_3/n225 ,
         \sub_x_10_3/n224 , \sub_x_10_3/n223 , \sub_x_10_3/n222 ,
         \sub_x_10_3/n221 , \sub_x_10_3/n220 , \sub_x_10_3/n219 ,
         \sub_x_10_3/n218 , \sub_x_10_3/n217 , \sub_x_10_3/n216 ,
         \sub_x_10_3/n215 , \sub_x_10_3/n214 , \sub_x_10_3/n213 ,
         \sub_x_10_3/n212 , \sub_x_10_3/n211 , \sub_x_10_3/n210 ,
         \sub_x_10_3/n209 , \sub_x_10_3/n208 , \sub_x_10_3/n207 ,
         \sub_x_10_3/n206 , \sub_x_10_3/n205 , \sub_x_10_3/n201 ,
         \sub_x_10_3/n194 , \sub_x_10_3/n193 , \sub_x_10_3/n192 ,
         \sub_x_10_3/n191 , \sub_x_10_3/n190 , \sub_x_10_3/n189 ,
         \sub_x_10_3/n188 , \sub_x_10_3/n187 , \sub_x_10_3/n186 ,
         \sub_x_10_3/n185 , \sub_x_10_3/n184 , \sub_x_10_3/n183 ,
         \sub_x_10_3/n182 , \sub_x_10_3/n181 , \sub_x_10_3/n180 ,
         \sub_x_10_3/n179 , \sub_x_10_3/n178 , \sub_x_10_3/n176 ,
         \sub_x_10_3/n175 , \sub_x_10_3/n174 , \sub_x_10_3/n173 ,
         \sub_x_10_3/n172 , \sub_x_10_3/n171 , \sub_x_10_3/n170 ,
         \sub_x_10_3/n169 , \sub_x_10_3/n168 , \sub_x_10_3/n167 ,
         \sub_x_10_3/n166 , \sub_x_10_3/n165 , \sub_x_10_3/n164 ,
         \sub_x_10_3/n163 , \sub_x_10_3/n162 , \sub_x_10_3/n161 ,
         \sub_x_10_3/n160 , \sub_x_10_3/n159 , \sub_x_10_3/n158 ,
         \sub_x_10_3/n157 , \sub_x_10_3/n156 , \sub_x_10_3/n155 ,
         \sub_x_10_3/n154 , \sub_x_10_3/n153 , \sub_x_10_3/n150 ,
         \sub_x_10_3/n149 , \sub_x_10_3/n148 , \sub_x_10_3/n147 ,
         \sub_x_10_3/n145 , \sub_x_10_3/n144 , \sub_x_10_3/n143 ,
         \sub_x_10_3/n142 , \sub_x_10_3/n141 , \sub_x_10_3/n140 ,
         \sub_x_10_3/n139 , \sub_x_10_3/n138 , \sub_x_10_3/n137 ,
         \sub_x_10_3/n136 , \sub_x_10_3/n135 , \sub_x_10_3/n134 ,
         \sub_x_10_3/n132 , \sub_x_10_3/n131 , \sub_x_10_3/n130 ,
         \sub_x_10_3/n129 , \sub_x_10_3/n128 , \sub_x_10_3/n125 ,
         \sub_x_10_3/n124 , \sub_x_10_3/n123 , \sub_x_10_3/n122 ,
         \sub_x_10_3/n120 , \sub_x_10_3/n119 , \sub_x_10_3/n118 ,
         \sub_x_10_3/n117 , \sub_x_10_3/n116 , \sub_x_10_3/n115 ,
         \sub_x_10_3/n114 , \sub_x_10_3/n113 , \sub_x_10_3/n112 ,
         \sub_x_10_3/n111 , \sub_x_10_3/n110 , \sub_x_10_3/n109 ,
         \sub_x_10_3/n108 , \sub_x_10_3/n107 , \sub_x_10_3/n105 ,
         \sub_x_10_3/n104 , \sub_x_10_3/n103 , \sub_x_10_3/n102 ,
         \sub_x_10_3/n101 , \sub_x_10_3/n100 , \sub_x_10_3/n99 ,
         \sub_x_10_3/n98 , \sub_x_10_3/n97 , \sub_x_10_3/n96 ,
         \sub_x_10_3/n95 , \sub_x_10_3/n94 , \sub_x_10_3/n93 ,
         \sub_x_10_3/n92 , \sub_x_10_3/n91 , \sub_x_10_3/n88 ,
         \sub_x_10_3/n87 , \sub_x_10_3/n86 , \sub_x_10_3/n85 ,
         \sub_x_10_3/n84 , \sub_x_10_3/n83 , \sub_x_10_3/n82 ,
         \sub_x_10_3/n81 , \sub_x_10_3/n80 , \sub_x_10_3/n79 ,
         \sub_x_10_3/n78 , \sub_x_10_3/n76 , \sub_x_10_3/n74 ,
         \sub_x_10_3/n73 , \sub_x_10_3/n72 , \sub_x_10_3/n71 ,
         \sub_x_10_3/n69 , \sub_x_10_3/n67 , \sub_x_10_3/n65 ,
         \sub_x_10_3/n64 , \sub_x_10_3/n63 , \sub_x_10_3/n62 ,
         \sub_x_10_3/n58 , \sub_x_10_3/n57 , \sub_x_10_3/n56 ,
         \sub_x_10_3/n55 , \sub_x_10_3/n50 , \sub_x_10_3/n49 ,
         \sub_x_10_3/n48 , \sub_x_10_3/n47 , \sub_x_10_3/n42 ,
         \sub_x_10_3/n41 , \sub_x_10_3/n40 , \sub_x_10_3/n39 ,
         \sub_x_10_3/n38 , \sub_x_10_3/n34 , \sub_x_10_3/n33 ,
         \sub_x_10_3/n31 , \sub_x_10_3/n30 , \sub_x_10_3/n29 ,
         \sub_x_10_3/n28 , \sub_x_10_3/n27 , \sub_x_10_3/n26 ,
         \sub_x_10_3/n25 , \sub_x_10_3/n24 , \sub_x_10_3/n23 ,
         \sub_x_10_3/n22 , \sub_x_10_3/n21 , \sub_x_10_3/n20 ,
         \sub_x_10_3/n19 , \sub_x_10_3/n18 , \sub_x_10_3/n17 ,
         \sub_x_10_3/n16 , \sub_x_10_3/n15 , \sub_x_10_3/n14 ,
         \sub_x_10_3/n13 , \sub_x_10_3/n12 , \sub_x_10_3/n11 ,
         \sub_x_10_3/n10 , \sub_x_10_3/n7 , \sub_x_10_3/n4 , \sub_x_10_3/n3 ,
         \sub_x_10_3/n2 , \sub_x_10_3/n1 , \add_x_10_1/n227 ,
         \add_x_10_1/n226 , \add_x_10_1/n225 , \add_x_10_1/n224 ,
         \add_x_10_1/n223 , \add_x_10_1/n222 , \add_x_10_1/n221 ,
         \add_x_10_1/n220 , \add_x_10_1/n219 , \add_x_10_1/n218 ,
         \add_x_10_1/n217 , \add_x_10_1/n216 , \add_x_10_1/n215 ,
         \add_x_10_1/n214 , \add_x_10_1/n213 , \add_x_10_1/n212 ,
         \add_x_10_1/n211 , \add_x_10_1/n210 , \add_x_10_1/n209 ,
         \add_x_10_1/n208 , \add_x_10_1/n207 , \add_x_10_1/n203 ,
         \add_x_10_1/n196 , \add_x_10_1/n194 , \add_x_10_1/n193 ,
         \add_x_10_1/n192 , \add_x_10_1/n191 , \add_x_10_1/n190 ,
         \add_x_10_1/n189 , \add_x_10_1/n188 , \add_x_10_1/n187 ,
         \add_x_10_1/n186 , \add_x_10_1/n185 , \add_x_10_1/n184 ,
         \add_x_10_1/n183 , \add_x_10_1/n182 , \add_x_10_1/n181 ,
         \add_x_10_1/n180 , \add_x_10_1/n179 , \add_x_10_1/n177 ,
         \add_x_10_1/n176 , \add_x_10_1/n175 , \add_x_10_1/n174 ,
         \add_x_10_1/n173 , \add_x_10_1/n172 , \add_x_10_1/n171 ,
         \add_x_10_1/n170 , \add_x_10_1/n169 , \add_x_10_1/n168 ,
         \add_x_10_1/n167 , \add_x_10_1/n166 , \add_x_10_1/n165 ,
         \add_x_10_1/n164 , \add_x_10_1/n163 , \add_x_10_1/n162 ,
         \add_x_10_1/n161 , \add_x_10_1/n160 , \add_x_10_1/n159 ,
         \add_x_10_1/n158 , \add_x_10_1/n157 , \add_x_10_1/n156 ,
         \add_x_10_1/n155 , \add_x_10_1/n154 , \add_x_10_1/n151 ,
         \add_x_10_1/n150 , \add_x_10_1/n149 , \add_x_10_1/n148 ,
         \add_x_10_1/n146 , \add_x_10_1/n145 , \add_x_10_1/n144 ,
         \add_x_10_1/n143 , \add_x_10_1/n142 , \add_x_10_1/n141 ,
         \add_x_10_1/n140 , \add_x_10_1/n139 , \add_x_10_1/n138 ,
         \add_x_10_1/n137 , \add_x_10_1/n136 , \add_x_10_1/n135 ,
         \add_x_10_1/n133 , \add_x_10_1/n132 , \add_x_10_1/n131 ,
         \add_x_10_1/n130 , \add_x_10_1/n129 , \add_x_10_1/n126 ,
         \add_x_10_1/n125 , \add_x_10_1/n124 , \add_x_10_1/n123 ,
         \add_x_10_1/n121 , \add_x_10_1/n120 , \add_x_10_1/n119 ,
         \add_x_10_1/n118 , \add_x_10_1/n117 , \add_x_10_1/n116 ,
         \add_x_10_1/n115 , \add_x_10_1/n114 , \add_x_10_1/n113 ,
         \add_x_10_1/n112 , \add_x_10_1/n111 , \add_x_10_1/n110 ,
         \add_x_10_1/n109 , \add_x_10_1/n108 , \add_x_10_1/n106 ,
         \add_x_10_1/n105 , \add_x_10_1/n104 , \add_x_10_1/n103 ,
         \add_x_10_1/n102 , \add_x_10_1/n101 , \add_x_10_1/n100 ,
         \add_x_10_1/n99 , \add_x_10_1/n98 , \add_x_10_1/n97 ,
         \add_x_10_1/n96 , \add_x_10_1/n95 , \add_x_10_1/n94 ,
         \add_x_10_1/n93 , \add_x_10_1/n92 , \add_x_10_1/n91 ,
         \add_x_10_1/n90 , \add_x_10_1/n89 , \add_x_10_1/n88 ,
         \add_x_10_1/n87 , \add_x_10_1/n86 , \add_x_10_1/n85 ,
         \add_x_10_1/n84 , \add_x_10_1/n83 , \add_x_10_1/n82 ,
         \add_x_10_1/n81 , \add_x_10_1/n80 , \add_x_10_1/n79 ,
         \add_x_10_1/n77 , \add_x_10_1/n75 , \add_x_10_1/n74 ,
         \add_x_10_1/n73 , \add_x_10_1/n72 , \add_x_10_1/n70 ,
         \add_x_10_1/n68 , \add_x_10_1/n66 , \add_x_10_1/n65 ,
         \add_x_10_1/n64 , \add_x_10_1/n63 , \add_x_10_1/n61 ,
         \add_x_10_1/n59 , \add_x_10_1/n58 , \add_x_10_1/n57 ,
         \add_x_10_1/n56 , \add_x_10_1/n55 , \add_x_10_1/n51 ,
         \add_x_10_1/n50 , \add_x_10_1/n49 , \add_x_10_1/n48 ,
         \add_x_10_1/n47 , \add_x_10_1/n45 , \add_x_10_1/n43 ,
         \add_x_10_1/n42 , \add_x_10_1/n41 , \add_x_10_1/n40 ,
         \add_x_10_1/n39 , \add_x_10_1/n37 , \add_x_10_1/n35 ,
         \add_x_10_1/n34 , \add_x_10_1/n31 , \add_x_10_1/n30 ,
         \add_x_10_1/n29 , \add_x_10_1/n28 , \add_x_10_1/n27 ,
         \add_x_10_1/n26 , \add_x_10_1/n25 , \add_x_10_1/n24 ,
         \add_x_10_1/n23 , \add_x_10_1/n22 , \add_x_10_1/n21 ,
         \add_x_10_1/n20 , \add_x_10_1/n19 , \add_x_10_1/n18 ,
         \add_x_10_1/n17 , \add_x_10_1/n16 , \add_x_10_1/n15 ,
         \add_x_10_1/n14 , \add_x_10_1/n13 , \add_x_10_1/n12 ,
         \add_x_10_1/n11 , \add_x_10_1/n10 , \add_x_10_1/n7 , \add_x_10_1/n4 ,
         \add_x_10_1/n3 , \add_x_10_1/n2 , \add_x_10_1/n1 , \cmp6_10_0/n134 ,
         \cmp6_10_0/n133 , \cmp6_10_0/n132 , \cmp6_10_0/n131 ,
         \cmp6_10_0/n130 , \cmp6_10_0/n129 , \cmp6_10_0/n127 ,
         \cmp6_10_0/n126 , \cmp6_10_0/n125 , \cmp6_10_0/n124 ,
         \cmp6_10_0/n123 , \cmp6_10_0/n122 , \cmp6_10_0/n121 ,
         \cmp6_10_0/n118 , \cmp6_10_0/n116 , \cmp6_10_0/n115 ,
         \cmp6_10_0/n114 , \cmp6_10_0/n112 , \cmp6_10_0/n110 ,
         \cmp6_10_0/n109 , \cmp6_10_0/n108 , \cmp6_10_0/n107 ,
         \cmp6_10_0/n106 , \cmp6_10_0/n105 , \cmp6_10_0/n100 , \cmp6_10_0/n99 ,
         \cmp6_10_0/n97 , \cmp6_10_0/n96 , \cmp6_10_0/n95 , \cmp6_10_0/n94 ,
         \cmp6_10_0/n93 , \cmp6_10_0/n92 , \cmp6_10_0/n91 , \cmp6_10_0/n89 ,
         \cmp6_10_0/n88 , \cmp6_10_0/n87 , \cmp6_10_0/n86 , \cmp6_10_0/n85 ,
         \cmp6_10_0/n84 , \cmp6_10_0/n83 , \cmp6_10_0/n82 , \cmp6_10_0/n81 ,
         \cmp6_10_0/n80 , \cmp6_10_0/n79 , \cmp6_10_0/n78 , \cmp6_10_0/n77 ,
         \cmp6_10_0/n76 , \cmp6_10_0/n75 , \cmp6_10_0/n74 , \cmp6_10_0/n73 ,
         \cmp6_10_0/n72 , \cmp6_10_0/n71 , \cmp6_10_0/n69 , \cmp6_10_0/n68 ,
         \cmp6_10_0/n67 , \cmp6_10_0/n65 , \cmp6_10_0/n64 , \cmp6_10_0/n63 ,
         \cmp6_10_0/n62 , \cmp6_10_0/n61 , \cmp6_10_0/n60 , \cmp6_10_0/n59 ,
         \cmp6_10_0/n56 , \cmp6_10_0/n54 , \cmp6_10_0/n53 , \cmp6_10_0/n52 ,
         \cmp6_10_0/n50 , \cmp6_10_0/n48 , \cmp6_10_0/n47 , \cmp6_10_0/n46 ,
         \cmp6_10_0/n45 , \cmp6_10_0/n44 , \cmp6_10_0/n43 , \cmp6_10_0/n40 ,
         \cmp6_10_0/n38 , \cmp6_10_0/n37 , \cmp6_10_0/n36 , \cmp6_10_0/n35 ,
         \cmp6_10_0/n34 , \cmp6_10_0/n33 , \cmp6_10_0/n32 , \cmp6_10_0/n27 ,
         \cmp6_10_0/n26 , \cmp6_10_0/n25 , \cmp6_10_0/n24 , \cmp6_10_0/n23 ,
         \cmp6_10_0/n22 , \cmp6_10_0/n17 , \cmp6_10_0/n16 , \cmp6_10_0/n15 ,
         \cmp6_10_0/n14 , \cmp6_10_0/n13 , \cmp6_10_0/n12 , \cmp6_10_0/n7 ,
         \cmp6_10_0/n6 , \cmp6_10_0/n5 , \cmp6_10_0/n4 , n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615;

  SEN_NR2_1 \add_x_10_2/U124  ( .A1(\add_x_10_2/n101 ), .A2(A[4]), .X(
        \add_x_10_2/n97 ) );
  SEN_NR2_1 \add_x_10_2/U81  ( .A1(\add_x_10_2/n67 ), .A2(A[12]), .X(
        \add_x_10_2/n62 ) );
  SEN_NR2_1 \add_x_10_2/U57  ( .A1(\add_x_10_2/n46 ), .A2(A[16]), .X(
        \add_x_10_2/n42 ) );
  SEN_ND2_G_1 \add_x_10_2/U87  ( .A1(\add_x_10_2/n84 ), .A2(\add_x_10_2/n68 ), 
        .X(\add_x_10_2/n67 ) );
  SEN_NR2_1 \add_x_10_2/U32  ( .A1(\add_x_10_2/n46 ), .A2(\add_x_10_2/n23 ), 
        .X(\add_x_10_2/n22 ) );
  SEN_ND2_G_1 \add_x_10_2/U7  ( .A1(\add_x_10_2/n7 ), .A2(\add_x_10_2/n5 ), 
        .X(\add_x_10_2/n4 ) );
  SEN_ND2_G_1 \add_x_10_2/U14  ( .A1(\add_x_10_2/n12 ), .A2(\add_x_10_2/n10 ), 
        .X(\add_x_10_2/n9 ) );
  SEN_ND2_G_1 \add_x_10_2/U21  ( .A1(\add_x_10_2/n17 ), .A2(\add_x_10_2/n15 ), 
        .X(\add_x_10_2/n14 ) );
  SEN_ND2_G_1 \add_x_10_2/U53  ( .A1(\add_x_10_2/n44 ), .A2(\add_x_10_2/n40 ), 
        .X(\add_x_10_2/n39 ) );
  SEN_ND2_G_1 \add_x_10_2/U109  ( .A1(\add_x_10_2/n86 ), .A2(\add_x_10_2/n102 ), .X(\add_x_10_2/n85 ) );
  SEN_ND2_G_1 \add_x_10_2/U140  ( .A1(\add_x_10_2/n111 ), .A2(
        \add_x_10_2/n113 ), .X(\add_x_10_2/n110 ) );
  SEN_ND2_G_1 \add_x_10_2/U111  ( .A1(\add_x_10_2/n91 ), .A2(\add_x_10_2/n88 ), 
        .X(\add_x_10_2/n87 ) );
  SEN_ND2_G_1 \add_x_10_2/U120  ( .A1(\add_x_10_2/n99 ), .A2(\add_x_10_2/n95 ), 
        .X(\add_x_10_2/n94 ) );
  SEN_ND2_G_1 \add_x_10_2/U64  ( .A1(\add_x_10_2/n68 ), .A2(\add_x_10_2/n49 ), 
        .X(\add_x_10_2/n48 ) );
  SEN_ND2_G_1 \add_x_10_2/U77  ( .A1(\add_x_10_2/n64 ), .A2(\add_x_10_2/n60 ), 
        .X(\add_x_10_2/n59 ) );
  SEN_ND2_G_1 \add_x_10_2/U100  ( .A1(\add_x_10_2/n82 ), .A2(\add_x_10_2/n79 ), 
        .X(\add_x_10_2/n78 ) );
  SEN_EN2_0P5 \add_x_10_2/U138  ( .A1(\add_x_10_2/n113 ), .A2(A[1]), .X(N157)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U128  ( .A1(A[3]), .A2(\add_x_10_2/n106 ), .X(N159) );
  SEN_EN2_0P5 \add_x_10_2/U118  ( .A1(A[5]), .A2(\add_x_10_2/n97 ), .X(N161)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U123  ( .A1(A[4]), .A2(\add_x_10_2/n101 ), .X(N160) );
  SEN_EN2_0P5 \add_x_10_2/U134  ( .A1(A[2]), .A2(\add_x_10_2/n109 ), .X(N158)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U97  ( .A1(A[9]), .A2(\add_x_10_2/n81 ), .X(N165)
         );
  SEN_EN2_0P5 \add_x_10_2/U114  ( .A1(A[6]), .A2(\add_x_10_2/n93 ), .X(N162)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U107  ( .A1(A[7]), .A2(\add_x_10_2/n90 ), .X(N163)
         );
  SEN_EN2_0P5 \add_x_10_2/U103  ( .A1(A[8]), .A2(\add_x_10_2/n84 ), .X(N164)
         );
  SEN_EN2_0P5 \add_x_10_2/U74  ( .A1(A[13]), .A2(\add_x_10_2/n62 ), .X(N169)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U92  ( .A1(A[10]), .A2(\add_x_10_2/n76 ), .X(N166)
         );
  SEN_EN2_0P5 \add_x_10_2/U85  ( .A1(A[11]), .A2(\add_x_10_2/n72 ), .X(N167)
         );
  SEN_EN2_0P5 \add_x_10_2/U80  ( .A1(A[12]), .A2(\add_x_10_2/n66 ), .X(N168)
         );
  SEN_EN2_0P5 \add_x_10_2/U6  ( .A1(A[28]), .A2(\add_x_10_2/n7 ), .X(N184) );
  SEN_EO2_S_0P5 \add_x_10_2/U69  ( .A1(A[14]), .A2(\add_x_10_2/n57 ), .X(N170)
         );
  SEN_EN2_0P5 \add_x_10_2/U51  ( .A1(A[17]), .A2(\add_x_10_2/n42 ), .X(N173)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U56  ( .A1(A[16]), .A2(\add_x_10_2/n46 ), .X(N172)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U17  ( .A1(A[25]), .A2(\add_x_10_2/n14 ), .X(N181)
         );
  SEN_EN2_0P5 \add_x_10_2/U47  ( .A1(A[18]), .A2(\add_x_10_2/n38 ), .X(N174)
         );
  SEN_EN2_0P5 \add_x_10_2/U61  ( .A1(A[15]), .A2(\add_x_10_2/n53 ), .X(N171)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U31  ( .A1(A[21]), .A2(\add_x_10_2/n26 ), .X(N177)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U40  ( .A1(A[19]), .A2(\add_x_10_2/n35 ), .X(N175)
         );
  SEN_EO2_S_0P5 \add_x_10_2/U3  ( .A1(A[29]), .A2(\add_x_10_2/n4 ), .X(N185)
         );
  SEN_EN2_0P5 \add_x_10_2/U36  ( .A1(A[20]), .A2(\add_x_10_2/n29 ), .X(N176)
         );
  SEN_EN2_0P5 \add_x_10_2/U27  ( .A1(A[22]), .A2(\add_x_10_2/n22 ), .X(N178)
         );
  SEN_AOI21_S_1 \sub_x_10_3/U236  ( .A1(\sub_x_10_3/n183 ), .A2(
        \sub_x_10_3/n191 ), .B(\sub_x_10_3/n184 ), .X(\sub_x_10_3/n182 ) );
  SEN_ND2_G_1 \sub_x_10_3/U252  ( .A1(\sub_x_10_3/n225 ), .A2(
        \sub_x_10_3/n193 ), .X(\sub_x_10_3/n31 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U244  ( .A1(\sub_x_10_3/n190 ), .A2(
        \sub_x_10_3/n188 ), .B(\sub_x_10_3/n189 ), .X(\sub_x_10_3/n187 ) );
  SEN_ND2_G_1 \sub_x_10_3/U239  ( .A1(\sub_x_10_3/n223 ), .A2(
        \sub_x_10_3/n186 ), .X(\sub_x_10_3/n29 ) );
  SEN_ND2_G_1 \sub_x_10_3/U222  ( .A1(\sub_x_10_3/n221 ), .A2(
        \sub_x_10_3/n175 ), .X(\sub_x_10_3/n27 ) );
  SEN_ND2_G_1 \sub_x_10_3/U230  ( .A1(\sub_x_10_3/n222 ), .A2(
        \sub_x_10_3/n180 ), .X(\sub_x_10_3/n28 ) );
  SEN_ND2_G_1 \sub_x_10_3/U245  ( .A1(\sub_x_10_3/n224 ), .A2(
        \sub_x_10_3/n189 ), .X(\sub_x_10_3/n30 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U196  ( .A1(\sub_x_10_3/n160 ), .A2(
        \sub_x_10_3/n158 ), .B(\sub_x_10_3/n159 ), .X(\sub_x_10_3/n157 ) );
  SEN_ND2_G_1 \sub_x_10_3/U191  ( .A1(\sub_x_10_3/n217 ), .A2(
        \sub_x_10_3/n156 ), .X(\sub_x_10_3/n23 ) );
  SEN_ND2_G_1 \sub_x_10_3/U214  ( .A1(\sub_x_10_3/n220 ), .A2(
        \sub_x_10_3/n170 ), .X(\sub_x_10_3/n26 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U213  ( .A1(\sub_x_10_3/n171 ), .A2(
        \sub_x_10_3/n169 ), .B(\sub_x_10_3/n170 ), .X(\sub_x_10_3/n168 ) );
  SEN_ND2_G_1 \sub_x_10_3/U208  ( .A1(\sub_x_10_3/n219 ), .A2(
        \sub_x_10_3/n167 ), .X(\sub_x_10_3/n25 ) );
  SEN_ND2_G_1 \sub_x_10_3/U197  ( .A1(\sub_x_10_3/n218 ), .A2(
        \sub_x_10_3/n159 ), .X(\sub_x_10_3/n24 ) );
  SEN_ND2_G_1 \sub_x_10_3/U154  ( .A1(\sub_x_10_3/n213 ), .A2(
        \sub_x_10_3/n131 ), .X(\sub_x_10_3/n19 ) );
  SEN_ND2_G_1 \sub_x_10_3/U181  ( .A1(\sub_x_10_3/n216 ), .A2(
        \sub_x_10_3/n149 ), .X(\sub_x_10_3/n22 ) );
  SEN_ND2_G_1 \sub_x_10_3/U173  ( .A1(\sub_x_10_3/n215 ), .A2(
        \sub_x_10_3/n144 ), .X(\sub_x_10_3/n21 ) );
  SEN_ND2_G_1 \sub_x_10_3/U162  ( .A1(\sub_x_10_3/n214 ), .A2(
        \sub_x_10_3/n136 ), .X(\sub_x_10_3/n20 ) );
  SEN_ND2_G_1 \sub_x_10_3/U144  ( .A1(\sub_x_10_3/n212 ), .A2(
        \sub_x_10_3/n124 ), .X(\sub_x_10_3/n18 ) );
  SEN_ND2_G_1 \sub_x_10_3/U115  ( .A1(\sub_x_10_3/n209 ), .A2(
        \sub_x_10_3/n104 ), .X(\sub_x_10_3/n15 ) );
  SEN_ND2_G_1 \sub_x_10_3/U123  ( .A1(\sub_x_10_3/n210 ), .A2(
        \sub_x_10_3/n109 ), .X(\sub_x_10_3/n16 ) );
  SEN_ND2_G_1 \sub_x_10_3/U107  ( .A1(\sub_x_10_3/n208 ), .A2(\sub_x_10_3/n99 ), .X(\sub_x_10_3/n14 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U168  ( .A1(\sub_x_10_3/n160 ), .A2(
        \sub_x_10_3/n139 ), .B(\sub_x_10_3/n140 ), .X(\sub_x_10_3/n138 ) );
  SEN_ND2_G_1 \sub_x_10_3/U136  ( .A1(\sub_x_10_3/n211 ), .A2(
        \sub_x_10_3/n119 ), .X(\sub_x_10_3/n17 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U87  ( .A1(\sub_x_10_3/n88 ), .A2(\sub_x_10_3/n85 ), .B(\sub_x_10_3/n86 ), .X(\sub_x_10_3/n84 ) );
  SEN_ND2_G_1 \sub_x_10_3/U82  ( .A1(\sub_x_10_3/n205 ), .A2(\sub_x_10_3/n83 ), 
        .X(\sub_x_10_3/n11 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U106  ( .A1(\sub_x_10_3/n100 ), .A2(
        \sub_x_10_3/n98 ), .B(\sub_x_10_3/n99 ), .X(\sub_x_10_3/n97 ) );
  SEN_ND2_G_1 \sub_x_10_3/U101  ( .A1(\sub_x_10_3/n207 ), .A2(\sub_x_10_3/n96 ), .X(\sub_x_10_3/n13 ) );
  SEN_ND2_G_1 \sub_x_10_3/U88  ( .A1(\sub_x_10_3/n206 ), .A2(\sub_x_10_3/n86 ), 
        .X(\sub_x_10_3/n12 ) );
  SEN_ND2_G_1 \sub_x_10_3/U10  ( .A1(n356), .A2(\sub_x_10_3/n38 ), .X(
        \sub_x_10_3/n2 ) );
  SEN_ND2_G_1 \sub_x_10_3/U74  ( .A1(n361), .A2(\sub_x_10_3/n78 ), .X(
        \sub_x_10_3/n10 ) );
  SEN_ND2_G_1 \sub_x_10_3/U13  ( .A1(n335), .A2(A[30]), .X(\sub_x_10_3/n38 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U19  ( .A1(n327), .A2(A[29]), .X(\sub_x_10_3/n41 )
         );
  SEN_NR2_1 \sub_x_10_3/U18  ( .A1(n327), .A2(A[29]), .X(\sub_x_10_3/n40 ) );
  SEN_ND2_G_1 \sub_x_10_3/U33  ( .A1(n332), .A2(A[27]), .X(\sub_x_10_3/n49 )
         );
  SEN_NR2_1 \sub_x_10_3/U32  ( .A1(n332), .A2(A[27]), .X(\sub_x_10_3/n48 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U43  ( .A1(\sub_x_10_3/n58 ), .A2(\sub_x_10_3/n56 ), .B(\sub_x_10_3/n57 ), .X(\sub_x_10_3/n55 ) );
  SEN_ND2_G_1 \sub_x_10_3/U47  ( .A1(n330), .A2(A[25]), .X(\sub_x_10_3/n57 )
         );
  SEN_NR2_1 \sub_x_10_3/U46  ( .A1(n330), .A2(A[25]), .X(\sub_x_10_3/n56 ) );
  SEN_ND2_G_1 \sub_x_10_3/U55  ( .A1(n336), .A2(A[24]), .X(\sub_x_10_3/n62 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U65  ( .A1(n319), .A2(A[23]), .X(\sub_x_10_3/n69 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U69  ( .A1(\sub_x_10_3/n92 ), .A2(\sub_x_10_3/n73 ), .B(\sub_x_10_3/n74 ), .X(\sub_x_10_3/n72 ) );
  SEN_ND2_G_1 \sub_x_10_3/U77  ( .A1(n320), .A2(A[22]), .X(\sub_x_10_3/n78 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U81  ( .A1(\sub_x_10_3/n82 ), .A2(\sub_x_10_3/n86 ), .B(\sub_x_10_3/n83 ), .X(\sub_x_10_3/n81 ) );
  SEN_ND2_G_1 \sub_x_10_3/U85  ( .A1(n317), .A2(A[21]), .X(\sub_x_10_3/n83 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U91  ( .A1(n314), .A2(A[20]), .X(\sub_x_10_3/n86 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U100  ( .A1(\sub_x_10_3/n95 ), .A2(
        \sub_x_10_3/n99 ), .B(\sub_x_10_3/n96 ), .X(\sub_x_10_3/n94 ) );
  SEN_ND2_G_1 \sub_x_10_3/U104  ( .A1(n311), .A2(A[19]), .X(\sub_x_10_3/n96 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U110  ( .A1(n310), .A2(A[18]), .X(\sub_x_10_3/n99 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U118  ( .A1(n315), .A2(A[17]), .X(\sub_x_10_3/n104 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U126  ( .A1(n325), .A2(A[16]), .X(\sub_x_10_3/n109 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U58  ( .A1(\sub_x_10_3/n71 ), .A2(n360), .X(
        \sub_x_10_3/n64 ) );
  SEN_ND2_G_1 \sub_x_10_3/U70  ( .A1(\sub_x_10_3/n80 ), .A2(n361), .X(
        \sub_x_10_3/n73 ) );
  SEN_ND2_G_1 \sub_x_10_3/U97  ( .A1(\sub_x_10_3/n101 ), .A2(\sub_x_10_3/n93 ), 
        .X(\sub_x_10_3/n91 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U131  ( .A1(\sub_x_10_3/n140 ), .A2(
        \sub_x_10_3/n114 ), .B(\sub_x_10_3/n115 ), .X(\sub_x_10_3/n113 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U135  ( .A1(\sub_x_10_3/n118 ), .A2(
        \sub_x_10_3/n124 ), .B(\sub_x_10_3/n119 ), .X(\sub_x_10_3/n117 ) );
  SEN_ND2_G_1 \sub_x_10_3/U139  ( .A1(n309), .A2(A[15]), .X(\sub_x_10_3/n119 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U147  ( .A1(n308), .A2(A[14]), .X(\sub_x_10_3/n124 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U153  ( .A1(\sub_x_10_3/n130 ), .A2(
        \sub_x_10_3/n136 ), .B(\sub_x_10_3/n131 ), .X(\sub_x_10_3/n129 ) );
  SEN_ND2_G_1 \sub_x_10_3/U157  ( .A1(n318), .A2(A[13]), .X(\sub_x_10_3/n131 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U165  ( .A1(n313), .A2(A[12]), .X(\sub_x_10_3/n136 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U172  ( .A1(\sub_x_10_3/n143 ), .A2(
        \sub_x_10_3/n149 ), .B(\sub_x_10_3/n144 ), .X(\sub_x_10_3/n142 ) );
  SEN_ND2_G_1 \sub_x_10_3/U176  ( .A1(n316), .A2(A[11]), .X(\sub_x_10_3/n144 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U184  ( .A1(n326), .A2(A[10]), .X(\sub_x_10_3/n149 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U190  ( .A1(\sub_x_10_3/n155 ), .A2(
        \sub_x_10_3/n159 ), .B(\sub_x_10_3/n156 ), .X(\sub_x_10_3/n154 ) );
  SEN_ND2_G_1 \sub_x_10_3/U194  ( .A1(n312), .A2(A[9]), .X(\sub_x_10_3/n156 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U200  ( .A1(n329), .A2(A[8]), .X(\sub_x_10_3/n159 )
         );
  SEN_NR2_1 \sub_x_10_3/U130  ( .A1(\sub_x_10_3/n139 ), .A2(\sub_x_10_3/n114 ), 
        .X(\sub_x_10_3/n112 ) );
  SEN_ND2_G_1 \sub_x_10_3/U132  ( .A1(\sub_x_10_3/n128 ), .A2(
        \sub_x_10_3/n116 ), .X(\sub_x_10_3/n114 ) );
  SEN_ND2_G_1 \sub_x_10_3/U169  ( .A1(\sub_x_10_3/n153 ), .A2(
        \sub_x_10_3/n141 ), .X(\sub_x_10_3/n139 ) );
  SEN_NR2_1 \sub_x_10_3/U183  ( .A1(n326), .A2(A[10]), .X(\sub_x_10_3/n148 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U203  ( .A1(\sub_x_10_3/n182 ), .A2(
        \sub_x_10_3/n162 ), .B(\sub_x_10_3/n163 ), .X(\sub_x_10_3/n161 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U207  ( .A1(\sub_x_10_3/n166 ), .A2(
        \sub_x_10_3/n170 ), .B(\sub_x_10_3/n167 ), .X(\sub_x_10_3/n165 ) );
  SEN_ND2_G_1 \sub_x_10_3/U211  ( .A1(n324), .A2(A[7]), .X(\sub_x_10_3/n167 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U217  ( .A1(n323), .A2(A[6]), .X(\sub_x_10_3/n170 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U221  ( .A1(\sub_x_10_3/n174 ), .A2(
        \sub_x_10_3/n180 ), .B(\sub_x_10_3/n175 ), .X(\sub_x_10_3/n173 ) );
  SEN_ND2_G_1 \sub_x_10_3/U225  ( .A1(n322), .A2(A[5]), .X(\sub_x_10_3/n175 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U233  ( .A1(n328), .A2(A[4]), .X(\sub_x_10_3/n180 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U204  ( .A1(\sub_x_10_3/n172 ), .A2(
        \sub_x_10_3/n164 ), .X(\sub_x_10_3/n162 ) );
  SEN_NR2_1 \sub_x_10_3/U232  ( .A1(n328), .A2(A[4]), .X(\sub_x_10_3/n179 ) );
  SEN_OAI21_G_1 \sub_x_10_3/U238  ( .A1(\sub_x_10_3/n185 ), .A2(
        \sub_x_10_3/n189 ), .B(\sub_x_10_3/n186 ), .X(\sub_x_10_3/n184 ) );
  SEN_ND2_G_1 \sub_x_10_3/U242  ( .A1(n321), .A2(A[3]), .X(\sub_x_10_3/n186 )
         );
  SEN_ND2_G_1 \sub_x_10_3/U248  ( .A1(n337), .A2(A[2]), .X(\sub_x_10_3/n189 )
         );
  SEN_OAI21_G_1 \sub_x_10_3/U251  ( .A1(\sub_x_10_3/n192 ), .A2(
        \sub_x_10_3/n194 ), .B(\sub_x_10_3/n193 ), .X(\sub_x_10_3/n191 ) );
  SEN_ND2_G_1 \sub_x_10_3/U255  ( .A1(n307), .A2(A[1]), .X(\sub_x_10_3/n193 )
         );
  SEN_NR2_1 \sub_x_10_3/U254  ( .A1(n307), .A2(A[1]), .X(\sub_x_10_3/n192 ) );
  SEN_NR2_1 \sub_x_10_3/U237  ( .A1(\sub_x_10_3/n188 ), .A2(\sub_x_10_3/n185 ), 
        .X(\sub_x_10_3/n183 ) );
  SEN_NR2_1 \sub_x_10_3/U247  ( .A1(n337), .A2(A[2]), .X(\sub_x_10_3/n188 ) );
  SEN_ND2_G_1 \sub_x_10_3/U2  ( .A1(n355), .A2(\sub_x_10_3/n33 ), .X(
        \sub_x_10_3/n1 ) );
  SEN_EO2_S_0P5 \sub_x_10_3/U249  ( .A1(\sub_x_10_3/n194 ), .A2(
        \sub_x_10_3/n31 ), .X(N349) );
  SEN_EN2_0P5 \sub_x_10_3/U234  ( .A1(\sub_x_10_3/n29 ), .A2(\sub_x_10_3/n187 ), .X(N351) );
  SEN_EO2_S_0P5 \sub_x_10_3/U218  ( .A1(\sub_x_10_3/n27 ), .A2(
        \sub_x_10_3/n176 ), .X(N353) );
  SEN_EN2_0P5 \sub_x_10_3/U226  ( .A1(\sub_x_10_3/n28 ), .A2(\sub_x_10_3/n181 ), .X(N352) );
  SEN_EO2_S_0P5 \sub_x_10_3/U243  ( .A1(\sub_x_10_3/n30 ), .A2(
        \sub_x_10_3/n190 ), .X(N350) );
  SEN_EN2_0P5 \sub_x_10_3/U185  ( .A1(\sub_x_10_3/n23 ), .A2(\sub_x_10_3/n157 ), .X(N357) );
  SEN_EO2_S_0P5 \sub_x_10_3/U212  ( .A1(\sub_x_10_3/n26 ), .A2(
        \sub_x_10_3/n171 ), .X(N354) );
  SEN_EN2_0P5 \sub_x_10_3/U201  ( .A1(\sub_x_10_3/n25 ), .A2(\sub_x_10_3/n168 ), .X(N355) );
  SEN_EO2_S_0P5 \sub_x_10_3/U195  ( .A1(\sub_x_10_3/n24 ), .A2(
        \sub_x_10_3/n160 ), .X(N356) );
  SEN_EO2_S_0P5 \sub_x_10_3/U148  ( .A1(\sub_x_10_3/n19 ), .A2(
        \sub_x_10_3/n132 ), .X(N361) );
  SEN_EN2_0P5 \sub_x_10_3/U177  ( .A1(\sub_x_10_3/n22 ), .A2(\sub_x_10_3/n150 ), .X(N358) );
  SEN_EO2_S_0P5 \sub_x_10_3/U166  ( .A1(\sub_x_10_3/n21 ), .A2(
        \sub_x_10_3/n145 ), .X(N359) );
  SEN_EO2_S_0P5 \sub_x_10_3/U158  ( .A1(\sub_x_10_3/n20 ), .A2(
        \sub_x_10_3/n137 ), .X(N360) );
  SEN_EN2_0P5 \sub_x_10_3/U20  ( .A1(\sub_x_10_3/n4 ), .A2(\sub_x_10_3/n47 ), 
        .X(N376) );
  SEN_EN2_0P5 \sub_x_10_3/U140  ( .A1(\sub_x_10_3/n18 ), .A2(\sub_x_10_3/n125 ), .X(N362) );
  SEN_EO2_S_0P5 \sub_x_10_3/U111  ( .A1(\sub_x_10_3/n15 ), .A2(
        \sub_x_10_3/n105 ), .X(N365) );
  SEN_EN2_0P5 \sub_x_10_3/U119  ( .A1(\sub_x_10_3/n16 ), .A2(\sub_x_10_3/n110 ), .X(N364) );
  SEN_EO2_S_0P5 \sub_x_10_3/U42  ( .A1(\sub_x_10_3/n7 ), .A2(\sub_x_10_3/n58 ), 
        .X(N373) );
  SEN_EO2_S_0P5 \sub_x_10_3/U105  ( .A1(\sub_x_10_3/n14 ), .A2(
        \sub_x_10_3/n100 ), .X(N366) );
  SEN_EO2_S_0P5 \sub_x_10_3/U127  ( .A1(\sub_x_10_3/n17 ), .A2(
        \sub_x_10_3/n120 ), .X(N363) );
  SEN_EN2_0P5 \sub_x_10_3/U78  ( .A1(\sub_x_10_3/n11 ), .A2(\sub_x_10_3/n84 ), 
        .X(N369) );
  SEN_EN2_0P5 \sub_x_10_3/U92  ( .A1(\sub_x_10_3/n13 ), .A2(\sub_x_10_3/n97 ), 
        .X(N367) );
  SEN_EN2_0P5 \sub_x_10_3/U86  ( .A1(\sub_x_10_3/n12 ), .A2(\sub_x_10_3/n87 ), 
        .X(N368) );
  SEN_EN2_0P5 \sub_x_10_3/U6  ( .A1(\sub_x_10_3/n2 ), .A2(\sub_x_10_3/n39 ), 
        .X(N378) );
  SEN_EO2_S_0P5 \sub_x_10_3/U66  ( .A1(\sub_x_10_3/n10 ), .A2(\sub_x_10_3/n79 ), .X(N370) );
  SEN_AOI21_S_1 \sub_x_10_3/U133  ( .A1(\sub_x_10_3/n116 ), .A2(
        \sub_x_10_3/n129 ), .B(\sub_x_10_3/n117 ), .X(\sub_x_10_3/n115 ) );
  SEN_AOI21_S_1 \sub_x_10_3/U170  ( .A1(\sub_x_10_3/n141 ), .A2(
        \sub_x_10_3/n154 ), .B(\sub_x_10_3/n142 ), .X(\sub_x_10_3/n140 ) );
  SEN_AOI21_S_1 \sub_x_10_3/U205  ( .A1(\sub_x_10_3/n164 ), .A2(
        \sub_x_10_3/n173 ), .B(\sub_x_10_3/n165 ), .X(\sub_x_10_3/n163 ) );
  SEN_EN2_0P5 \sub_x_10_3/U256  ( .A1(n339), .A2(A[0]), .X(N348) );
  SEN_ND2_G_1 \add_x_10_1/U252  ( .A1(\add_x_10_1/n227 ), .A2(
        \add_x_10_1/n194 ), .X(\add_x_10_1/n31 ) );
  SEN_OAI21_G_1 \add_x_10_1/U244  ( .A1(\add_x_10_1/n191 ), .A2(
        \add_x_10_1/n189 ), .B(\add_x_10_1/n190 ), .X(\add_x_10_1/n188 ) );
  SEN_ND2_G_1 \add_x_10_1/U239  ( .A1(\add_x_10_1/n225 ), .A2(
        \add_x_10_1/n187 ), .X(\add_x_10_1/n29 ) );
  SEN_ND2_G_1 \add_x_10_1/U222  ( .A1(\add_x_10_1/n223 ), .A2(
        \add_x_10_1/n176 ), .X(\add_x_10_1/n27 ) );
  SEN_ND2_G_1 \add_x_10_1/U230  ( .A1(\add_x_10_1/n224 ), .A2(
        \add_x_10_1/n181 ), .X(\add_x_10_1/n28 ) );
  SEN_ND2_G_1 \add_x_10_1/U245  ( .A1(\add_x_10_1/n226 ), .A2(
        \add_x_10_1/n190 ), .X(\add_x_10_1/n30 ) );
  SEN_OAI21_G_1 \add_x_10_1/U196  ( .A1(\add_x_10_1/n161 ), .A2(
        \add_x_10_1/n159 ), .B(\add_x_10_1/n160 ), .X(\add_x_10_1/n158 ) );
  SEN_ND2_G_1 \add_x_10_1/U191  ( .A1(\add_x_10_1/n219 ), .A2(
        \add_x_10_1/n157 ), .X(\add_x_10_1/n23 ) );
  SEN_ND2_G_1 \add_x_10_1/U214  ( .A1(\add_x_10_1/n222 ), .A2(
        \add_x_10_1/n171 ), .X(\add_x_10_1/n26 ) );
  SEN_OAI21_G_1 \add_x_10_1/U213  ( .A1(\add_x_10_1/n172 ), .A2(
        \add_x_10_1/n170 ), .B(\add_x_10_1/n171 ), .X(\add_x_10_1/n169 ) );
  SEN_ND2_G_1 \add_x_10_1/U208  ( .A1(\add_x_10_1/n221 ), .A2(
        \add_x_10_1/n168 ), .X(\add_x_10_1/n25 ) );
  SEN_ND2_G_1 \add_x_10_1/U197  ( .A1(\add_x_10_1/n220 ), .A2(
        \add_x_10_1/n160 ), .X(\add_x_10_1/n24 ) );
  SEN_ND2_G_1 \add_x_10_1/U154  ( .A1(\add_x_10_1/n215 ), .A2(
        \add_x_10_1/n132 ), .X(\add_x_10_1/n19 ) );
  SEN_ND2_G_1 \add_x_10_1/U181  ( .A1(\add_x_10_1/n218 ), .A2(
        \add_x_10_1/n150 ), .X(\add_x_10_1/n22 ) );
  SEN_ND2_G_1 \add_x_10_1/U173  ( .A1(\add_x_10_1/n217 ), .A2(
        \add_x_10_1/n145 ), .X(\add_x_10_1/n21 ) );
  SEN_ND2_G_1 \add_x_10_1/U162  ( .A1(\add_x_10_1/n216 ), .A2(
        \add_x_10_1/n137 ), .X(\add_x_10_1/n20 ) );
  SEN_ND2_G_1 \add_x_10_1/U144  ( .A1(\add_x_10_1/n214 ), .A2(
        \add_x_10_1/n125 ), .X(\add_x_10_1/n18 ) );
  SEN_ND2_G_1 \add_x_10_1/U115  ( .A1(\add_x_10_1/n211 ), .A2(
        \add_x_10_1/n105 ), .X(\add_x_10_1/n15 ) );
  SEN_ND2_G_1 \add_x_10_1/U123  ( .A1(\add_x_10_1/n212 ), .A2(
        \add_x_10_1/n110 ), .X(\add_x_10_1/n16 ) );
  SEN_ND2_G_1 \add_x_10_1/U107  ( .A1(\add_x_10_1/n210 ), .A2(
        \add_x_10_1/n100 ), .X(\add_x_10_1/n14 ) );
  SEN_OAI21_G_1 \add_x_10_1/U168  ( .A1(\add_x_10_1/n161 ), .A2(
        \add_x_10_1/n140 ), .B(\add_x_10_1/n141 ), .X(\add_x_10_1/n139 ) );
  SEN_ND2_G_1 \add_x_10_1/U136  ( .A1(\add_x_10_1/n213 ), .A2(
        \add_x_10_1/n120 ), .X(\add_x_10_1/n17 ) );
  SEN_OAI21_G_1 \add_x_10_1/U87  ( .A1(\add_x_10_1/n89 ), .A2(\add_x_10_1/n86 ), .B(\add_x_10_1/n87 ), .X(\add_x_10_1/n85 ) );
  SEN_ND2_G_1 \add_x_10_1/U82  ( .A1(\add_x_10_1/n207 ), .A2(\add_x_10_1/n84 ), 
        .X(\add_x_10_1/n11 ) );
  SEN_OAI21_G_1 \add_x_10_1/U106  ( .A1(\add_x_10_1/n101 ), .A2(
        \add_x_10_1/n99 ), .B(\add_x_10_1/n100 ), .X(\add_x_10_1/n98 ) );
  SEN_ND2_G_1 \add_x_10_1/U101  ( .A1(\add_x_10_1/n209 ), .A2(\add_x_10_1/n97 ), .X(\add_x_10_1/n13 ) );
  SEN_ND2_G_1 \add_x_10_1/U88  ( .A1(\add_x_10_1/n208 ), .A2(\add_x_10_1/n87 ), 
        .X(\add_x_10_1/n12 ) );
  SEN_ND2_G_1 \add_x_10_1/U10  ( .A1(n349), .A2(\add_x_10_1/n39 ), .X(
        \add_x_10_1/n2 ) );
  SEN_ND2_G_1 \add_x_10_1/U74  ( .A1(n354), .A2(\add_x_10_1/n79 ), .X(
        \add_x_10_1/n10 ) );
  SEN_ND2_G_1 \add_x_10_1/U13  ( .A1(A[30]), .A2(B[30]), .X(\add_x_10_1/n39 )
         );
  SEN_ND2_G_1 \add_x_10_1/U19  ( .A1(A[29]), .A2(B[29]), .X(\add_x_10_1/n42 )
         );
  SEN_NR2_1 \add_x_10_1/U18  ( .A1(A[29]), .A2(B[29]), .X(\add_x_10_1/n41 ) );
  SEN_ND2_G_1 \add_x_10_1/U27  ( .A1(A[28]), .A2(B[28]), .X(\add_x_10_1/n47 )
         );
  SEN_OAI21_G_1 \add_x_10_1/U29  ( .A1(\add_x_10_1/n51 ), .A2(\add_x_10_1/n49 ), .B(\add_x_10_1/n50 ), .X(\add_x_10_1/n48 ) );
  SEN_ND2_G_1 \add_x_10_1/U33  ( .A1(A[27]), .A2(B[27]), .X(\add_x_10_1/n50 )
         );
  SEN_NR2_1 \add_x_10_1/U32  ( .A1(A[27]), .A2(B[27]), .X(\add_x_10_1/n49 ) );
  SEN_ND2_G_1 \add_x_10_1/U41  ( .A1(A[26]), .A2(B[26]), .X(\add_x_10_1/n55 )
         );
  SEN_ND2_G_1 \add_x_10_1/U47  ( .A1(A[25]), .A2(B[25]), .X(\add_x_10_1/n58 )
         );
  SEN_NR2_1 \add_x_10_1/U46  ( .A1(A[25]), .A2(B[25]), .X(\add_x_10_1/n57 ) );
  SEN_ND2_G_1 \add_x_10_1/U55  ( .A1(A[24]), .A2(B[24]), .X(\add_x_10_1/n63 )
         );
  SEN_ND2_G_1 \add_x_10_1/U65  ( .A1(A[23]), .A2(B[23]), .X(\add_x_10_1/n70 )
         );
  SEN_OAI21_G_1 \add_x_10_1/U69  ( .A1(\add_x_10_1/n93 ), .A2(\add_x_10_1/n74 ), .B(\add_x_10_1/n75 ), .X(\add_x_10_1/n73 ) );
  SEN_ND2_G_1 \add_x_10_1/U77  ( .A1(A[22]), .A2(B[22]), .X(\add_x_10_1/n79 )
         );
  SEN_OAI21_G_1 \add_x_10_1/U81  ( .A1(\add_x_10_1/n83 ), .A2(\add_x_10_1/n87 ), .B(\add_x_10_1/n84 ), .X(\add_x_10_1/n82 ) );
  SEN_ND2_G_1 \add_x_10_1/U85  ( .A1(A[21]), .A2(B[21]), .X(\add_x_10_1/n84 )
         );
  SEN_ND2_G_1 \add_x_10_1/U91  ( .A1(A[20]), .A2(B[20]), .X(\add_x_10_1/n87 )
         );
  SEN_OAI21_G_1 \add_x_10_1/U100  ( .A1(\add_x_10_1/n96 ), .A2(
        \add_x_10_1/n100 ), .B(\add_x_10_1/n97 ), .X(\add_x_10_1/n95 ) );
  SEN_ND2_G_1 \add_x_10_1/U104  ( .A1(A[19]), .A2(B[19]), .X(\add_x_10_1/n97 )
         );
  SEN_ND2_G_1 \add_x_10_1/U110  ( .A1(A[18]), .A2(B[18]), .X(\add_x_10_1/n100 ) );
  SEN_OAI21_G_1 \add_x_10_1/U114  ( .A1(\add_x_10_1/n104 ), .A2(
        \add_x_10_1/n110 ), .B(\add_x_10_1/n105 ), .X(\add_x_10_1/n103 ) );
  SEN_ND2_G_1 \add_x_10_1/U118  ( .A1(A[17]), .A2(B[17]), .X(\add_x_10_1/n105 ) );
  SEN_ND2_G_1 \add_x_10_1/U126  ( .A1(A[16]), .A2(B[16]), .X(\add_x_10_1/n110 ) );
  SEN_ND2_G_1 \add_x_10_1/U58  ( .A1(\add_x_10_1/n72 ), .A2(n353), .X(
        \add_x_10_1/n65 ) );
  SEN_ND2_G_1 \add_x_10_1/U70  ( .A1(\add_x_10_1/n81 ), .A2(n354), .X(
        \add_x_10_1/n74 ) );
  SEN_NR2_1 \add_x_10_1/U84  ( .A1(A[21]), .A2(B[21]), .X(\add_x_10_1/n83 ) );
  SEN_NR2_1 \add_x_10_1/U90  ( .A1(A[20]), .A2(B[20]), .X(\add_x_10_1/n86 ) );
  SEN_ND2_G_1 \add_x_10_1/U97  ( .A1(\add_x_10_1/n102 ), .A2(\add_x_10_1/n94 ), 
        .X(\add_x_10_1/n92 ) );
  SEN_NR2_1 \add_x_10_1/U109  ( .A1(A[18]), .A2(B[18]), .X(\add_x_10_1/n99 )
         );
  SEN_NR2_1 \add_x_10_1/U117  ( .A1(A[17]), .A2(B[17]), .X(\add_x_10_1/n104 )
         );
  SEN_NR2_1 \add_x_10_1/U125  ( .A1(A[16]), .A2(B[16]), .X(\add_x_10_1/n109 )
         );
  SEN_OAI21_G_1 \add_x_10_1/U131  ( .A1(\add_x_10_1/n141 ), .A2(
        \add_x_10_1/n115 ), .B(\add_x_10_1/n116 ), .X(\add_x_10_1/n114 ) );
  SEN_OAI21_G_1 \add_x_10_1/U135  ( .A1(\add_x_10_1/n119 ), .A2(
        \add_x_10_1/n125 ), .B(\add_x_10_1/n120 ), .X(\add_x_10_1/n118 ) );
  SEN_ND2_G_1 \add_x_10_1/U139  ( .A1(A[15]), .A2(B[15]), .X(\add_x_10_1/n120 ) );
  SEN_ND2_G_1 \add_x_10_1/U147  ( .A1(A[14]), .A2(B[14]), .X(\add_x_10_1/n125 ) );
  SEN_OAI21_G_1 \add_x_10_1/U153  ( .A1(\add_x_10_1/n131 ), .A2(
        \add_x_10_1/n137 ), .B(\add_x_10_1/n132 ), .X(\add_x_10_1/n130 ) );
  SEN_ND2_G_1 \add_x_10_1/U157  ( .A1(A[13]), .A2(B[13]), .X(\add_x_10_1/n132 ) );
  SEN_ND2_G_1 \add_x_10_1/U165  ( .A1(A[12]), .A2(B[12]), .X(\add_x_10_1/n137 ) );
  SEN_OAI21_G_1 \add_x_10_1/U172  ( .A1(\add_x_10_1/n144 ), .A2(
        \add_x_10_1/n150 ), .B(\add_x_10_1/n145 ), .X(\add_x_10_1/n143 ) );
  SEN_ND2_G_1 \add_x_10_1/U176  ( .A1(A[11]), .A2(B[11]), .X(\add_x_10_1/n145 ) );
  SEN_ND2_G_1 \add_x_10_1/U184  ( .A1(A[10]), .A2(B[10]), .X(\add_x_10_1/n150 ) );
  SEN_OAI21_G_1 \add_x_10_1/U190  ( .A1(\add_x_10_1/n156 ), .A2(
        \add_x_10_1/n160 ), .B(\add_x_10_1/n157 ), .X(\add_x_10_1/n155 ) );
  SEN_ND2_G_1 \add_x_10_1/U194  ( .A1(A[9]), .A2(B[9]), .X(\add_x_10_1/n157 )
         );
  SEN_ND2_G_1 \add_x_10_1/U200  ( .A1(A[8]), .A2(B[8]), .X(\add_x_10_1/n160 )
         );
  SEN_NR2_1 \add_x_10_1/U130  ( .A1(\add_x_10_1/n140 ), .A2(\add_x_10_1/n115 ), 
        .X(\add_x_10_1/n113 ) );
  SEN_ND2_G_1 \add_x_10_1/U132  ( .A1(\add_x_10_1/n129 ), .A2(
        \add_x_10_1/n117 ), .X(\add_x_10_1/n115 ) );
  SEN_NR2_1 \add_x_10_1/U146  ( .A1(A[14]), .A2(B[14]), .X(\add_x_10_1/n124 )
         );
  SEN_NR2_1 \add_x_10_1/U164  ( .A1(A[12]), .A2(B[12]), .X(\add_x_10_1/n136 )
         );
  SEN_ND2_G_1 \add_x_10_1/U169  ( .A1(\add_x_10_1/n154 ), .A2(
        \add_x_10_1/n142 ), .X(\add_x_10_1/n140 ) );
  SEN_NR2_1 \add_x_10_1/U183  ( .A1(A[10]), .A2(B[10]), .X(\add_x_10_1/n149 )
         );
  SEN_NR2_1 \add_x_10_1/U193  ( .A1(A[9]), .A2(B[9]), .X(\add_x_10_1/n156 ) );
  SEN_OAI21_G_1 \add_x_10_1/U203  ( .A1(\add_x_10_1/n183 ), .A2(
        \add_x_10_1/n163 ), .B(\add_x_10_1/n164 ), .X(\add_x_10_1/n162 ) );
  SEN_OAI21_G_1 \add_x_10_1/U207  ( .A1(\add_x_10_1/n167 ), .A2(
        \add_x_10_1/n171 ), .B(\add_x_10_1/n168 ), .X(\add_x_10_1/n166 ) );
  SEN_ND2_G_1 \add_x_10_1/U211  ( .A1(A[7]), .A2(B[7]), .X(\add_x_10_1/n168 )
         );
  SEN_ND2_G_1 \add_x_10_1/U217  ( .A1(A[6]), .A2(B[6]), .X(\add_x_10_1/n171 )
         );
  SEN_OAI21_G_1 \add_x_10_1/U221  ( .A1(\add_x_10_1/n175 ), .A2(
        \add_x_10_1/n181 ), .B(\add_x_10_1/n176 ), .X(\add_x_10_1/n174 ) );
  SEN_ND2_G_1 \add_x_10_1/U225  ( .A1(A[5]), .A2(B[5]), .X(\add_x_10_1/n176 )
         );
  SEN_ND2_G_1 \add_x_10_1/U233  ( .A1(A[4]), .A2(B[4]), .X(\add_x_10_1/n181 )
         );
  SEN_ND2_G_1 \add_x_10_1/U204  ( .A1(\add_x_10_1/n173 ), .A2(
        \add_x_10_1/n165 ), .X(\add_x_10_1/n163 ) );
  SEN_NR2_1 \add_x_10_1/U216  ( .A1(A[6]), .A2(B[6]), .X(\add_x_10_1/n170 ) );
  SEN_NR2_1 \add_x_10_1/U224  ( .A1(A[5]), .A2(B[5]), .X(\add_x_10_1/n175 ) );
  SEN_NR2_1 \add_x_10_1/U232  ( .A1(A[4]), .A2(B[4]), .X(\add_x_10_1/n180 ) );
  SEN_OAI21_G_1 \add_x_10_1/U238  ( .A1(\add_x_10_1/n186 ), .A2(
        \add_x_10_1/n190 ), .B(\add_x_10_1/n187 ), .X(\add_x_10_1/n185 ) );
  SEN_ND2_G_1 \add_x_10_1/U242  ( .A1(A[3]), .A2(B[3]), .X(\add_x_10_1/n187 )
         );
  SEN_ND2_G_1 \add_x_10_1/U248  ( .A1(A[2]), .A2(B[2]), .X(\add_x_10_1/n190 )
         );
  SEN_OAI21_G_1 \add_x_10_1/U251  ( .A1(\add_x_10_1/n193 ), .A2(
        \add_x_10_1/n196 ), .B(\add_x_10_1/n194 ), .X(\add_x_10_1/n192 ) );
  SEN_ND2_G_1 \add_x_10_1/U255  ( .A1(A[1]), .A2(B[1]), .X(\add_x_10_1/n194 )
         );
  SEN_NR2_1 \add_x_10_1/U254  ( .A1(A[1]), .A2(B[1]), .X(\add_x_10_1/n193 ) );
  SEN_NR2_1 \add_x_10_1/U237  ( .A1(\add_x_10_1/n189 ), .A2(\add_x_10_1/n186 ), 
        .X(\add_x_10_1/n184 ) );
  SEN_NR2_1 \add_x_10_1/U241  ( .A1(A[3]), .A2(B[3]), .X(\add_x_10_1/n186 ) );
  SEN_NR2_1 \add_x_10_1/U247  ( .A1(A[2]), .A2(B[2]), .X(\add_x_10_1/n189 ) );
  SEN_ND2_G_1 \add_x_10_1/U2  ( .A1(n347), .A2(\add_x_10_1/n34 ), .X(
        \add_x_10_1/n1 ) );
  SEN_ND2_G_1 \add_x_10_1/U260  ( .A1(A[0]), .A2(B[0]), .X(\add_x_10_1/n196 )
         );
  SEN_EO2_S_0P5 \add_x_10_1/U249  ( .A1(\add_x_10_1/n196 ), .A2(
        \add_x_10_1/n31 ), .X(N125) );
  SEN_EN2_0P5 \add_x_10_1/U234  ( .A1(\add_x_10_1/n29 ), .A2(\add_x_10_1/n188 ), .X(N127) );
  SEN_EO2_S_0P5 \add_x_10_1/U218  ( .A1(\add_x_10_1/n27 ), .A2(
        \add_x_10_1/n177 ), .X(N129) );
  SEN_EN2_0P5 \add_x_10_1/U226  ( .A1(\add_x_10_1/n28 ), .A2(\add_x_10_1/n182 ), .X(N128) );
  SEN_EO2_S_0P5 \add_x_10_1/U243  ( .A1(\add_x_10_1/n30 ), .A2(
        \add_x_10_1/n191 ), .X(N126) );
  SEN_EN2_0P5 \add_x_10_1/U185  ( .A1(\add_x_10_1/n23 ), .A2(\add_x_10_1/n158 ), .X(N133) );
  SEN_EO2_S_0P5 \add_x_10_1/U212  ( .A1(\add_x_10_1/n26 ), .A2(
        \add_x_10_1/n172 ), .X(N130) );
  SEN_EN2_0P5 \add_x_10_1/U201  ( .A1(\add_x_10_1/n25 ), .A2(\add_x_10_1/n169 ), .X(N131) );
  SEN_EO2_S_0P5 \add_x_10_1/U195  ( .A1(\add_x_10_1/n24 ), .A2(
        \add_x_10_1/n161 ), .X(N132) );
  SEN_EO2_S_0P5 \add_x_10_1/U148  ( .A1(\add_x_10_1/n19 ), .A2(
        \add_x_10_1/n133 ), .X(N137) );
  SEN_EN2_0P5 \add_x_10_1/U177  ( .A1(\add_x_10_1/n22 ), .A2(\add_x_10_1/n151 ), .X(N134) );
  SEN_EO2_S_0P5 \add_x_10_1/U166  ( .A1(\add_x_10_1/n21 ), .A2(
        \add_x_10_1/n146 ), .X(N135) );
  SEN_EO2_S_0P5 \add_x_10_1/U158  ( .A1(\add_x_10_1/n20 ), .A2(
        \add_x_10_1/n138 ), .X(N136) );
  SEN_EN2_0P5 \add_x_10_1/U20  ( .A1(\add_x_10_1/n4 ), .A2(\add_x_10_1/n48 ), 
        .X(N152) );
  SEN_EN2_0P5 \add_x_10_1/U140  ( .A1(\add_x_10_1/n18 ), .A2(\add_x_10_1/n126 ), .X(N138) );
  SEN_EO2_S_0P5 \add_x_10_1/U111  ( .A1(\add_x_10_1/n15 ), .A2(
        \add_x_10_1/n106 ), .X(N141) );
  SEN_EN2_0P5 \add_x_10_1/U119  ( .A1(\add_x_10_1/n16 ), .A2(\add_x_10_1/n111 ), .X(N140) );
  SEN_EO2_S_0P5 \add_x_10_1/U42  ( .A1(\add_x_10_1/n7 ), .A2(\add_x_10_1/n59 ), 
        .X(N149) );
  SEN_EO2_S_0P5 \add_x_10_1/U105  ( .A1(\add_x_10_1/n14 ), .A2(
        \add_x_10_1/n101 ), .X(N142) );
  SEN_EO2_S_0P5 \add_x_10_1/U127  ( .A1(\add_x_10_1/n17 ), .A2(
        \add_x_10_1/n121 ), .X(N139) );
  SEN_EN2_0P5 \add_x_10_1/U78  ( .A1(\add_x_10_1/n11 ), .A2(\add_x_10_1/n85 ), 
        .X(N145) );
  SEN_EN2_0P5 \add_x_10_1/U92  ( .A1(\add_x_10_1/n13 ), .A2(\add_x_10_1/n98 ), 
        .X(N143) );
  SEN_EN2_0P5 \add_x_10_1/U86  ( .A1(\add_x_10_1/n12 ), .A2(\add_x_10_1/n88 ), 
        .X(N144) );
  SEN_EN2_0P5 \add_x_10_1/U6  ( .A1(\add_x_10_1/n2 ), .A2(\add_x_10_1/n40 ), 
        .X(N154) );
  SEN_EO2_S_0P5 \add_x_10_1/U66  ( .A1(\add_x_10_1/n10 ), .A2(\add_x_10_1/n80 ), .X(N146) );
  SEN_ND2_G_1 \cmp6_10_0/U34  ( .A1(\cmp6_10_0/n32 ), .A2(n346), .X(
        \cmp6_10_0/n26 ) );
  SEN_ND2_G_1 \cmp6_10_0/U13  ( .A1(n331), .A2(A[31]), .X(\cmp6_10_0/n5 ) );
  SEN_OAI21_G_1 \cmp6_10_0/U41  ( .A1(\cmp6_10_0/n73 ), .A2(\cmp6_10_0/n34 ), 
        .B(\cmp6_10_0/n35 ), .X(\cmp6_10_0/n33 ) );
  SEN_OAI21_G_1 \cmp6_10_0/U51  ( .A1(\cmp6_10_0/n59 ), .A2(\cmp6_10_0/n44 ), 
        .B(\cmp6_10_0/n45 ), .X(\cmp6_10_0/n43 ) );
  SEN_OAI21_G_1 \cmp6_10_0/U69  ( .A1(\cmp6_10_0/n62 ), .A2(\cmp6_10_0/n65 ), 
        .B(\cmp6_10_0/n63 ), .X(\cmp6_10_0/n61 ) );
  SEN_ND2_G_1 \cmp6_10_0/U52  ( .A1(\cmp6_10_0/n52 ), .A2(\cmp6_10_0/n46 ), 
        .X(\cmp6_10_0/n44 ) );
  SEN_OAI21_G_1 \cmp6_10_0/U83  ( .A1(\cmp6_10_0/n91 ), .A2(\cmp6_10_0/n76 ), 
        .B(\cmp6_10_0/n77 ), .X(\cmp6_10_0/n75 ) );
  SEN_ND2_G_1 \cmp6_10_0/U84  ( .A1(\cmp6_10_0/n84 ), .A2(\cmp6_10_0/n78 ), 
        .X(\cmp6_10_0/n76 ) );
  SEN_OAI21_G_1 \cmp6_10_0/U113  ( .A1(\cmp6_10_0/n121 ), .A2(\cmp6_10_0/n106 ), .B(\cmp6_10_0/n107 ), .X(\cmp6_10_0/n105 ) );
  SEN_ND2_G_1 \cmp6_10_0/U114  ( .A1(\cmp6_10_0/n114 ), .A2(\cmp6_10_0/n108 ), 
        .X(\cmp6_10_0/n106 ) );
  SEN_OAI21_G_1 \cmp6_10_0/U137  ( .A1(\cmp6_10_0/n133 ), .A2(\cmp6_10_0/n130 ), .B(\cmp6_10_0/n131 ), .X(\cmp6_10_0/n129 ) );
  SEN_EN2_0P5 \cmp6_10_0/U12  ( .A1(A[31]), .A2(n331), .X(\cmp6_10_0/n4 ) );
  SEN_EN2_0P5 \cmp6_10_0/U22  ( .A1(A[29]), .A2(n327), .X(\cmp6_10_0/n14 ) );
  SEN_EN2_0P5 \cmp6_10_0/U32  ( .A1(A[27]), .A2(n332), .X(\cmp6_10_0/n24 ) );
  SEN_AOI21_S_1 \cmp6_10_0/U43  ( .A1(\cmp6_10_0/n43 ), .A2(\cmp6_10_0/n36 ), 
        .B(\cmp6_10_0/n37 ), .X(\cmp6_10_0/n35 ) );
  SEN_AOI21_S_1 \cmp6_10_0/U53  ( .A1(\cmp6_10_0/n46 ), .A2(\cmp6_10_0/n53 ), 
        .B(\cmp6_10_0/n47 ), .X(\cmp6_10_0/n45 ) );
  SEN_AOI21_S_1 \cmp6_10_0/U67  ( .A1(\cmp6_10_0/n60 ), .A2(\cmp6_10_0/n67 ), 
        .B(\cmp6_10_0/n61 ), .X(\cmp6_10_0/n59 ) );
  SEN_EN2_0P5 \cmp6_10_0/U46  ( .A1(A[25]), .A2(n330), .X(\cmp6_10_0/n38 ) );
  SEN_EN2_0P5 \cmp6_10_0/U48  ( .A1(A[24]), .A2(n336), .X(\cmp6_10_0/n40 ) );
  SEN_EN2_0P5 \cmp6_10_0/U58  ( .A1(A[22]), .A2(n320), .X(\cmp6_10_0/n50 ) );
  SEN_EN2_0P5 \cmp6_10_0/U62  ( .A1(A[21]), .A2(n317), .X(\cmp6_10_0/n54 ) );
  SEN_EN2_0P5 \cmp6_10_0/U64  ( .A1(A[20]), .A2(n314), .X(\cmp6_10_0/n56 ) );
  SEN_EN2_0P5 \cmp6_10_0/U70  ( .A1(A[19]), .A2(n311), .X(\cmp6_10_0/n62 ) );
  SEN_EN2_0P5 \cmp6_10_0/U72  ( .A1(A[18]), .A2(n310), .X(\cmp6_10_0/n64 ) );
  SEN_EN2_0P5 \cmp6_10_0/U76  ( .A1(A[17]), .A2(n315), .X(\cmp6_10_0/n68 ) );
  SEN_AOI21_S_1 \cmp6_10_0/U81  ( .A1(\cmp6_10_0/n105 ), .A2(\cmp6_10_0/n74 ), 
        .B(\cmp6_10_0/n75 ), .X(\cmp6_10_0/n73 ) );
  SEN_AOI21_S_1 \cmp6_10_0/U85  ( .A1(\cmp6_10_0/n78 ), .A2(\cmp6_10_0/n85 ), 
        .B(\cmp6_10_0/n79 ), .X(\cmp6_10_0/n77 ) );
  SEN_AOI21_S_1 \cmp6_10_0/U99  ( .A1(\cmp6_10_0/n92 ), .A2(\cmp6_10_0/n99 ), 
        .B(\cmp6_10_0/n93 ), .X(\cmp6_10_0/n91 ) );
  SEN_EN2_0P5 \cmp6_10_0/U96  ( .A1(A[12]), .A2(n313), .X(\cmp6_10_0/n88 ) );
  SEN_EN2_0P5 \cmp6_10_0/U104  ( .A1(A[10]), .A2(n326), .X(\cmp6_10_0/n96 ) );
  SEN_EN2_0P5 \cmp6_10_0/U108  ( .A1(A[9]), .A2(n312), .X(\cmp6_10_0/n100 ) );
  SEN_AOI21_S_1 \cmp6_10_0/U115  ( .A1(\cmp6_10_0/n108 ), .A2(\cmp6_10_0/n115 ), .B(\cmp6_10_0/n109 ), .X(\cmp6_10_0/n107 ) );
  SEN_EN2_0P5 \cmp6_10_0/U120  ( .A1(A[6]), .A2(n323), .X(\cmp6_10_0/n112 ) );
  SEN_EN2_0P5 \cmp6_10_0/U124  ( .A1(A[5]), .A2(n322), .X(\cmp6_10_0/n116 ) );
  SEN_EN2_0P5 \cmp6_10_0/U126  ( .A1(A[4]), .A2(n328), .X(\cmp6_10_0/n118 ) );
  SEN_AOI21_S_1 \cmp6_10_0/U129  ( .A1(\cmp6_10_0/n129 ), .A2(\cmp6_10_0/n122 ), .B(\cmp6_10_0/n123 ), .X(\cmp6_10_0/n121 ) );
  SEN_EN2_0P5 \cmp6_10_0/U134  ( .A1(A[2]), .A2(n337), .X(\cmp6_10_0/n126 ) );
  SEN_EN2_0P5 \cmp6_10_0/U138  ( .A1(A[1]), .A2(n307), .X(\cmp6_10_0/n130 ) );
  SEN_NR2_G_1 \add_x_10_1/U210  ( .A1(A[7]), .A2(B[7]), .X(\add_x_10_1/n167 )
         );
  SEN_NR2_G_1 \add_x_10_1/U175  ( .A1(A[11]), .A2(B[11]), .X(\add_x_10_1/n144 ) );
  SEN_NR2_G_1 \add_x_10_1/U156  ( .A1(A[13]), .A2(B[13]), .X(\add_x_10_1/n131 ) );
  SEN_NR2_G_1 \add_x_10_1/U138  ( .A1(A[15]), .A2(B[15]), .X(\add_x_10_1/n119 ) );
  SEN_NR2_G_1 \sub_x_10_3/U199  ( .A1(n329), .A2(A[8]), .X(\sub_x_10_3/n158 )
         );
  SEN_NR2_G_1 \cmp6_10_0/U44  ( .A1(\cmp6_10_0/n40 ), .A2(\cmp6_10_0/n38 ), 
        .X(\cmp6_10_0/n36 ) );
  SEN_NR2_G_1 \add_x_10_1/U206  ( .A1(\add_x_10_1/n170 ), .A2(
        \add_x_10_1/n167 ), .X(\add_x_10_1/n165 ) );
  SEN_NR2_G_1 \add_x_10_1/U152  ( .A1(\add_x_10_1/n136 ), .A2(
        \add_x_10_1/n131 ), .X(\add_x_10_1/n129 ) );
  SEN_NR2_G_1 \sub_x_10_3/U84  ( .A1(n317), .A2(A[21]), .X(\sub_x_10_3/n82 )
         );
  SEN_NR2_G_1 \sub_x_10_3/U103  ( .A1(n311), .A2(A[19]), .X(\sub_x_10_3/n95 )
         );
  SEN_NR2_G_1 \sub_x_10_3/U175  ( .A1(n316), .A2(A[11]), .X(\sub_x_10_3/n143 )
         );
  SEN_ND2_S_1 \add_x_10_2/U44  ( .A1(\add_x_10_2/n36 ), .A2(\add_x_10_2/n33 ), 
        .X(\add_x_10_2/n32 ) );
  SEN_NR2_G_1 \sub_x_10_3/U117  ( .A1(n315), .A2(A[17]), .X(\sub_x_10_3/n103 )
         );
  SEN_NR2_G_1 \add_x_10_1/U99  ( .A1(\add_x_10_1/n99 ), .A2(\add_x_10_1/n96 ), 
        .X(\add_x_10_1/n94 ) );
  SEN_NR2_G_1 \add_x_10_1/U171  ( .A1(\add_x_10_1/n149 ), .A2(
        \add_x_10_1/n144 ), .X(\add_x_10_1/n142 ) );
  SEN_NR2_G_1 \sub_x_10_3/U210  ( .A1(n324), .A2(A[7]), .X(\sub_x_10_3/n166 )
         );
  SEN_NR2_G_1 \sub_x_10_3/U146  ( .A1(n308), .A2(A[14]), .X(\sub_x_10_3/n123 )
         );
  SEN_NR2_G_1 \sub_x_10_3/U193  ( .A1(n312), .A2(A[9]), .X(\sub_x_10_3/n155 )
         );
  SEN_NR2_G_1 \add_x_10_1/U189  ( .A1(\add_x_10_1/n159 ), .A2(
        \add_x_10_1/n156 ), .X(\add_x_10_1/n154 ) );
  SEN_NR2_G_1 \sub_x_10_3/U156  ( .A1(n318), .A2(A[13]), .X(\sub_x_10_3/n130 )
         );
  SEN_NR2_G_1 \sub_x_10_3/U138  ( .A1(n309), .A2(A[15]), .X(\sub_x_10_3/n118 )
         );
  SEN_AOI21_G_1 \add_x_10_1/U236  ( .A1(\add_x_10_1/n184 ), .A2(
        \add_x_10_1/n192 ), .B(\add_x_10_1/n185 ), .X(\add_x_10_1/n183 ) );
  SEN_NR2_G_1 \sub_x_10_3/U99  ( .A1(\sub_x_10_3/n98 ), .A2(\sub_x_10_3/n95 ), 
        .X(\sub_x_10_3/n93 ) );
  SEN_NR2_G_1 \cmp6_10_0/U122  ( .A1(\cmp6_10_0/n118 ), .A2(\cmp6_10_0/n116 ), 
        .X(\cmp6_10_0/n114 ) );
  SEN_OAI21_1 \cmp6_10_0/U131  ( .A1(\cmp6_10_0/n124 ), .A2(\cmp6_10_0/n127 ), 
        .B(\cmp6_10_0/n125 ), .X(\cmp6_10_0/n123 ) );
  SEN_NR2_G_1 \sub_x_10_3/U189  ( .A1(\sub_x_10_3/n158 ), .A2(
        \sub_x_10_3/n155 ), .X(\sub_x_10_3/n153 ) );
  SEN_AOI21_G_1 \add_x_10_1/U71  ( .A1(\add_x_10_1/n82 ), .A2(n354), .B(
        \add_x_10_1/n77 ), .X(\add_x_10_1/n75 ) );
  SEN_NR2_G_1 \sub_x_10_3/U113  ( .A1(\sub_x_10_3/n108 ), .A2(
        \sub_x_10_3/n103 ), .X(\sub_x_10_3/n101 ) );
  SEN_NR2_G_1 \cmp6_10_0/U141  ( .A1(\cmp6_10_0/n134 ), .A2(n343), .X(
        \cmp6_10_0/n133 ) );
  SEN_NR2_G_1 \sub_x_10_3/U206  ( .A1(\sub_x_10_3/n169 ), .A2(
        \sub_x_10_3/n166 ), .X(\sub_x_10_3/n164 ) );
  SEN_NR2_G_1 \add_x_10_2/U110  ( .A1(\add_x_10_2/n94 ), .A2(\add_x_10_2/n87 ), 
        .X(\add_x_10_2/n86 ) );
  SEN_AOI21_G_1 \add_x_10_1/U133  ( .A1(\add_x_10_1/n117 ), .A2(
        \add_x_10_1/n130 ), .B(\add_x_10_1/n118 ), .X(\add_x_10_1/n116 ) );
  SEN_AOI21_G_1 \add_x_10_1/U170  ( .A1(\add_x_10_1/n142 ), .A2(
        \add_x_10_1/n155 ), .B(\add_x_10_1/n143 ), .X(\add_x_10_1/n141 ) );
  SEN_AOI21_G_1 \add_x_10_1/U205  ( .A1(\add_x_10_1/n165 ), .A2(
        \add_x_10_1/n174 ), .B(\add_x_10_1/n166 ), .X(\add_x_10_1/n164 ) );
  SEN_NR2_G_1 \sub_x_10_3/U152  ( .A1(\sub_x_10_3/n135 ), .A2(
        \sub_x_10_3/n130 ), .X(\sub_x_10_3/n128 ) );
  SEN_NR2_G_1 \cmp6_10_0/U54  ( .A1(\cmp6_10_0/n50 ), .A2(\cmp6_10_0/n48 ), 
        .X(\cmp6_10_0/n46 ) );
  SEN_NR2_G_1 \cmp6_10_0/U86  ( .A1(\cmp6_10_0/n82 ), .A2(\cmp6_10_0/n80 ), 
        .X(\cmp6_10_0/n78 ) );
  SEN_NR2_G_1 \add_x_10_2/U43  ( .A1(\add_x_10_2/n39 ), .A2(\add_x_10_2/n32 ), 
        .X(\add_x_10_2/n31 ) );
  SEN_NR2_G_1 \cmp6_10_0/U92  ( .A1(\cmp6_10_0/n88 ), .A2(\cmp6_10_0/n86 ), 
        .X(\cmp6_10_0/n84 ) );
  SEN_NR2_G_1 \cmp6_10_0/U68  ( .A1(\cmp6_10_0/n64 ), .A2(\cmp6_10_0/n62 ), 
        .X(\cmp6_10_0/n60 ) );
  SEN_NR2_G_1 \cmp6_10_0/U60  ( .A1(\cmp6_10_0/n56 ), .A2(\cmp6_10_0/n54 ), 
        .X(\cmp6_10_0/n52 ) );
  SEN_NR2_G_1 \add_x_10_2/U65  ( .A1(\add_x_10_2/n59 ), .A2(\add_x_10_2/n50 ), 
        .X(\add_x_10_2/n49 ) );
  SEN_NR2_G_1 \sub_x_10_3/U171  ( .A1(\sub_x_10_3/n148 ), .A2(
        \sub_x_10_3/n143 ), .X(\sub_x_10_3/n141 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U71  ( .A1(\sub_x_10_3/n81 ), .A2(n361), .B(
        \sub_x_10_3/n76 ), .X(\sub_x_10_3/n74 ) );
  SEN_AOI21_G_1 \add_x_10_1/U59  ( .A1(\add_x_10_1/n73 ), .A2(n353), .B(
        \add_x_10_1/n68 ), .X(\add_x_10_1/n66 ) );
  SEN_NR2_G_1 \add_x_10_2/U29  ( .A1(\add_x_10_2/n23 ), .A2(A[22]), .X(
        \add_x_10_2/n20 ) );
  SEN_AOI21_G_1 \add_x_10_1/U219  ( .A1(\add_x_10_1/n182 ), .A2(
        \add_x_10_1/n173 ), .B(\add_x_10_1/n174 ), .X(\add_x_10_1/n172 ) );
  SEN_AOI21_G_1 \add_x_10_1/U227  ( .A1(\add_x_10_1/n182 ), .A2(
        \add_x_10_1/n224 ), .B(\add_x_10_1/n179 ), .X(\add_x_10_1/n177 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U219  ( .A1(\sub_x_10_3/n181 ), .A2(
        \sub_x_10_3/n172 ), .B(\sub_x_10_3/n173 ), .X(\sub_x_10_3/n171 ) );
  SEN_ND2_S_1 \add_x_10_2/U115  ( .A1(\add_x_10_2/n93 ), .A2(\add_x_10_2/n91 ), 
        .X(\add_x_10_2/n90 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U227  ( .A1(\sub_x_10_3/n181 ), .A2(
        \sub_x_10_3/n222 ), .B(\sub_x_10_3/n178 ), .X(\sub_x_10_3/n176 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U59  ( .A1(\sub_x_10_3/n72 ), .A2(n360), .B(
        \sub_x_10_3/n67 ), .X(\sub_x_10_3/n65 ) );
  SEN_AOI21_G_1 \add_x_10_1/U159  ( .A1(\add_x_10_1/n139 ), .A2(
        \add_x_10_1/n216 ), .B(\add_x_10_1/n135 ), .X(\add_x_10_1/n133 ) );
  SEN_NR2_G_1 \add_x_10_2/U52  ( .A1(\add_x_10_2/n46 ), .A2(\add_x_10_2/n39 ), 
        .X(\add_x_10_2/n38 ) );
  SEN_AOI21_G_1 \add_x_10_1/U120  ( .A1(\add_x_10_1/n111 ), .A2(
        \add_x_10_1/n212 ), .B(\add_x_10_1/n108 ), .X(\add_x_10_1/n106 ) );
  SEN_AOI21_G_1 \add_x_10_1/U112  ( .A1(\add_x_10_1/n111 ), .A2(
        \add_x_10_1/n102 ), .B(\add_x_10_1/n103 ), .X(\add_x_10_1/n101 ) );
  SEN_AOI21_G_1 \add_x_10_1/U94  ( .A1(\add_x_10_1/n111 ), .A2(
        \add_x_10_1/n90 ), .B(\add_x_10_1/n91 ), .X(\add_x_10_1/n89 ) );
  SEN_AOI21_G_1 \add_x_10_1/U178  ( .A1(\add_x_10_1/n151 ), .A2(
        \add_x_10_1/n218 ), .B(\add_x_10_1/n148 ), .X(\add_x_10_1/n146 ) );
  SEN_NR2_G_1 \cmp6_10_0/U40  ( .A1(\cmp6_10_0/n72 ), .A2(\cmp6_10_0/n34 ), 
        .X(\cmp6_10_0/n32 ) );
  SEN_NR2_G_1 \add_x_10_2/U93  ( .A1(\add_x_10_2/n76 ), .A2(A[10]), .X(
        \add_x_10_2/n72 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U120  ( .A1(\sub_x_10_3/n110 ), .A2(
        \sub_x_10_3/n210 ), .B(\sub_x_10_3/n107 ), .X(\sub_x_10_3/n105 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U112  ( .A1(\sub_x_10_3/n110 ), .A2(
        \sub_x_10_3/n101 ), .B(\sub_x_10_3/n102 ), .X(\sub_x_10_3/n100 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U159  ( .A1(\sub_x_10_3/n138 ), .A2(
        \sub_x_10_3/n214 ), .B(\sub_x_10_3/n134 ), .X(\sub_x_10_3/n132 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U178  ( .A1(\sub_x_10_3/n150 ), .A2(
        \sub_x_10_3/n216 ), .B(\sub_x_10_3/n147 ), .X(\sub_x_10_3/n145 ) );
  SEN_AOI21_G_1 \add_x_10_1/U141  ( .A1(\add_x_10_1/n126 ), .A2(
        \add_x_10_1/n214 ), .B(\add_x_10_1/n123 ), .X(\add_x_10_1/n121 ) );
  SEN_AOI21_G_1 \add_x_10_1/U79  ( .A1(\add_x_10_1/n88 ), .A2(\add_x_10_1/n81 ), .B(\add_x_10_1/n82 ), .X(\add_x_10_1/n80 ) );
  SEN_NR2_G_1 \add_x_10_2/U70  ( .A1(\add_x_10_2/n57 ), .A2(A[14]), .X(
        \add_x_10_2/n53 ) );
  SEN_NR2_G_1 \cmp6_10_0/U30  ( .A1(\cmp6_10_0/n26 ), .A2(\cmp6_10_0/n24 ), 
        .X(\cmp6_10_0/n22 ) );
  SEN_NR2_G_1 \add_x_10_2/U18  ( .A1(\add_x_10_2/n14 ), .A2(A[25]), .X(
        \add_x_10_2/n12 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U79  ( .A1(\sub_x_10_3/n87 ), .A2(\sub_x_10_3/n80 ), .B(\sub_x_10_3/n81 ), .X(\sub_x_10_3/n79 ) );
  SEN_AOI21_G_1 \sub_x_10_3/U141  ( .A1(\sub_x_10_3/n125 ), .A2(
        \sub_x_10_3/n212 ), .B(\sub_x_10_3/n122 ), .X(\sub_x_10_3/n120 ) );
  SEN_NR2_G_1 \cmp6_10_0/U20  ( .A1(\cmp6_10_0/n16 ), .A2(\cmp6_10_0/n14 ), 
        .X(\cmp6_10_0/n12 ) );
  SEN_NR2_G_1 \add_x_10_2/U11  ( .A1(\add_x_10_2/n9 ), .A2(A[27]), .X(
        \add_x_10_2/n7 ) );
  SEN_AOI21_G_1 \add_x_10_1/U7  ( .A1(\add_x_10_1/n40 ), .A2(n349), .B(
        \add_x_10_1/n37 ), .X(\add_x_10_1/n35 ) );
  SEN_AN2_1 \cmp6_10_0/U5  ( .A1(N56), .A2(N57), .X(N53) );
  SEN_NR2_G_1 \sub_x_10_3/U257  ( .A1(A[0]), .A2(n339), .X(\sub_x_10_3/n194 )
         );
  SEN_NR2_G_1 \add_x_10_1/U134  ( .A1(\add_x_10_1/n124 ), .A2(
        \add_x_10_1/n119 ), .X(\add_x_10_1/n117 ) );
  SEN_NR2_G_1 \add_x_10_1/U103  ( .A1(A[19]), .A2(B[19]), .X(\add_x_10_1/n96 )
         );
  SEN_NR2_G_1 \add_x_10_1/U113  ( .A1(\add_x_10_1/n109 ), .A2(
        \add_x_10_1/n104 ), .X(\add_x_10_1/n102 ) );
  SEN_NR2_G_1 \add_x_10_1/U220  ( .A1(\add_x_10_1/n180 ), .A2(
        \add_x_10_1/n175 ), .X(\add_x_10_1/n173 ) );
  SEN_NR2_G_1 \sub_x_10_3/U134  ( .A1(\sub_x_10_3/n123 ), .A2(
        \sub_x_10_3/n118 ), .X(\sub_x_10_3/n116 ) );
  SEN_NR2_G_1 \sub_x_10_3/U220  ( .A1(\sub_x_10_3/n179 ), .A2(
        \sub_x_10_3/n174 ), .X(\sub_x_10_3/n172 ) );
  SEN_NR2_G_1 \sub_x_10_3/U80  ( .A1(\sub_x_10_3/n85 ), .A2(\sub_x_10_3/n82 ), 
        .X(\sub_x_10_3/n80 ) );
  SEN_NR2_1 \add_x_10_1/U68  ( .A1(\add_x_10_1/n92 ), .A2(\add_x_10_1/n74 ), 
        .X(\add_x_10_1/n72 ) );
  SEN_NR2_1 \add_x_10_2/U119  ( .A1(\add_x_10_2/n101 ), .A2(\add_x_10_2/n94 ), 
        .X(\add_x_10_2/n93 ) );
  SEN_NR2_1 \sub_x_10_3/U68  ( .A1(\sub_x_10_3/n91 ), .A2(\sub_x_10_3/n73 ), 
        .X(\sub_x_10_3/n71 ) );
  SEN_NR2_G_1 \add_x_10_1/U199  ( .A1(A[8]), .A2(B[8]), .X(\add_x_10_1/n159 )
         );
  SEN_NR2_1 \sub_x_10_3/U125  ( .A1(n325), .A2(A[16]), .X(\sub_x_10_3/n108 )
         );
  SEN_ND2_G_0P65 \add_x_10_1/U24  ( .A1(n350), .A2(\add_x_10_1/n47 ), .X(
        \add_x_10_1/n4 ) );
  SEN_ND2_0P8 \cmp6_10_0/U135  ( .A1(n337), .A2(A[2]), .X(\cmp6_10_0/n127 ) );
  SEN_ND2_S_0P5 \cmp6_10_0/U33  ( .A1(n332), .A2(A[27]), .X(\cmp6_10_0/n25 )
         );
  SEN_NR2_G_1 \sub_x_10_3/U216  ( .A1(n323), .A2(A[6]), .X(\sub_x_10_3/n169 )
         );
  SEN_NR2_G_1 \add_x_10_1/U80  ( .A1(\add_x_10_1/n86 ), .A2(\add_x_10_1/n83 ), 
        .X(\add_x_10_1/n81 ) );
  SEN_NR2_G_1 \sub_x_10_3/U164  ( .A1(n313), .A2(A[12]), .X(\sub_x_10_3/n135 )
         );
  SEN_OAI21_S_1 \cmp6_10_0/U87  ( .A1(\cmp6_10_0/n80 ), .A2(\cmp6_10_0/n83 ), 
        .B(\cmp6_10_0/n81 ), .X(\cmp6_10_0/n79 ) );
  SEN_NR2_G_1 \sub_x_10_3/U224  ( .A1(n322), .A2(A[5]), .X(\sub_x_10_3/n174 )
         );
  SEN_NR2_G_1 \sub_x_10_3/U109  ( .A1(n310), .A2(A[18]), .X(\sub_x_10_3/n98 )
         );
  SEN_ND2_G_0P65 \add_x_10_2/U135  ( .A1(\add_x_10_2/n109 ), .A2(
        \add_x_10_2/n107 ), .X(\add_x_10_2/n106 ) );
  SEN_ND2_S_1 \add_x_10_2/U104  ( .A1(\add_x_10_2/n84 ), .A2(\add_x_10_2/n82 ), 
        .X(\add_x_10_2/n81 ) );
  SEN_ND2_S_1 \add_x_10_2/U48  ( .A1(\add_x_10_2/n38 ), .A2(\add_x_10_2/n36 ), 
        .X(\add_x_10_2/n35 ) );
  SEN_ND2_G_1 \cmp6_10_0/U24  ( .A1(\cmp6_10_0/n22 ), .A2(n345), .X(
        \cmp6_10_0/n16 ) );
  SEN_ND2_S_0P65 \add_x_10_1/U5  ( .A1(A[31]), .A2(B[31]), .X(\add_x_10_1/n34 ) );
  SEN_ND2_0P5 \cmp6_10_0/U79  ( .A1(n325), .A2(A[16]), .X(\cmp6_10_0/n71 ) );
  SEN_ND2_0P5 \cmp6_10_0/U91  ( .A1(n308), .A2(A[14]), .X(\cmp6_10_0/n83 ) );
  SEN_ND2_0P5 \sub_x_10_3/U5  ( .A1(n331), .A2(A[31]), .X(\sub_x_10_3/n33 ) );
  SEN_ND2_0P5 \cmp6_10_0/U105  ( .A1(n326), .A2(A[10]), .X(\cmp6_10_0/n97 ) );
  SEN_ND2_S_0P8 \cmp6_10_0/U23  ( .A1(n327), .A2(A[29]), .X(\cmp6_10_0/n15 )
         );
  SEN_ND2_0P5 \cmp6_10_0/U89  ( .A1(n309), .A2(A[15]), .X(\cmp6_10_0/n81 ) );
  SEN_NR2_1 \sub_x_10_3/U90  ( .A1(n314), .A2(A[20]), .X(\sub_x_10_3/n85 ) );
  SEN_ND2_S_1 \add_x_10_2/U66  ( .A1(\add_x_10_2/n55 ), .A2(\add_x_10_2/n51 ), 
        .X(\add_x_10_2/n50 ) );
  SEN_ND2_G_0P65 \add_x_10_1/U44  ( .A1(\add_x_10_1/n203 ), .A2(
        \add_x_10_1/n58 ), .X(\add_x_10_1/n7 ) );
  SEN_ND2_0P5 \cmp6_10_0/U133  ( .A1(n321), .A2(A[3]), .X(\cmp6_10_0/n125 ) );
  SEN_ND2_0P5 \cmp6_10_0/U95  ( .A1(n318), .A2(A[13]), .X(\cmp6_10_0/n87 ) );
  SEN_ND2_0P5 \cmp6_10_0/U97  ( .A1(n313), .A2(A[12]), .X(\cmp6_10_0/n89 ) );
  SEN_NR2_1 \sub_x_10_3/U241  ( .A1(n321), .A2(A[3]), .X(\sub_x_10_3/n185 ) );
  SEN_ND2_0P5 \cmp6_10_0/U103  ( .A1(n316), .A2(A[11]), .X(\cmp6_10_0/n95 ) );
  SEN_ND2_0P5 \cmp6_10_0/U77  ( .A1(n315), .A2(A[17]), .X(\cmp6_10_0/n69 ) );
  SEN_ND2_0P5 \cmp6_10_0/U139  ( .A1(n307), .A2(A[1]), .X(\cmp6_10_0/n131 ) );
  SEN_ND2_0P5 \cmp6_10_0/U73  ( .A1(n310), .A2(A[18]), .X(\cmp6_10_0/n65 ) );
  SEN_ND2_0P5 \cmp6_10_0/U71  ( .A1(n311), .A2(A[19]), .X(\cmp6_10_0/n63 ) );
  SEN_ND2_G_0P65 \sub_x_10_3/U44  ( .A1(\sub_x_10_3/n201 ), .A2(
        \sub_x_10_3/n57 ), .X(\sub_x_10_3/n7 ) );
  SEN_OAI21_0P75 \cmp6_10_0/U101  ( .A1(\cmp6_10_0/n94 ), .A2(\cmp6_10_0/n97 ), 
        .B(\cmp6_10_0/n95 ), .X(\cmp6_10_0/n93 ) );
  SEN_OAI21_0P75 \cmp6_10_0/U93  ( .A1(\cmp6_10_0/n86 ), .A2(\cmp6_10_0/n89 ), 
        .B(\cmp6_10_0/n87 ), .X(\cmp6_10_0/n85 ) );
  SEN_NR2_1 \add_x_10_2/U63  ( .A1(\add_x_10_2/n48 ), .A2(\add_x_10_2/n85 ), 
        .X(\add_x_10_2/n47 ) );
  SEN_ND2_G_1 \add_x_10_2/U37  ( .A1(\add_x_10_2/n29 ), .A2(\add_x_10_2/n27 ), 
        .X(\add_x_10_2/n26 ) );
  SEN_EN2_0P5 U263 ( .A1(A[15]), .A2(n309), .X(\cmp6_10_0/n80 ) );
  SEN_EO2_S_0P5 U264 ( .A1(\add_x_10_2/A[31] ), .A2(\add_x_10_2/n1 ), .X(N187)
         );
  SEN_EN2_0P5 U265 ( .A1(A[11]), .A2(n316), .X(\cmp6_10_0/n94 ) );
  SEN_EN2_0P5 U266 ( .A1(A[13]), .A2(n318), .X(\cmp6_10_0/n86 ) );
  SEN_EN2_0P5 U267 ( .A1(A[14]), .A2(n308), .X(\cmp6_10_0/n82 ) );
  SEN_EN2_0P5 U268 ( .A1(A[23]), .A2(n319), .X(\cmp6_10_0/n48 ) );
  SEN_EN2_0P5 U269 ( .A1(A[3]), .A2(n321), .X(\cmp6_10_0/n124 ) );
  SEN_INV_S_1 U270 ( .A(B[7]), .X(n324) );
  SEN_INV_S_1 U271 ( .A(B[12]), .X(n313) );
  SEN_INV_S_1 U272 ( .A(B[13]), .X(n318) );
  SEN_INV_S_1 U273 ( .A(n387), .X(n385) );
  SEN_INV_S_1 U274 ( .A(n365), .X(n363) );
  SEN_INV_S_1 U275 ( .A(B[21]), .X(n317) );
  SEN_INV_S_1 U276 ( .A(n387), .X(n386) );
  SEN_INV_S_1 U277 ( .A(n365), .X(n364) );
  SEN_AOI211_0P5 U278 ( .A1(N187), .A2(n383), .B1(n610), .B2(n609), .X(n614)
         );
  SEN_EO2_S_0P5 U279 ( .A1(A[23]), .A2(\add_x_10_2/n19 ), .X(n229) );
  SEN_OAOI211_0P5 U280 ( .A1(A[23]), .A2(n371), .B(n367), .C(n319), .X(n230)
         );
  SEN_NR2_0P5 U281 ( .A1(n371), .A2(B[23]), .X(n231) );
  SEN_AOI211_0P5 U282 ( .A1(B[23]), .A2(n376), .B1(n373), .B2(n231), .X(n232)
         );
  SEN_INV_0P5 U283 ( .A(A[23]), .X(n233) );
  SEN_AOI22_0P5 U284 ( .A1(A[23]), .A2(n232), .B1(n381), .B2(n233), .X(n234)
         );
  SEN_AOI211_0P5 U285 ( .A1(n383), .A2(n229), .B1(n230), .B2(n234), .X(n235)
         );
  SEN_AOI21_0P5 U286 ( .A1(\add_x_10_1/n72 ), .A2(\add_x_10_1/n111 ), .B(
        \add_x_10_1/n73 ), .X(n236) );
  SEN_ND2_0P5 U287 ( .A1(n353), .A2(\add_x_10_1/n70 ), .X(n237) );
  SEN_ND2_0P5 U288 ( .A1(n237), .A2(n236), .X(n238) );
  SEN_OAI211_0P5 U289 ( .A1(n237), .A2(n236), .B1(n238), .B2(n386), .X(n239)
         );
  SEN_AOI21_0P5 U290 ( .A1(\sub_x_10_3/n71 ), .A2(\sub_x_10_3/n110 ), .B(
        \sub_x_10_3/n72 ), .X(n240) );
  SEN_ND2_0P5 U291 ( .A1(n360), .A2(\sub_x_10_3/n69 ), .X(n241) );
  SEN_ND2_0P5 U292 ( .A1(n241), .A2(n240), .X(n242) );
  SEN_OAI211_0P5 U293 ( .A1(n241), .A2(n240), .B1(n242), .B2(n364), .X(n243)
         );
  SEN_ND3_S_0P5 U294 ( .A1(n235), .A2(n239), .A3(n243), .X(Z[23]) );
  SEN_AOI21_S_1 U295 ( .A1(A[8]), .A2(n329), .B(\cmp6_10_0/n100 ), .X(n244) );
  SEN_OAI211_0P5 U296 ( .A1(A[8]), .A2(n329), .B1(\cmp6_10_0/n92 ), .B2(n244), 
        .X(n245) );
  SEN_NR2_1 U297 ( .A1(\cmp6_10_0/n76 ), .A2(n245), .X(\cmp6_10_0/n74 ) );
  SEN_AN3B_1 U298 ( .B1(\add_x_10_2/n107 ), .B2(\add_x_10_2/n104 ), .A(
        \add_x_10_2/n110 ), .X(\add_x_10_2/n102 ) );
  SEN_AOI21B_1 U299 ( .A1(\add_x_10_1/n56 ), .A2(n351), .B(\add_x_10_1/n55 ), 
        .X(\add_x_10_1/n51 ) );
  SEN_AOAI211_0P5 U300 ( .A1(n352), .A2(\add_x_10_1/n63 ), .B(\add_x_10_1/n64 ), .C(n386), .X(n246) );
  SEN_AOI31_0P5 U301 ( .A1(\add_x_10_1/n64 ), .A2(n352), .A3(\add_x_10_1/n63 ), 
        .B(n246), .X(n247) );
  SEN_AOAI211_0P5 U302 ( .A1(n359), .A2(\sub_x_10_3/n62 ), .B(\sub_x_10_3/n63 ), .C(n364), .X(n248) );
  SEN_AOI31_0P5 U303 ( .A1(\sub_x_10_3/n63 ), .A2(n359), .A3(\sub_x_10_3/n62 ), 
        .B(n248), .X(n249) );
  SEN_EN2_0P5 U304 ( .A1(A[24]), .A2(\add_x_10_2/n17 ), .X(n250) );
  SEN_OAOI211_0P5 U305 ( .A1(A[24]), .A2(n370), .B(n367), .C(n336), .X(n251)
         );
  SEN_NR2_0P5 U306 ( .A1(n371), .A2(B[24]), .X(n252) );
  SEN_AOI211_0P5 U307 ( .A1(B[24]), .A2(n376), .B1(n373), .B2(n252), .X(n253)
         );
  SEN_INV_0P5 U308 ( .A(\add_x_10_2/n15 ), .X(n254) );
  SEN_AOI22_0P5 U309 ( .A1(\add_x_10_2/n15 ), .A2(n381), .B1(n253), .B2(n254), 
        .X(n255) );
  SEN_AOI211_0P5 U310 ( .A1(n383), .A2(n250), .B1(n251), .B2(n255), .X(n256)
         );
  SEN_OR3B_0P5 U311 ( .B1(n247), .B2(n249), .A(n256), .X(Z[24]) );
  SEN_NR4B_1 U312 ( .A(\cmp6_10_0/n122 ), .B1(\cmp6_10_0/n132 ), .B2(
        \cmp6_10_0/n130 ), .B3(\cmp6_10_0/n106 ), .X(n257) );
  SEN_ND2_0P5 U313 ( .A1(\cmp6_10_0/n74 ), .A2(n257), .X(\cmp6_10_0/n72 ) );
  SEN_ND2B_1 U314 ( .A(\add_x_10_2/n78 ), .B(\add_x_10_2/n84 ), .X(
        \add_x_10_2/n76 ) );
  SEN_ND2B_1 U315 ( .A(\add_x_10_2/n59 ), .B(\add_x_10_2/n66 ), .X(
        \add_x_10_2/n57 ) );
  SEN_OA21_1 U316 ( .A1(n258), .A2(\sub_x_10_3/n91 ), .B(\sub_x_10_3/n92 ), 
        .X(\sub_x_10_3/n88 ) );
  SEN_INV_0P5 U317 ( .A(\sub_x_10_3/n110 ), .X(n258) );
  SEN_ND2B_1 U318 ( .A(\add_x_10_1/n41 ), .B(\add_x_10_1/n42 ), .X(
        \add_x_10_1/n3 ) );
  SEN_NR2_1 U319 ( .A1(\add_x_10_2/n4 ), .A2(A[29]), .X(n259) );
  SEN_EO2_S_0P5 U320 ( .A1(n259), .A2(\add_x_10_2/A[30] ), .X(N186) );
  SEN_AN2_1 U321 ( .A1(n259), .A2(\add_x_10_2/A[30] ), .X(\add_x_10_2/n1 ) );
  SEN_EO2_S_0P5 U322 ( .A1(A[27]), .A2(\add_x_10_2/n9 ), .X(n260) );
  SEN_OAOI211_0P5 U323 ( .A1(A[27]), .A2(n370), .B(n367), .C(n332), .X(n261)
         );
  SEN_AOI211_0P5 U324 ( .A1(B[27]), .A2(n376), .B1(n586), .B2(n373), .X(n262)
         );
  SEN_INV_0P5 U325 ( .A(A[27]), .X(n263) );
  SEN_AOI22_0P5 U326 ( .A1(A[27]), .A2(n262), .B1(n381), .B2(n263), .X(n264)
         );
  SEN_AOI211_0P5 U327 ( .A1(n383), .A2(n260), .B1(n261), .B2(n264), .X(n265)
         );
  SEN_ND2B_1 U328 ( .A(\add_x_10_1/n49 ), .B(\add_x_10_1/n50 ), .X(n266) );
  SEN_ND2_0P5 U329 ( .A1(n266), .A2(\add_x_10_1/n51 ), .X(n267) );
  SEN_OAI211_0P5 U330 ( .A1(\add_x_10_1/n51 ), .A2(n266), .B1(n267), .B2(n386), 
        .X(n268) );
  SEN_ND2B_1 U331 ( .A(\sub_x_10_3/n48 ), .B(\sub_x_10_3/n49 ), .X(n269) );
  SEN_ND2_0P5 U332 ( .A1(n269), .A2(\sub_x_10_3/n50 ), .X(n270) );
  SEN_OAI211_0P5 U333 ( .A1(\sub_x_10_3/n50 ), .A2(n269), .B1(n270), .B2(n364), 
        .X(n271) );
  SEN_ND3_S_0P5 U334 ( .A1(n265), .A2(n268), .A3(n271), .X(Z[27]) );
  SEN_ND2_0P5 U335 ( .A1(A[4]), .A2(n328), .X(n272) );
  SEN_AO2BB2_0P5 U336 ( .A1(\cmp6_10_0/n116 ), .A2(n272), .B1(A[5]), .B2(n322), 
        .X(\cmp6_10_0/n115 ) );
  SEN_ND2_0P5 U337 ( .A1(A[20]), .A2(n314), .X(n273) );
  SEN_AO2BB2_0P5 U338 ( .A1(\cmp6_10_0/n54 ), .A2(n273), .B1(A[21]), .B2(n317), 
        .X(\cmp6_10_0/n53 ) );
  SEN_OAI21_G_1 U339 ( .A1(n325), .A2(A[16]), .B(\cmp6_10_0/n60 ), .X(n274) );
  SEN_AOI211_G_1 U340 ( .A1(n325), .A2(A[16]), .B1(\cmp6_10_0/n68 ), .B2(n274), 
        .X(n275) );
  SEN_ND3B_1 U341 ( .A(\cmp6_10_0/n44 ), .B1(n275), .B2(\cmp6_10_0/n36 ), .X(
        \cmp6_10_0/n34 ) );
  SEN_AN3B_0P5 U342 ( .B1(INST[1]), .B2(n408), .A(n404), .X(n606) );
  SEN_INV_0P5 U343 ( .A(\add_x_10_1/n154 ), .X(n276) );
  SEN_OAI21B_0P5 U344 ( .A1(\add_x_10_1/n161 ), .A2(n276), .B(
        \add_x_10_1/n155 ), .X(\add_x_10_1/n151 ) );
  SEN_INV_0P5 U345 ( .A(\add_x_10_1/n129 ), .X(n277) );
  SEN_OAI21B_0P5 U346 ( .A1(\add_x_10_1/n138 ), .A2(n277), .B(
        \add_x_10_1/n130 ), .X(\add_x_10_1/n126 ) );
  SEN_NR2B_1 U347 ( .A(\add_x_10_2/n31 ), .B(\add_x_10_2/n46 ), .X(
        \add_x_10_2/n29 ) );
  SEN_AOI21B_1 U348 ( .A1(\sub_x_10_3/n63 ), .A2(n359), .B(\sub_x_10_3/n62 ), 
        .X(\sub_x_10_3/n58 ) );
  SEN_OAOI211_0P5 U349 ( .A1(A[29]), .A2(n369), .B(n367), .C(n327), .X(n278)
         );
  SEN_AOI211_0P5 U350 ( .A1(n383), .A2(N185), .B1(n278), .B2(n596), .X(n279)
         );
  SEN_ND2_0P5 U351 ( .A1(\add_x_10_1/n3 ), .A2(\add_x_10_1/n43 ), .X(n280) );
  SEN_OAI211_0P5 U352 ( .A1(\add_x_10_1/n3 ), .A2(\add_x_10_1/n43 ), .B1(n280), 
        .B2(n386), .X(n281) );
  SEN_ND2_0P5 U353 ( .A1(\sub_x_10_3/n3 ), .A2(\sub_x_10_3/n42 ), .X(n282) );
  SEN_OAI211_0P5 U354 ( .A1(\sub_x_10_3/n3 ), .A2(\sub_x_10_3/n42 ), .B1(n282), 
        .B2(n364), .X(n283) );
  SEN_ND3_S_0P5 U355 ( .A1(n279), .A2(n281), .A3(n283), .X(Z[29]) );
  SEN_ND2_0P5 U356 ( .A1(A[6]), .A2(n323), .X(n284) );
  SEN_AO2BB2_0P5 U357 ( .A1(\cmp6_10_0/n110 ), .A2(n284), .B1(A[7]), .B2(n324), 
        .X(\cmp6_10_0/n109 ) );
  SEN_ND2_0P5 U358 ( .A1(A[8]), .A2(n329), .X(n285) );
  SEN_AO2BB2_0P5 U359 ( .A1(\cmp6_10_0/n100 ), .A2(n285), .B1(A[9]), .B2(n312), 
        .X(\cmp6_10_0/n99 ) );
  SEN_ND2_0P5 U360 ( .A1(A[22]), .A2(n320), .X(n286) );
  SEN_AO2BB2_0P5 U361 ( .A1(\cmp6_10_0/n48 ), .A2(n286), .B1(A[23]), .B2(n319), 
        .X(\cmp6_10_0/n47 ) );
  SEN_ND2_0P5 U362 ( .A1(A[24]), .A2(n336), .X(n287) );
  SEN_AO2BB2_0P5 U363 ( .A1(\cmp6_10_0/n38 ), .A2(n287), .B1(A[25]), .B2(n330), 
        .X(\cmp6_10_0/n37 ) );
  SEN_AN3B_0P5 U364 ( .B1(\add_x_10_2/n70 ), .B2(\add_x_10_2/n74 ), .A(
        \add_x_10_2/n78 ), .X(\add_x_10_2/n68 ) );
  SEN_INV_0P5 U365 ( .A(INST[1]), .X(n288) );
  SEN_AOI22_0P5 U366 ( .A1(INST[1]), .A2(N57), .B1(N56), .B2(n288), .X(n289)
         );
  SEN_AOI21_0P5 U367 ( .A1(N54), .A2(n288), .B(n393), .X(n290) );
  SEN_AOAI211_0P5 U368 ( .A1(n393), .A2(n289), .B(n290), .C(INST[2]), .X(n391)
         );
  SEN_INV_0P5 U369 ( .A(\sub_x_10_3/n153 ), .X(n291) );
  SEN_OAI21B_0P5 U370 ( .A1(\sub_x_10_3/n160 ), .A2(n291), .B(
        \sub_x_10_3/n154 ), .X(\sub_x_10_3/n150 ) );
  SEN_OAI21B_0P5 U371 ( .A1(\sub_x_10_3/n137 ), .A2(n292), .B(
        \sub_x_10_3/n129 ), .X(\sub_x_10_3/n125 ) );
  SEN_INV_0P5 U372 ( .A(\sub_x_10_3/n128 ), .X(n292) );
  SEN_OR3B_0P5 U373 ( .B1(A[21]), .B2(A[20]), .A(\add_x_10_2/n31 ), .X(
        \add_x_10_2/n23 ) );
  SEN_AO21B_1 U374 ( .A1(n334), .A2(A[28]), .B(n357), .X(\sub_x_10_3/n4 ) );
  SEN_ND2B_1 U375 ( .A(\sub_x_10_3/n40 ), .B(\sub_x_10_3/n41 ), .X(
        \sub_x_10_3/n3 ) );
  SEN_AOAI211_0P5 U376 ( .A1(n351), .A2(\add_x_10_1/n55 ), .B(\add_x_10_1/n56 ), .C(n386), .X(n293) );
  SEN_AOI31_0P5 U377 ( .A1(\add_x_10_1/n56 ), .A2(n351), .A3(\add_x_10_1/n55 ), 
        .B(n293), .X(n294) );
  SEN_ND2_0P5 U378 ( .A1(n333), .A2(A[26]), .X(n295) );
  SEN_AOAI211_0P5 U379 ( .A1(n358), .A2(n295), .B(\sub_x_10_3/n55 ), .C(n364), 
        .X(n296) );
  SEN_AOI31_0P5 U380 ( .A1(\sub_x_10_3/n55 ), .A2(n358), .A3(n295), .B(n296), 
        .X(n297) );
  SEN_EN2_0P5 U381 ( .A1(\add_x_10_2/n12 ), .A2(A[26]), .X(n298) );
  SEN_OAOI211_0P5 U382 ( .A1(A[26]), .A2(n370), .B(n367), .C(n333), .X(n299)
         );
  SEN_NR2_0P5 U383 ( .A1(n371), .A2(B[26]), .X(n300) );
  SEN_AOI211_0P5 U384 ( .A1(B[26]), .A2(n376), .B1(n373), .B2(n300), .X(n301)
         );
  SEN_INV_0P5 U385 ( .A(\add_x_10_2/n10 ), .X(n302) );
  SEN_AOI22_0P5 U386 ( .A1(\add_x_10_2/n10 ), .A2(n381), .B1(n301), .B2(n302), 
        .X(n303) );
  SEN_AOI211_0P5 U387 ( .A1(n611), .A2(n298), .B1(n299), .B2(n303), .X(n304)
         );
  SEN_OR3B_0P5 U388 ( .B1(n294), .B2(n297), .A(n304), .X(Z[26]) );
  SEN_ND2_0P5 U389 ( .A1(N378), .A2(n602), .X(n305) );
  SEN_AOI211_0P5 U390 ( .A1(n383), .A2(N186), .B1(n600), .B2(n599), .X(n306)
         );
  SEN_ND3_S_0P5 U391 ( .A1(n305), .A2(n306), .A3(n601), .X(Z[30]) );
  SEN_ND2_S_1 U392 ( .A1(N154), .A2(n612), .X(n601) );
  SEN_NR2_T_1 U393 ( .A1(\cmp6_10_0/n6 ), .A2(\cmp6_10_0/n4 ), .X(N54) );
  SEN_OAI21_S_2 U394 ( .A1(\add_x_10_1/n59 ), .A2(\add_x_10_1/n57 ), .B(
        \add_x_10_1/n58 ), .X(\add_x_10_1/n56 ) );
  SEN_OAOI211_1 U395 ( .A1(A[25]), .A2(n370), .B(n367), .C(n330), .X(n582) );
  SEN_OAOI211_1 U396 ( .A1(A[22]), .A2(n371), .B(n367), .C(n320), .X(n575) );
  SEN_AOI211_0P5 U397 ( .A1(n376), .A2(B[30]), .B1(n373), .B2(n597), .X(n598)
         );
  SEN_NR2_G_0P5 U398 ( .A1(n372), .A2(B[10]), .X(n488) );
  SEN_NR2_0P65 U399 ( .A1(n371), .A2(B[29]), .X(n594) );
  SEN_INV_0P8 U400 ( .A(\add_x_10_2/n110 ), .X(\add_x_10_2/n109 ) );
  SEN_INV_0P8 U401 ( .A(\sub_x_10_3/n174 ), .X(\sub_x_10_3/n221 ) );
  SEN_INV_0P8 U402 ( .A(\sub_x_10_3/n185 ), .X(\sub_x_10_3/n223 ) );
  SEN_INV_0P8 U403 ( .A(\sub_x_10_3/n95 ), .X(\sub_x_10_3/n207 ) );
  SEN_INV_0P8 U404 ( .A(n409), .X(n405) );
  SEN_INV_0P8 U405 ( .A(\sub_x_10_3/n85 ), .X(\sub_x_10_3/n206 ) );
  SEN_INV_0P8 U406 ( .A(\add_x_10_1/n86 ), .X(\add_x_10_1/n208 ) );
  SEN_INV_0P65 U407 ( .A(\sub_x_10_3/n56 ), .X(\sub_x_10_3/n201 ) );
  SEN_INV_0P8 U408 ( .A(\sub_x_10_3/n118 ), .X(\sub_x_10_3/n211 ) );
  SEN_EN2_S_1 U409 ( .A1(A[7]), .A2(n324), .X(\cmp6_10_0/n110 ) );
  SEN_INV_0P8 U410 ( .A(\add_x_10_1/n186 ), .X(\add_x_10_1/n225 ) );
  SEN_INV_1 U411 ( .A(B[22]), .X(n320) );
  SEN_INV_2 U412 ( .A(B[1]), .X(n307) );
  SEN_INV_0P8 U413 ( .A(\add_x_10_1/n119 ), .X(\add_x_10_1/n213 ) );
  SEN_AN2_1 U414 ( .A1(n335), .A2(A[30]), .X(n340) );
  SEN_INV_1 U415 ( .A(B[15]), .X(n309) );
  SEN_INV_1 U416 ( .A(B[14]), .X(n308) );
  SEN_INV_1 U417 ( .A(B[0]), .X(n339) );
  SEN_ND2_G_0P65 U418 ( .A1(INST[0]), .A2(INST[2]), .X(n399) );
  SEN_INV_1 U419 ( .A(B[2]), .X(n337) );
  SEN_INV_1 U420 ( .A(N56), .X(N52) );
  SEN_ND2_G_1 U421 ( .A1(N363), .A2(n364), .X(n529) );
  SEN_ND2_G_1 U422 ( .A1(\cmp6_10_0/n12 ), .A2(n344), .X(\cmp6_10_0/n6 ) );
  SEN_ND2_G_1 U423 ( .A1(N370), .A2(n364), .X(n578) );
  SEN_OAI21_S_2 U424 ( .A1(\cmp6_10_0/n17 ), .A2(\cmp6_10_0/n14 ), .B(
        \cmp6_10_0/n15 ), .X(\cmp6_10_0/n13 ) );
  SEN_ND2_G_1 U425 ( .A1(N367), .A2(n364), .X(n557) );
  SEN_ND2_G_1 U426 ( .A1(N362), .A2(n363), .X(n522) );
  SEN_ND2_G_1 U427 ( .A1(N146), .A2(n386), .X(n576) );
  SEN_ND2_G_1 U428 ( .A1(N139), .A2(n386), .X(n527) );
  SEN_ND2_G_1 U429 ( .A1(N369), .A2(n364), .X(n571) );
  SEN_ND2_G_1 U430 ( .A1(N368), .A2(n364), .X(n564) );
  SEN_ND2_G_1 U431 ( .A1(N365), .A2(n364), .X(n543) );
  SEN_ND2_G_1 U432 ( .A1(N361), .A2(n363), .X(n515) );
  SEN_ND2_G_1 U433 ( .A1(N144), .A2(n386), .X(n562) );
  SEN_ND2_G_1 U434 ( .A1(N366), .A2(n364), .X(n550) );
  SEN_ND2_G_1 U435 ( .A1(N138), .A2(n385), .X(n520) );
  SEN_ND2_G_1 U436 ( .A1(N360), .A2(n363), .X(n508) );
  SEN_ND2_G_1 U437 ( .A1(N359), .A2(n363), .X(n501) );
  SEN_ND2_G_1 U438 ( .A1(N373), .A2(n364), .X(n585) );
  SEN_ND2_G_1 U439 ( .A1(N145), .A2(n386), .X(n569) );
  SEN_ND2_G_1 U440 ( .A1(N143), .A2(n386), .X(n555) );
  SEN_ND2_G_1 U441 ( .A1(N357), .A2(n363), .X(n487) );
  SEN_ND2_G_1 U442 ( .A1(N136), .A2(n385), .X(n506) );
  SEN_ND2_G_1 U443 ( .A1(N141), .A2(n386), .X(n541) );
  SEN_ND2_G_1 U444 ( .A1(N137), .A2(n385), .X(n513) );
  SEN_ND2_G_1 U445 ( .A1(N135), .A2(n385), .X(n499) );
  SEN_ND2_G_1 U446 ( .A1(N355), .A2(n363), .X(n473) );
  SEN_ND2_G_1 U447 ( .A1(N142), .A2(n386), .X(n548) );
  SEN_ND2_G_1 U448 ( .A1(N149), .A2(n386), .X(n583) );
  SEN_ND2_G_1 U449 ( .A1(N364), .A2(n364), .X(n536) );
  SEN_ND2_G_1 U450 ( .A1(N358), .A2(n363), .X(n494) );
  SEN_OAOI211_1 U451 ( .A1(A[19]), .A2(n371), .B(n367), .C(n311), .X(n554) );
  SEN_ND2_G_1 U452 ( .A1(N354), .A2(n363), .X(n466) );
  SEN_ND2_G_1 U453 ( .A1(N134), .A2(n385), .X(n492) );
  SEN_OAOI211_1 U454 ( .A1(A[21]), .A2(n371), .B(n367), .C(n317), .X(n568) );
  SEN_OAOI211_1 U455 ( .A1(A[20]), .A2(n371), .B(n367), .C(n314), .X(n561) );
  SEN_ND2_G_1 U456 ( .A1(N353), .A2(n363), .X(n459) );
  SEN_ND2_G_1 U457 ( .A1(N356), .A2(n363), .X(n480) );
  SEN_ND2_G_1 U458 ( .A1(N133), .A2(n385), .X(n485) );
  SEN_OAOI211_1 U459 ( .A1(A[7]), .A2(n369), .B(n366), .C(n324), .X(n470) );
  SEN_ND2_G_1 U460 ( .A1(N131), .A2(n385), .X(n471) );
  SEN_ND2_G_1 U461 ( .A1(N140), .A2(n386), .X(n534) );
  SEN_ND2_G_1 U462 ( .A1(N130), .A2(n385), .X(n464) );
  SEN_ND2_G_1 U463 ( .A1(N132), .A2(n385), .X(n478) );
  SEN_ND2_G_1 U464 ( .A1(N351), .A2(n363), .X(n445) );
  SEN_AOI211_0P5 U465 ( .A1(n376), .A2(B[28]), .B1(n373), .B2(n587), .X(n588)
         );
  SEN_ND2_G_1 U466 ( .A1(N129), .A2(n385), .X(n457) );
  SEN_ND2_G_1 U467 ( .A1(N352), .A2(n363), .X(n452) );
  SEN_OAI21_S_2 U468 ( .A1(\sub_x_10_3/n111 ), .A2(\sub_x_10_3/n64 ), .B(
        \sub_x_10_3/n65 ), .X(\sub_x_10_3/n63 ) );
  SEN_AOI211_0P5 U469 ( .A1(n376), .A2(B[29]), .B1(n373), .B2(n594), .X(n595)
         );
  SEN_NR2_T_1 U470 ( .A1(\add_x_10_2/n19 ), .A2(A[23]), .X(\add_x_10_2/n17 )
         );
  SEN_OAOI211_0P5 U471 ( .A1(A[28]), .A2(n370), .B(n603), .C(n334), .X(n590)
         );
  SEN_ND2_G_1 U472 ( .A1(N349), .A2(n363), .X(n430) );
  SEN_ND2_G_1 U473 ( .A1(N127), .A2(n385), .X(n443) );
  SEN_ND2_G_1 U474 ( .A1(N350), .A2(n363), .X(n438) );
  SEN_NR2_G_0P8 U475 ( .A1(n372), .A2(B[1]), .X(n423) );
  SEN_ND2_G_1 U476 ( .A1(N128), .A2(n385), .X(n450) );
  SEN_ND2_G_1 U477 ( .A1(N125), .A2(n385), .X(n429) );
  SEN_ND2_G_1 U478 ( .A1(N126), .A2(n385), .X(n436) );
  SEN_NR2_G_1 U479 ( .A1(\cmp6_10_0/n112 ), .A2(\cmp6_10_0/n110 ), .X(
        \cmp6_10_0/n108 ) );
  SEN_OAI21_G_1 U480 ( .A1(\sub_x_10_3/n103 ), .A2(\sub_x_10_3/n109 ), .B(
        \sub_x_10_3/n104 ), .X(\sub_x_10_3/n102 ) );
  SEN_INV_0P8 U481 ( .A(\sub_x_10_3/n103 ), .X(\sub_x_10_3/n209 ) );
  SEN_INV_0P8 U482 ( .A(\sub_x_10_3/n98 ), .X(\sub_x_10_3/n208 ) );
  SEN_INV_0P8 U483 ( .A(\sub_x_10_3/n169 ), .X(\sub_x_10_3/n220 ) );
  SEN_INV_0P8 U484 ( .A(\sub_x_10_3/n155 ), .X(\sub_x_10_3/n217 ) );
  SEN_NR2_G_1 U485 ( .A1(\cmp6_10_0/n126 ), .A2(\cmp6_10_0/n124 ), .X(
        \cmp6_10_0/n122 ) );
  SEN_INV_0P8 U486 ( .A(\sub_x_10_3/n143 ), .X(\sub_x_10_3/n215 ) );
  SEN_INV_0P8 U487 ( .A(\sub_x_10_3/n166 ), .X(\sub_x_10_3/n219 ) );
  SEN_INV_0P8 U488 ( .A(\add_x_10_1/n96 ), .X(\add_x_10_1/n209 ) );
  SEN_INV_0P8 U489 ( .A(\add_x_10_1/n175 ), .X(\add_x_10_1/n223 ) );
  SEN_INV_0P8 U490 ( .A(\add_x_10_1/n170 ), .X(\add_x_10_1/n222 ) );
  SEN_INV_0P8 U491 ( .A(\add_x_10_1/n144 ), .X(\add_x_10_1/n217 ) );
  SEN_INV_0P8 U492 ( .A(\add_x_10_1/n167 ), .X(\add_x_10_1/n221 ) );
  SEN_AN2_DG_1 U493 ( .A1(n334), .A2(A[28]), .X(n341) );
  SEN_INV_1 U494 ( .A(B[20]), .X(n314) );
  SEN_AN2_S_0P5 U495 ( .A1(n333), .A2(A[26]), .X(n342) );
  SEN_INV_1 U496 ( .A(B[23]), .X(n319) );
  SEN_EN2_1 U497 ( .A1(A[0]), .A2(n339), .X(\cmp6_10_0/n132 ) );
  SEN_INV_0P8 U498 ( .A(\add_x_10_1/n57 ), .X(\add_x_10_1/n203 ) );
  SEN_INV_1 U499 ( .A(B[10]), .X(n326) );
  SEN_INV_1 U500 ( .A(B[16]), .X(n325) );
  SEN_INV_1 U501 ( .A(B[31]), .X(n331) );
  SEN_INV_1 U502 ( .A(B[24]), .X(n336) );
  SEN_INV_1 U503 ( .A(B[25]), .X(n330) );
  SEN_INV_1 U504 ( .A(B[26]), .X(n333) );
  SEN_INV_1 U505 ( .A(B[27]), .X(n332) );
  SEN_INV_1 U506 ( .A(B[28]), .X(n334) );
  SEN_INV_1 U507 ( .A(B[29]), .X(n327) );
  SEN_INV_1 U508 ( .A(B[30]), .X(n335) );
  SEN_INV_1 U509 ( .A(B[8]), .X(n329) );
  SEN_INV_1 U510 ( .A(B[4]), .X(n328) );
  SEN_AOI21_G_2 U511 ( .A1(\cmp6_10_0/n13 ), .A2(n344), .B(n340), .X(
        \cmp6_10_0/n7 ) );
  SEN_AOI211_G_0P5 U512 ( .A1(N181), .A2(n383), .B1(n582), .B2(n581), .X(n584)
         );
  SEN_OAI21_S_1P5 U513 ( .A1(\cmp6_10_0/n27 ), .A2(\cmp6_10_0/n24 ), .B(
        \cmp6_10_0/n25 ), .X(\cmp6_10_0/n23 ) );
  SEN_AOI211_G_0P5 U514 ( .A1(N172), .A2(n382), .B1(n533), .B2(n532), .X(n535)
         );
  SEN_AOI211_G_0P5 U515 ( .A1(N176), .A2(n383), .B1(n561), .B2(n560), .X(n563)
         );
  SEN_AOI211_G_0P5 U516 ( .A1(N173), .A2(n382), .B1(n540), .B2(n539), .X(n542)
         );
  SEN_AOI211_G_0P5 U517 ( .A1(N174), .A2(n382), .B1(n547), .B2(n546), .X(n549)
         );
  SEN_NR2_G_0P5 U518 ( .A1(n372), .A2(B[12]), .X(n502) );
  SEN_NR2_G_0P5 U519 ( .A1(n372), .A2(B[14]), .X(n516) );
  SEN_NR2_G_0P5 U520 ( .A1(n372), .A2(B[15]), .X(n523) );
  SEN_NR2_G_0P5 U521 ( .A1(n372), .A2(B[16]), .X(n530) );
  SEN_NR2_G_0P5 U522 ( .A1(n372), .A2(B[11]), .X(n495) );
  SEN_NR2_G_0P5 U523 ( .A1(n372), .A2(B[13]), .X(n509) );
  SEN_NR2_G_0P5 U524 ( .A1(n372), .A2(B[9]), .X(n481) );
  SEN_NR2_G_0P5 U525 ( .A1(n372), .A2(B[21]), .X(n565) );
  SEN_NR2_G_0P5 U526 ( .A1(n371), .A2(B[22]), .X(n572) );
  SEN_ND2_S_1 U527 ( .A1(\add_x_10_2/n47 ), .A2(\add_x_10_2/n20 ), .X(
        \add_x_10_2/n19 ) );
  SEN_NR2_G_0P5 U528 ( .A1(n372), .A2(B[20]), .X(n558) );
  SEN_NR2_G_0P5 U529 ( .A1(n371), .A2(B[27]), .X(n586) );
  SEN_NR2_G_0P5 U530 ( .A1(n372), .A2(B[19]), .X(n551) );
  SEN_NR2_G_0P5 U531 ( .A1(n372), .A2(B[18]), .X(n544) );
  SEN_NR2_G_0P5 U532 ( .A1(n371), .A2(B[28]), .X(n587) );
  SEN_NR2_G_0P5 U533 ( .A1(n371), .A2(B[25]), .X(n579) );
  SEN_NR2_G_0P5 U534 ( .A1(n372), .A2(B[17]), .X(n537) );
  SEN_INV_1 U535 ( .A(n338), .X(n369) );
  SEN_INV_1 U536 ( .A(n338), .X(n370) );
  SEN_INV_1 U537 ( .A(n338), .X(n371) );
  SEN_INV_1 U538 ( .A(n338), .X(n372) );
  SEN_AOI22_0P5 U539 ( .A1(n338), .A2(A[0]), .B1(SEL), .B2(n425), .X(n417) );
  SEN_INV_1 U540 ( .A(n604), .X(n338) );
  SEN_NR2_S_0P5 U541 ( .A1(n604), .A2(B[6]), .X(n460) );
  SEN_AOI21_G_1 U542 ( .A1(\sub_x_10_3/n93 ), .A2(\sub_x_10_3/n102 ), .B(
        \sub_x_10_3/n94 ), .X(\sub_x_10_3/n92 ) );
  SEN_NR2_S_0P5 U543 ( .A1(n604), .A2(B[8]), .X(n474) );
  SEN_NR2_S_0P5 U544 ( .A1(n604), .A2(B[7]), .X(n467) );
  SEN_NR2_S_0P5 U545 ( .A1(n604), .A2(B[5]), .X(n453) );
  SEN_INV_1 U546 ( .A(n380), .X(n379) );
  SEN_NR2_S_0P5 U547 ( .A1(n604), .A2(B[4]), .X(n446) );
  SEN_INV_0P8 U548 ( .A(\sub_x_10_3/n130 ), .X(\sub_x_10_3/n213 ) );
  SEN_NR2_G_1 U549 ( .A1(\cmp6_10_0/n96 ), .A2(\cmp6_10_0/n94 ), .X(
        \cmp6_10_0/n92 ) );
  SEN_INV_0P8 U550 ( .A(\add_x_10_1/n156 ), .X(\add_x_10_1/n219 ) );
  SEN_INV_0P8 U551 ( .A(\add_x_10_1/n99 ), .X(\add_x_10_1/n210 ) );
  SEN_INV_0P8 U552 ( .A(\sub_x_10_3/n158 ), .X(\sub_x_10_3/n218 ) );
  SEN_INV_0P8 U553 ( .A(\add_x_10_1/n104 ), .X(\add_x_10_1/n211 ) );
  SEN_INV_0P65 U554 ( .A(\cmp6_10_0/n132 ), .X(\cmp6_10_0/n134 ) );
  SEN_INV_0P8 U555 ( .A(\add_x_10_1/n159 ), .X(\add_x_10_1/n220 ) );
  SEN_INV_2 U556 ( .A(B[18]), .X(n310) );
  SEN_INV_2 U557 ( .A(B[19]), .X(n311) );
  SEN_INV_2 U558 ( .A(B[9]), .X(n312) );
  SEN_INV_2 U559 ( .A(B[17]), .X(n315) );
  SEN_INV_2 U560 ( .A(B[11]), .X(n316) );
  SEN_INV_2 U561 ( .A(B[3]), .X(n321) );
  SEN_INV_2 U562 ( .A(B[5]), .X(n322) );
  SEN_INV_2 U563 ( .A(B[6]), .X(n323) );
  SEN_AN2_1 U564 ( .A1(INST[2]), .A2(SEL), .X(n394) );
  SEN_ND3_T_0P65 U565 ( .A1(n615), .A2(n614), .A3(n613), .X(Z[31]) );
  SEN_OR2_1 U566 ( .A1(N52), .A2(N54), .X(N55) );
  SEN_EO2_1 U567 ( .A1(\sub_x_10_3/n1 ), .A2(\sub_x_10_3/n34 ), .X(N379) );
  SEN_ND2_G_1 U568 ( .A1(N155), .A2(n612), .X(n613) );
  SEN_INV_1 U569 ( .A(N54), .X(N57) );
  SEN_AOI21_G_2 U570 ( .A1(\sub_x_10_3/n39 ), .A2(n356), .B(n340), .X(
        \sub_x_10_3/n34 ) );
  SEN_OAI21_S_3 U571 ( .A1(\cmp6_10_0/n7 ), .A2(\cmp6_10_0/n4 ), .B(
        \cmp6_10_0/n5 ), .X(N56) );
  SEN_AOI21_G_2 U572 ( .A1(\sub_x_10_3/n47 ), .A2(n357), .B(n341), .X(
        \sub_x_10_3/n42 ) );
  SEN_AOI21_G_2 U573 ( .A1(\add_x_10_1/n48 ), .A2(n350), .B(\add_x_10_1/n45 ), 
        .X(\add_x_10_1/n43 ) );
  SEN_AOI21_G_2 U574 ( .A1(\cmp6_10_0/n23 ), .A2(n345), .B(n341), .X(
        \cmp6_10_0/n17 ) );
  SEN_AOI211_G_0P5 U575 ( .A1(N170), .A2(n382), .B1(n519), .B2(n518), .X(n521)
         );
  SEN_AOI21_G_2 U576 ( .A1(\sub_x_10_3/n55 ), .A2(n358), .B(n342), .X(
        \sub_x_10_3/n50 ) );
  SEN_AOI211_G_0P5 U577 ( .A1(N164), .A2(n382), .B1(n477), .B2(n476), .X(n479)
         );
  SEN_AOI211_G_0P5 U578 ( .A1(N178), .A2(n382), .B1(n575), .B2(n574), .X(n577)
         );
  SEN_AOI211_G_0P5 U579 ( .A1(N162), .A2(n382), .B1(n463), .B2(n462), .X(n465)
         );
  SEN_AOI211_G_0P5 U580 ( .A1(N168), .A2(n382), .B1(n505), .B2(n504), .X(n507)
         );
  SEN_AOI211_G_0P5 U581 ( .A1(N159), .A2(n383), .B1(n442), .B2(n441), .X(n444)
         );
  SEN_AOI211_G_0P5 U582 ( .A1(N158), .A2(n383), .B1(n435), .B2(n434), .X(n437)
         );
  SEN_AOI211_G_0P5 U583 ( .A1(N166), .A2(n382), .B1(n491), .B2(n490), .X(n493)
         );
  SEN_AOI211_G_0P5 U584 ( .A1(n383), .A2(N157), .B1(n428), .B2(n427), .X(n431)
         );
  SEN_AOI211_G_0P5 U585 ( .A1(N163), .A2(n382), .B1(n470), .B2(n469), .X(n472)
         );
  SEN_AOI211_G_0P5 U586 ( .A1(N167), .A2(n382), .B1(n498), .B2(n497), .X(n500)
         );
  SEN_INV_1 U587 ( .A(\sub_x_10_3/n88 ), .X(\sub_x_10_3/n87 ) );
  SEN_AOI211_G_0P5 U588 ( .A1(N165), .A2(n382), .B1(n484), .B2(n483), .X(n486)
         );
  SEN_AOI211_G_0P5 U589 ( .A1(N169), .A2(n382), .B1(n512), .B2(n511), .X(n514)
         );
  SEN_AOI211_G_0P5 U590 ( .A1(N160), .A2(n383), .B1(n449), .B2(n448), .X(n451)
         );
  SEN_AOI211_G_0P5 U591 ( .A1(N161), .A2(n383), .B1(n456), .B2(n455), .X(n458)
         );
  SEN_AOI21_T_1 U592 ( .A1(\cmp6_10_0/n33 ), .A2(n346), .B(n342), .X(
        \cmp6_10_0/n27 ) );
  SEN_MUXI2_D_1 U593 ( .D0(n598), .D1(n379), .S(\add_x_10_2/A[30] ), .X(n599)
         );
  SEN_MUXI2_S_0P5 U594 ( .D0(n496), .D1(n607), .S(\add_x_10_2/n70 ), .X(n497)
         );
  SEN_INV_1 U595 ( .A(\sub_x_10_3/n138 ), .X(\sub_x_10_3/n137 ) );
  SEN_OAOI211_1 U596 ( .A1(A[14]), .A2(n370), .B(n367), .C(n308), .X(n519) );
  SEN_OAOI211_1 U597 ( .A1(A[15]), .A2(n370), .B(n367), .C(n309), .X(n526) );
  SEN_MUXI2_S_0P5 U598 ( .D0(n510), .D1(n607), .S(\add_x_10_2/n60 ), .X(n511)
         );
  SEN_MUXI2_S_0P5 U599 ( .D0(n489), .D1(n607), .S(\add_x_10_2/n74 ), .X(n490)
         );
  SEN_MUXI2_S_0P5 U600 ( .D0(n503), .D1(n607), .S(\add_x_10_2/n64 ), .X(n504)
         );
  SEN_MUXI2_D_1 U601 ( .D0(n517), .D1(n381), .S(\add_x_10_2/n55 ), .X(n518) );
  SEN_MUXI2_D_1 U602 ( .D0(n595), .D1(n379), .S(\add_x_10_2/A[29] ), .X(n596)
         );
  SEN_MUXI2_D_1 U603 ( .D0(n524), .D1(n381), .S(\add_x_10_2/n51 ), .X(n525) );
  SEN_MUXI2_S_0P5 U604 ( .D0(n482), .D1(n607), .S(\add_x_10_2/n79 ), .X(n483)
         );
  SEN_INV_1 U605 ( .A(\add_x_10_1/n89 ), .X(\add_x_10_1/n88 ) );
  SEN_MUXI2_D_1 U606 ( .D0(n573), .D1(n381), .S(\add_x_10_2/A[22] ), .X(n574)
         );
  SEN_MUXI2_D_1 U607 ( .D0(n588), .D1(n381), .S(\add_x_10_2/n5 ), .X(n589) );
  SEN_MUXI2_D_1 U608 ( .D0(n538), .D1(n381), .S(\add_x_10_2/n40 ), .X(n539) );
  SEN_MUXI2_D_1 U609 ( .D0(n545), .D1(n381), .S(\add_x_10_2/n36 ), .X(n546) );
  SEN_AOI211_G_0P5 U610 ( .A1(B[0]), .A2(n420), .B1(n419), .B2(n418), .X(n421)
         );
  SEN_MUXI2_D_1 U611 ( .D0(n566), .D1(n381), .S(\add_x_10_2/A[21] ), .X(n567)
         );
  SEN_MUXI2_D_1 U612 ( .D0(n552), .D1(n381), .S(\add_x_10_2/n33 ), .X(n553) );
  SEN_MUXI2_S_0P5 U613 ( .D0(n424), .D1(n607), .S(\add_x_10_2/n111 ), .X(n428)
         );
  SEN_MUXI2_D_1 U614 ( .D0(n608), .D1(n379), .S(\add_x_10_2/A[31] ), .X(n609)
         );
  SEN_MUXI2_D_1 U615 ( .D0(n531), .D1(n381), .S(\add_x_10_2/n44 ), .X(n532) );
  SEN_MUXI2_D_1 U616 ( .D0(n580), .D1(n381), .S(\add_x_10_2/A[25] ), .X(n581)
         );
  SEN_MUXI2_D_1 U617 ( .D0(n559), .D1(n381), .S(\add_x_10_2/n27 ), .X(n560) );
  SEN_MUXI2_S_0P5 U618 ( .D0(n468), .D1(n607), .S(\add_x_10_2/n88 ), .X(n469)
         );
  SEN_AOI21_G_2 U619 ( .A1(\add_x_10_1/n64 ), .A2(n352), .B(\add_x_10_1/n61 ), 
        .X(\add_x_10_1/n59 ) );
  SEN_MUXI2_S_0P5 U620 ( .D0(n475), .D1(n607), .S(\add_x_10_2/n82 ), .X(n476)
         );
  SEN_INV_1 U621 ( .A(n368), .X(n366) );
  SEN_INV_1 U622 ( .A(\sub_x_10_3/n111 ), .X(\sub_x_10_3/n110 ) );
  SEN_MUXI2_S_0P5 U623 ( .D0(n454), .D1(n607), .S(\add_x_10_2/n95 ), .X(n455)
         );
  SEN_MUXI2_S_0P5 U624 ( .D0(n461), .D1(n607), .S(\add_x_10_2/n91 ), .X(n462)
         );
  SEN_MUXI2_S_0P5 U625 ( .D0(n440), .D1(n607), .S(\add_x_10_2/n104 ), .X(n441)
         );
  SEN_INV_1 U626 ( .A(\add_x_10_1/n139 ), .X(\add_x_10_1/n138 ) );
  SEN_INV_1 U627 ( .A(n368), .X(n367) );
  SEN_MUXI2_S_0P5 U628 ( .D0(n447), .D1(n607), .S(\add_x_10_2/n99 ), .X(n448)
         );
  SEN_MUXI2_S_0P5 U629 ( .D0(n433), .D1(n607), .S(\add_x_10_2/n107 ), .X(n434)
         );
  SEN_INV_1 U630 ( .A(\add_x_10_2/n67 ), .X(\add_x_10_2/n66 ) );
  SEN_AOI22_0P5 U631 ( .A1(A[0]), .A2(n383), .B1(n380), .B2(\add_x_10_2/n113 ), 
        .X(n416) );
  SEN_AOI21_G_1 U632 ( .A1(\sub_x_10_3/n161 ), .A2(\sub_x_10_3/n112 ), .B(
        \sub_x_10_3/n113 ), .X(\sub_x_10_3/n111 ) );
  SEN_INV_1 U633 ( .A(n603), .X(n368) );
  SEN_INV_1 U634 ( .A(\add_x_10_1/n112 ), .X(\add_x_10_1/n111 ) );
  SEN_INV_1 U635 ( .A(\sub_x_10_3/n161 ), .X(\sub_x_10_3/n160 ) );
  SEN_NR2_0P65 U636 ( .A1(n372), .A2(B[31]), .X(n605) );
  SEN_NR2_0P65 U637 ( .A1(n371), .A2(B[30]), .X(n597) );
  SEN_INV_1 U638 ( .A(\add_x_10_2/n47 ), .X(\add_x_10_2/n46 ) );
  SEN_OAI21_S_2 U639 ( .A1(\add_x_10_1/n112 ), .A2(\add_x_10_1/n65 ), .B(
        \add_x_10_1/n66 ), .X(\add_x_10_1/n64 ) );
  SEN_INV_1 U640 ( .A(n384), .X(n382) );
  SEN_NR2_G_1 U641 ( .A1(n426), .A2(n425), .X(n603) );
  SEN_INV_1 U642 ( .A(n362), .X(n373) );
  SEN_AOI21_T_1 U643 ( .A1(\add_x_10_1/n162 ), .A2(\add_x_10_1/n113 ), .B(
        \add_x_10_1/n114 ), .X(\add_x_10_1/n112 ) );
  SEN_INV_1 U644 ( .A(\add_x_10_2/n85 ), .X(\add_x_10_2/n84 ) );
  SEN_INV_S_0P5 U645 ( .A(n426), .X(n402) );
  SEN_INV_1 U646 ( .A(\sub_x_10_3/n182 ), .X(\sub_x_10_3/n181 ) );
  SEN_INV_1 U647 ( .A(n362), .X(n375) );
  SEN_INV_1 U648 ( .A(n362), .X(n374) );
  SEN_INV_1 U649 ( .A(n384), .X(n383) );
  SEN_INV_1 U650 ( .A(\add_x_10_1/n162 ), .X(\add_x_10_1/n161 ) );
  SEN_INV_1 U651 ( .A(\sub_x_10_3/n191 ), .X(\sub_x_10_3/n190 ) );
  SEN_NR2_S_0P5 U652 ( .A1(n604), .A2(B[2]), .X(n432) );
  SEN_INV_1 U653 ( .A(n380), .X(n381) );
  SEN_INV_1 U654 ( .A(n378), .X(n377) );
  SEN_NR2_S_0P5 U655 ( .A1(n604), .A2(B[3]), .X(n439) );
  SEN_NR2_G_1 U656 ( .A1(n397), .A2(n396), .X(n426) );
  SEN_INV_1 U657 ( .A(\add_x_10_2/n102 ), .X(\add_x_10_2/n101 ) );
  SEN_INV_1 U658 ( .A(n611), .X(n384) );
  SEN_INV_1 U659 ( .A(\add_x_10_1/n92 ), .X(\add_x_10_1/n90 ) );
  SEN_INV_1 U660 ( .A(\add_x_10_1/n183 ), .X(\add_x_10_1/n182 ) );
  SEN_INV_1 U661 ( .A(n378), .X(n376) );
  SEN_INV_1 U662 ( .A(\add_x_10_1/n93 ), .X(\add_x_10_1/n91 ) );
  SEN_INV_1 U663 ( .A(\add_x_10_1/n192 ), .X(\add_x_10_1/n191 ) );
  SEN_OAI21_G_1 U664 ( .A1(\cmp6_10_0/n68 ), .A2(\cmp6_10_0/n71 ), .B(
        \cmp6_10_0/n69 ), .X(\cmp6_10_0/n67 ) );
  SEN_INV_1 U665 ( .A(n612), .X(n387) );
  SEN_INV_1 U666 ( .A(\sub_x_10_3/n69 ), .X(\sub_x_10_3/n67 ) );
  SEN_NR2_G_1 U667 ( .A1(n406), .A2(n405), .X(n611) );
  SEN_INV_1 U668 ( .A(\sub_x_10_3/n136 ), .X(\sub_x_10_3/n134 ) );
  SEN_INV_1 U669 ( .A(\sub_x_10_3/n192 ), .X(\sub_x_10_3/n225 ) );
  SEN_INV_1 U670 ( .A(n606), .X(n378) );
  SEN_NR2_G_1 U671 ( .A1(n412), .A2(n395), .X(n396) );
  SEN_AOI21_G_1 U672 ( .A1(\add_x_10_1/n94 ), .A2(\add_x_10_1/n103 ), .B(
        \add_x_10_1/n95 ), .X(\add_x_10_1/n93 ) );
  SEN_INV_1 U673 ( .A(\sub_x_10_3/n82 ), .X(\sub_x_10_3/n205 ) );
  SEN_AOI22_0P5 U674 ( .A1(n606), .A2(A[0]), .B1(n425), .B2(n400), .X(n401) );
  SEN_INV_1 U675 ( .A(n607), .X(n380) );
  SEN_INV_1 U676 ( .A(\sub_x_10_3/n124 ), .X(\sub_x_10_3/n122 ) );
  SEN_INV_1 U677 ( .A(\sub_x_10_3/n135 ), .X(\sub_x_10_3/n214 ) );
  SEN_INV_1 U678 ( .A(\sub_x_10_3/n123 ), .X(\sub_x_10_3/n212 ) );
  SEN_INV_1 U679 ( .A(\sub_x_10_3/n78 ), .X(\sub_x_10_3/n76 ) );
  SEN_INV_1 U680 ( .A(n410), .X(n411) );
  SEN_INV_1 U681 ( .A(\add_x_10_1/n70 ), .X(\add_x_10_1/n68 ) );
  SEN_INV_1 U682 ( .A(\add_x_10_1/n79 ), .X(\add_x_10_1/n77 ) );
  SEN_NR2_G_1 U683 ( .A1(n406), .A2(n404), .X(n612) );
  SEN_INV_1 U684 ( .A(\add_x_10_1/n39 ), .X(\add_x_10_1/n37 ) );
  SEN_INV_1 U685 ( .A(\add_x_10_1/n47 ), .X(\add_x_10_1/n45 ) );
  SEN_OAI21_S_1 U686 ( .A1(n409), .A2(n410), .B(INST[1]), .X(n414) );
  SEN_INV_1 U687 ( .A(\add_x_10_1/n63 ), .X(\add_x_10_1/n61 ) );
  SEN_OAI21_S_1 U688 ( .A1(n409), .A2(n394), .B(INST[1]), .X(n397) );
  SEN_INV_1 U689 ( .A(n404), .X(n412) );
  SEN_INV_1 U690 ( .A(n602), .X(n365) );
  SEN_INV_1 U691 ( .A(\add_x_10_1/n136 ), .X(\add_x_10_1/n216 ) );
  SEN_INV_0P8 U692 ( .A(\add_x_10_1/n131 ), .X(\add_x_10_1/n215 ) );
  SEN_INV_1 U693 ( .A(\add_x_10_1/n137 ), .X(\add_x_10_1/n135 ) );
  SEN_AN2_1 U694 ( .A1(n348), .A2(\add_x_10_1/n196 ), .X(N124) );
  SEN_INV_1 U695 ( .A(\add_x_10_1/n124 ), .X(\add_x_10_1/n214 ) );
  SEN_INV_1 U696 ( .A(\add_x_10_1/n150 ), .X(\add_x_10_1/n148 ) );
  SEN_INV_1 U697 ( .A(\add_x_10_1/n125 ), .X(\add_x_10_1/n123 ) );
  SEN_INV_1 U698 ( .A(\add_x_10_1/n149 ), .X(\add_x_10_1/n218 ) );
  SEN_INV_1 U699 ( .A(\sub_x_10_3/n108 ), .X(\sub_x_10_3/n210 ) );
  SEN_INV_1 U700 ( .A(\sub_x_10_3/n109 ), .X(\sub_x_10_3/n107 ) );
  SEN_INV_1 U701 ( .A(\add_x_10_1/n193 ), .X(\add_x_10_1/n227 ) );
  SEN_INV_1 U702 ( .A(\sub_x_10_3/n188 ), .X(\sub_x_10_3/n224 ) );
  SEN_INV_1 U703 ( .A(\sub_x_10_3/n149 ), .X(\sub_x_10_3/n147 ) );
  SEN_INV_1 U704 ( .A(\add_x_10_1/n109 ), .X(\add_x_10_1/n212 ) );
  SEN_INV_1 U705 ( .A(\sub_x_10_3/n148 ), .X(\sub_x_10_3/n216 ) );
  SEN_INV_1 U706 ( .A(\add_x_10_1/n110 ), .X(\add_x_10_1/n108 ) );
  SEN_INV_1 U707 ( .A(\add_x_10_1/n189 ), .X(\add_x_10_1/n226 ) );
  SEN_INV_1 U708 ( .A(\add_x_10_1/n83 ), .X(\add_x_10_1/n207 ) );
  SEN_INV_1 U709 ( .A(\sub_x_10_3/n179 ), .X(\sub_x_10_3/n222 ) );
  SEN_INV_1 U710 ( .A(\sub_x_10_3/n180 ), .X(\sub_x_10_3/n178 ) );
  SEN_INV_1 U711 ( .A(\add_x_10_1/n180 ), .X(\add_x_10_1/n224 ) );
  SEN_INV_1 U712 ( .A(\add_x_10_1/n181 ), .X(\add_x_10_1/n179 ) );
  SEN_INV_1 U713 ( .A(A[29]), .X(\add_x_10_2/A[29] ) );
  SEN_INV_1 U714 ( .A(A[0]), .X(\add_x_10_2/n113 ) );
  SEN_INV_1 U715 ( .A(A[30]), .X(\add_x_10_2/A[30] ) );
  SEN_INV_1 U716 ( .A(n403), .X(n406) );
  SEN_NR2_G_1 U717 ( .A1(n399), .A2(n398), .X(n425) );
  SEN_INV_1 U718 ( .A(n394), .X(n395) );
  SEN_INV_1 U719 ( .A(A[28]), .X(\add_x_10_2/n5 ) );
  SEN_INV_1 U720 ( .A(A[26]), .X(\add_x_10_2/n10 ) );
  SEN_INV_1 U721 ( .A(A[25]), .X(\add_x_10_2/A[25] ) );
  SEN_INV_1 U722 ( .A(A[24]), .X(\add_x_10_2/n15 ) );
  SEN_INV_1 U723 ( .A(A[8]), .X(\add_x_10_2/n82 ) );
  SEN_INV_1 U724 ( .A(A[9]), .X(\add_x_10_2/n79 ) );
  SEN_INV_1 U725 ( .A(A[10]), .X(\add_x_10_2/n74 ) );
  SEN_INV_1 U726 ( .A(A[11]), .X(\add_x_10_2/n70 ) );
  SEN_INV_1 U727 ( .A(A[22]), .X(\add_x_10_2/A[22] ) );
  SEN_INV_1 U728 ( .A(A[12]), .X(\add_x_10_2/n64 ) );
  SEN_INV_1 U729 ( .A(A[21]), .X(\add_x_10_2/A[21] ) );
  SEN_INV_1 U730 ( .A(A[13]), .X(\add_x_10_2/n60 ) );
  SEN_INV_1 U731 ( .A(A[14]), .X(\add_x_10_2/n55 ) );
  SEN_INV_1 U732 ( .A(A[20]), .X(\add_x_10_2/n27 ) );
  SEN_INV_1 U733 ( .A(A[15]), .X(\add_x_10_2/n51 ) );
  SEN_INV_1 U734 ( .A(A[4]), .X(\add_x_10_2/n99 ) );
  SEN_NR2_G_1 U735 ( .A1(n408), .A2(INST[1]), .X(n407) );
  SEN_INV_1 U736 ( .A(A[5]), .X(\add_x_10_2/n95 ) );
  SEN_INV_1 U737 ( .A(A[19]), .X(\add_x_10_2/n33 ) );
  SEN_NR2_G_1 U738 ( .A1(n393), .A2(INST[3]), .X(n409) );
  SEN_INV_1 U739 ( .A(A[6]), .X(\add_x_10_2/n91 ) );
  SEN_INV_1 U740 ( .A(A[18]), .X(\add_x_10_2/n36 ) );
  SEN_INV_1 U741 ( .A(A[7]), .X(\add_x_10_2/n88 ) );
  SEN_INV_1 U742 ( .A(A[17]), .X(\add_x_10_2/n40 ) );
  SEN_INV_1 U743 ( .A(A[16]), .X(\add_x_10_2/n44 ) );
  SEN_INV_1 U744 ( .A(A[2]), .X(\add_x_10_2/n107 ) );
  SEN_INV_1 U745 ( .A(A[3]), .X(\add_x_10_2/n104 ) );
  SEN_INV_1 U746 ( .A(A[1]), .X(\add_x_10_2/n111 ) );
  SEN_INV_1 U747 ( .A(INST[3]), .X(n392) );
  SEN_INV_1 U748 ( .A(A[31]), .X(\add_x_10_2/A[31] ) );
  SEN_INV_1 U749 ( .A(INST[2]), .X(n408) );
  SEN_ND2_G_0P65 U750 ( .A1(INST[1]), .A2(INST[3]), .X(n398) );
  SEN_NR2_G_1 U751 ( .A1(INST[2]), .A2(INST[1]), .X(n403) );
  SEN_INV_1 U752 ( .A(INST[0]), .X(n393) );
  SEN_INV_S_0P5 U753 ( .A(SEL), .X(n400) );
  SEN_AN2_S_1 U754 ( .A1(n339), .A2(A[0]), .X(n343) );
  SEN_EO2_S_0P5 U755 ( .A1(A[26]), .A2(n333), .X(n346) );
  SEN_EO2_S_0P5 U756 ( .A1(A[28]), .A2(n334), .X(n345) );
  SEN_EO2_S_0P5 U757 ( .A1(A[30]), .A2(n335), .X(n344) );
  SEN_OR2_1 U758 ( .A1(A[31]), .A2(B[31]), .X(n347) );
  SEN_OR2_1 U759 ( .A1(A[0]), .A2(B[0]), .X(n348) );
  SEN_OR2_1 U760 ( .A1(A[30]), .A2(B[30]), .X(n349) );
  SEN_OR2_1 U761 ( .A1(A[28]), .A2(B[28]), .X(n350) );
  SEN_OR2_1 U762 ( .A1(A[26]), .A2(B[26]), .X(n351) );
  SEN_OR2_1 U763 ( .A1(A[24]), .A2(B[24]), .X(n352) );
  SEN_OR2_1 U764 ( .A1(A[23]), .A2(B[23]), .X(n353) );
  SEN_OR2_1 U765 ( .A1(A[22]), .A2(B[22]), .X(n354) );
  SEN_OAI21_S_2 U766 ( .A1(\add_x_10_1/n43 ), .A2(\add_x_10_1/n41 ), .B(
        \add_x_10_1/n42 ), .X(\add_x_10_1/n40 ) );
  SEN_EO2_1 U767 ( .A1(\add_x_10_1/n1 ), .A2(\add_x_10_1/n35 ), .X(N155) );
  SEN_OR2_1 U768 ( .A1(n331), .A2(A[31]), .X(n355) );
  SEN_OR2_1 U769 ( .A1(n335), .A2(A[30]), .X(n356) );
  SEN_OR2_1 U770 ( .A1(n334), .A2(A[28]), .X(n357) );
  SEN_OR2_1 U771 ( .A1(n333), .A2(A[26]), .X(n358) );
  SEN_OR2_1 U772 ( .A1(n336), .A2(A[24]), .X(n359) );
  SEN_OR2_1 U773 ( .A1(n319), .A2(A[23]), .X(n360) );
  SEN_OR2_1 U774 ( .A1(n320), .A2(A[22]), .X(n361) );
  SEN_OAI21_S_3 U775 ( .A1(\sub_x_10_3/n42 ), .A2(\sub_x_10_3/n40 ), .B(
        \sub_x_10_3/n41 ), .X(\sub_x_10_3/n39 ) );
  SEN_OAI21_S_2 U776 ( .A1(\sub_x_10_3/n50 ), .A2(\sub_x_10_3/n48 ), .B(
        \sub_x_10_3/n49 ), .X(\sub_x_10_3/n47 ) );
  SEN_AOI21_2 U777 ( .A1(N55), .A2(INST[1]), .B(INST[0]), .X(n388) );
  SEN_AOAI211_2 U778 ( .A1(n389), .A2(INST[0]), .B(n388), .C(n408), .X(n390)
         );
  SEN_MUXI2_DG_1 U779 ( .D0(N52), .D1(N53), .S(INST[1]), .X(n389) );
  SEN_ND3_1 U780 ( .A1(n391), .A2(INST[3]), .A3(n390), .X(n422) );
  SEN_OAOI211_G_1 U781 ( .A1(A[1]), .A2(n369), .B(n366), .C(n307), .X(n427) );
  SEN_OAOI211_G_1 U782 ( .A1(A[3]), .A2(n369), .B(n366), .C(n321), .X(n442) );
  SEN_OAOI211_G_1 U783 ( .A1(A[5]), .A2(n369), .B(n366), .C(n322), .X(n456) );
  SEN_OAOI211_G_1 U784 ( .A1(A[4]), .A2(n369), .B(n366), .C(n328), .X(n449) );
  SEN_OAOI211_G_1 U785 ( .A1(A[2]), .A2(n369), .B(n366), .C(n337), .X(n435) );
  SEN_OAOI211_G_1 U786 ( .A1(A[9]), .A2(n369), .B(n366), .C(n312), .X(n484) );
  SEN_OAOI211_G_1 U787 ( .A1(A[6]), .A2(n369), .B(n366), .C(n323), .X(n463) );
  SEN_OAOI211_G_1 U788 ( .A1(A[8]), .A2(n369), .B(n366), .C(n329), .X(n477) );
  SEN_OAOI211_G_1 U789 ( .A1(A[13]), .A2(n369), .B(n366), .C(n318), .X(n512)
         );
  SEN_OAOI211_G_1 U790 ( .A1(A[10]), .A2(n370), .B(n366), .C(n326), .X(n491)
         );
  SEN_OAOI211_G_1 U791 ( .A1(A[11]), .A2(n370), .B(n366), .C(n316), .X(n498)
         );
  SEN_OAOI211_G_1 U792 ( .A1(A[12]), .A2(n370), .B(n366), .C(n313), .X(n505)
         );
  SEN_ND2_G_1 U793 ( .A1(N152), .A2(n386), .X(n591) );
  SEN_ND2_G_1 U794 ( .A1(N376), .A2(n364), .X(n593) );
  SEN_OAOI211_G_1 U795 ( .A1(A[17]), .A2(n370), .B(n367), .C(n315), .X(n540)
         );
  SEN_OAOI211_G_1 U796 ( .A1(A[16]), .A2(n370), .B(n367), .C(n325), .X(n533)
         );
  SEN_OAOI211_G_1 U797 ( .A1(A[18]), .A2(n370), .B(n367), .C(n310), .X(n547)
         );
  SEN_OAOI211_G_1 U798 ( .A1(A[30]), .A2(n369), .B(n366), .C(n335), .X(n600)
         );
  SEN_OAOI211_G_1 U799 ( .A1(A[31]), .A2(n369), .B(n366), .C(n331), .X(n610)
         );
  SEN_ND2_G_1 U800 ( .A1(N379), .A2(n602), .X(n615) );
  SEN_ND2_G_1 U801 ( .A1(n422), .A2(n421), .X(Z[0]) );
  SEN_OAI211_1 U802 ( .A1(n417), .A2(B[0]), .B1(n416), .B2(n415), .X(n418) );
  SEN_ND2_G_1 U803 ( .A1(n375), .A2(A[0]), .X(n415) );
  SEN_NR2_1 U804 ( .A1(n412), .A2(n411), .X(n413) );
  SEN_NR2_1 U805 ( .A1(n408), .A2(SEL), .X(n410) );
  SEN_ND2_G_1 U806 ( .A1(n409), .A2(n407), .X(n607) );
  SEN_AO22_1 U807 ( .A1(n363), .A2(N348), .B1(N124), .B2(n385), .X(n419) );
  SEN_OAI211_1 U808 ( .A1(A[0]), .A2(n371), .B1(n402), .B2(n401), .X(n420) );
  SEN_ND2_G_1 U809 ( .A1(n407), .A2(n412), .X(n604) );
  SEN_ND2_G_1 U810 ( .A1(n393), .A2(n392), .X(n404) );
  SEN_AN3B_1 U811 ( .B1(n403), .B2(INST[3]), .A(INST[0]), .X(n602) );
  SEN_ND3_S_0P5 U812 ( .A1(n431), .A2(n430), .A3(n429), .X(Z[1]) );
  SEN_AOI211_0P5 U813 ( .A1(n606), .A2(B[1]), .B1(n375), .B2(n423), .X(n424)
         );
  SEN_ND3_S_0P5 U814 ( .A1(n445), .A2(n444), .A3(n443), .X(Z[3]) );
  SEN_AOI211_0P5 U815 ( .A1(n377), .A2(B[3]), .B1(n375), .B2(n439), .X(n440)
         );
  SEN_ND3_S_0P5 U816 ( .A1(n459), .A2(n458), .A3(n457), .X(Z[5]) );
  SEN_AOI211_0P5 U817 ( .A1(n377), .A2(B[5]), .B1(n375), .B2(n453), .X(n454)
         );
  SEN_ND3_S_0P5 U818 ( .A1(n452), .A2(n451), .A3(n450), .X(Z[4]) );
  SEN_AOI211_0P5 U819 ( .A1(n377), .A2(B[4]), .B1(n375), .B2(n446), .X(n447)
         );
  SEN_ND3_S_0P5 U820 ( .A1(n438), .A2(n437), .A3(n436), .X(Z[2]) );
  SEN_AOI211_0P5 U821 ( .A1(n376), .A2(B[2]), .B1(n375), .B2(n432), .X(n433)
         );
  SEN_ND3_S_0P5 U822 ( .A1(n487), .A2(n486), .A3(n485), .X(Z[9]) );
  SEN_AOI211_0P5 U823 ( .A1(n377), .A2(B[9]), .B1(n374), .B2(n481), .X(n482)
         );
  SEN_ND3_S_0P5 U824 ( .A1(n466), .A2(n465), .A3(n464), .X(Z[6]) );
  SEN_AOI211_0P5 U825 ( .A1(n377), .A2(B[6]), .B1(n374), .B2(n460), .X(n461)
         );
  SEN_ND3_S_0P5 U826 ( .A1(n473), .A2(n472), .A3(n471), .X(Z[7]) );
  SEN_AOI211_0P5 U827 ( .A1(n377), .A2(B[7]), .B1(n374), .B2(n467), .X(n468)
         );
  SEN_ND3_S_0P5 U828 ( .A1(n480), .A2(n479), .A3(n478), .X(Z[8]) );
  SEN_AOI211_0P5 U829 ( .A1(n377), .A2(B[8]), .B1(n374), .B2(n474), .X(n475)
         );
  SEN_ND3_S_0P5 U830 ( .A1(n515), .A2(n514), .A3(n513), .X(Z[13]) );
  SEN_AOI211_0P5 U831 ( .A1(n377), .A2(B[13]), .B1(n374), .B2(n509), .X(n510)
         );
  SEN_ND3_S_0P5 U832 ( .A1(n494), .A2(n493), .A3(n492), .X(Z[10]) );
  SEN_AOI211_0P5 U833 ( .A1(n377), .A2(B[10]), .B1(n374), .B2(n488), .X(n489)
         );
  SEN_ND3_S_0P5 U834 ( .A1(n501), .A2(n500), .A3(n499), .X(Z[11]) );
  SEN_AOI211_0P5 U835 ( .A1(n377), .A2(B[11]), .B1(n374), .B2(n495), .X(n496)
         );
  SEN_ND3_S_0P5 U836 ( .A1(n508), .A2(n507), .A3(n506), .X(Z[12]) );
  SEN_AOI211_0P5 U837 ( .A1(n377), .A2(B[12]), .B1(n374), .B2(n502), .X(n503)
         );
  SEN_ND3_S_0P5 U838 ( .A1(n593), .A2(n592), .A3(n591), .X(Z[28]) );
  SEN_AOI211_0P5 U839 ( .A1(N184), .A2(n611), .B1(n590), .B2(n589), .X(n592)
         );
  SEN_ND3_S_0P5 U840 ( .A1(n522), .A2(n521), .A3(n520), .X(Z[14]) );
  SEN_AOI211_0P5 U841 ( .A1(n377), .A2(B[14]), .B1(n374), .B2(n516), .X(n517)
         );
  SEN_ND3_S_0P5 U842 ( .A1(n543), .A2(n542), .A3(n541), .X(Z[17]) );
  SEN_AOI211_0P5 U843 ( .A1(n377), .A2(B[17]), .B1(n374), .B2(n537), .X(n538)
         );
  SEN_ND3_S_0P5 U844 ( .A1(n536), .A2(n535), .A3(n534), .X(Z[16]) );
  SEN_AOI211_0P5 U845 ( .A1(n377), .A2(B[16]), .B1(n374), .B2(n530), .X(n531)
         );
  SEN_ND3_S_0P5 U846 ( .A1(n585), .A2(n584), .A3(n583), .X(Z[25]) );
  SEN_AOI211_0P5 U847 ( .A1(n376), .A2(B[25]), .B1(n373), .B2(n579), .X(n580)
         );
  SEN_ND3_S_0P5 U848 ( .A1(n550), .A2(n549), .A3(n548), .X(Z[18]) );
  SEN_AOI211_0P5 U849 ( .A1(n376), .A2(B[18]), .B1(n374), .B2(n544), .X(n545)
         );
  SEN_ND3_S_0P5 U850 ( .A1(n529), .A2(n528), .A3(n527), .X(Z[15]) );
  SEN_AOI211_0P5 U851 ( .A1(N171), .A2(n382), .B1(n526), .B2(n525), .X(n528)
         );
  SEN_AOI211_0P5 U852 ( .A1(n377), .A2(B[15]), .B1(n374), .B2(n523), .X(n524)
         );
  SEN_ND3_S_0P5 U853 ( .A1(n571), .A2(n570), .A3(n569), .X(Z[21]) );
  SEN_AOI211_0P5 U854 ( .A1(N177), .A2(n382), .B1(n568), .B2(n567), .X(n570)
         );
  SEN_AOI211_0P5 U855 ( .A1(n376), .A2(B[21]), .B1(n373), .B2(n565), .X(n566)
         );
  SEN_ND3_S_0P5 U856 ( .A1(n557), .A2(n556), .A3(n555), .X(Z[19]) );
  SEN_AOI211_0P5 U857 ( .A1(N175), .A2(n383), .B1(n554), .B2(n553), .X(n556)
         );
  SEN_AOI211_0P5 U858 ( .A1(n376), .A2(B[19]), .B1(n373), .B2(n551), .X(n552)
         );
  SEN_ND3_S_0P5 U859 ( .A1(n564), .A2(n563), .A3(n562), .X(Z[20]) );
  SEN_AOI211_0P5 U860 ( .A1(n376), .A2(B[20]), .B1(n373), .B2(n558), .X(n559)
         );
  SEN_ND3_S_0P5 U861 ( .A1(n578), .A2(n577), .A3(n576), .X(Z[22]) );
  SEN_AOI211_0P5 U862 ( .A1(n376), .A2(B[22]), .B1(n373), .B2(n572), .X(n573)
         );
  SEN_AOI211_0P5 U863 ( .A1(B[31]), .A2(n376), .B1(n373), .B2(n605), .X(n608)
         );
  SEN_OR2_1 U864 ( .A1(n414), .A2(n413), .X(n362) );
endmodule

