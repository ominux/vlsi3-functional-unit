
module Alu ( Z, A, B, INST, SEL );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  input SEL;
  wire   n216, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n288, n289, n290, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n370, n373, n374, n375, n376,
         n377, n378, n379, n380, n383, n384, n385, n386, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;

  SEN_ND2_4 U265 ( .A1(n1288), .A2(n272), .X(n1290) );
  SEN_AOI21B_3 U266 ( .A1(n1275), .A2(n1276), .B(n306), .X(n1288) );
  SEN_INV_1P5 U267 ( .A(n1287), .X(n1292) );
  SEN_INV_0P8 U268 ( .A(n256), .X(n1248) );
  SEN_ND3_T_0P8 U269 ( .A1(n1258), .A2(n1257), .A3(n1256), .X(Z[30]) );
  SEN_NR2_T_1 U272 ( .A1(n925), .A2(n924), .X(n929) );
  SEN_MUXI2_DG_1 U277 ( .D0(n1223), .D1(n1217), .S(A[29]), .X(n1228) );
  SEN_INV_2 U279 ( .A(n1152), .X(n1186) );
  SEN_ND2_G_1 U280 ( .A1(n373), .A2(n1214), .X(n1215) );
  SEN_ND2_T_0P5 U281 ( .A1(n343), .A2(n1076), .X(n1082) );
  SEN_AOI21B_0P5 U282 ( .A1(n272), .A2(n344), .B(n375), .X(n697) );
  SEN_OR2_1 U283 ( .A1(B[13]), .A2(A[13]), .X(n855) );
  SEN_ND3_T_1P5 U284 ( .A1(n437), .A2(n436), .A3(n435), .X(n500) );
  SEN_ND2_T_2 U290 ( .A1(n1299), .A2(n319), .X(n320) );
  SEN_INV_1P25 U291 ( .A(n235), .X(n289) );
  SEN_MUXI2_DG_3 U294 ( .D0(n1134), .D1(n1139), .S(B[25]), .X(n1135) );
  SEN_ND2B_S_0P5 U295 ( .A(n380), .B(n869), .X(n867) );
  SEN_OAI21_G_0P5 U296 ( .A1(n866), .A2(n891), .B(n959), .X(n869) );
  SEN_OAI211_4 U299 ( .A1(n1292), .A2(n379), .B1(n1290), .B2(n375), .X(n1299)
         );
  SEN_ND2_1P5 U302 ( .A1(n531), .A2(n458), .X(n620) );
  SEN_ND2B_V1_1 U305 ( .A(B[13]), .B(A[13]), .X(n865) );
  SEN_INV_S_3 U307 ( .A(n627), .X(n659) );
  SEN_OAI211_0P5 U312 ( .A1(n271), .A2(n868), .B1(n375), .B2(n867), .X(n873)
         );
  SEN_ND2_T_0P5 U314 ( .A1(n1046), .A2(n339), .X(n1015) );
  SEN_INV_1P5 U316 ( .A(n563), .X(n462) );
  SEN_OR3B_2 U317 ( .B1(A[7]), .B2(A[8]), .A(n691), .X(n701) );
  SEN_INV_S_4 U318 ( .A(n660), .X(n691) );
  SEN_ND2_2 U319 ( .A1(n758), .A2(n674), .X(n732) );
  SEN_MUXI2_S_1 U321 ( .D0(n1174), .D1(n1178), .S(B[27]), .X(n1175) );
  SEN_ND2_T_1 U322 ( .A1(n1169), .A2(n1168), .X(n1174) );
  SEN_ND2B_2 U323 ( .A(n703), .B(n702), .X(n704) );
  SEN_MUXI2_DG_2 U324 ( .D0(n700), .D1(n296), .S(B[9]), .X(n703) );
  SEN_INV_S_4 U325 ( .A(n902), .X(n949) );
  SEN_OR3B_4 U326 ( .B1(A[15]), .B2(A[16]), .A(n896), .X(n902) );
  SEN_AO2BB2_4 U327 ( .A1(B[18]), .A2(A[18]), .B1(n957), .B2(n1007), .X(n1000)
         );
  SEN_OAI21_T_0P5 U331 ( .A1(n1218), .A2(n385), .B(n1219), .X(n1197) );
  SEN_ND2_2 U332 ( .A1(n1179), .A2(n238), .X(n1180) );
  SEN_MUXI2_DG_3 U334 ( .D0(n1225), .D1(n1224), .S(A[29]), .X(n1226) );
  SEN_NR2_G_2 U336 ( .A1(n1138), .A2(n298), .X(n1141) );
  SEN_ND2_S_1 U337 ( .A1(n389), .A2(n1218), .X(n1200) );
  SEN_OR3B_1 U338 ( .B1(n298), .B2(n1253), .A(n1301), .X(n1255) );
  SEN_ND2B_V1_4 U339 ( .A(A[29]), .B(n1252), .X(n1301) );
  SEN_MUXI2_DG_1 U340 ( .D0(n1159), .D1(n1158), .S(A[26]), .X(n1160) );
  SEN_INV_S_6 U341 ( .A(n1222), .X(n1252) );
  SEN_INV_S_1 U343 ( .A(n1157), .X(n1138) );
  SEN_ND2B_S_8 U344 ( .A(n1221), .B(n388), .X(n1222) );
  SEN_OR3B_4 U345 ( .B1(A[27]), .B2(n268), .A(n1218), .X(n1221) );
  SEN_INV_S_2 U346 ( .A(n1197), .X(n1176) );
  SEN_ND2_T_2 U347 ( .A1(n1285), .A2(n1239), .X(n1191) );
  SEN_INV_0P65 U351 ( .A(n607), .X(n605) );
  SEN_OR3B_1 U354 ( .B1(A[21]), .B2(A[22]), .A(n1071), .X(n1072) );
  SEN_OAI211_3 U358 ( .A1(n324), .A2(n370), .B1(n375), .B2(n1133), .X(n1139)
         );
  SEN_AN2_S_2 U364 ( .A1(n1283), .A2(n415), .X(n345) );
  SEN_ND2_G_1 U365 ( .A1(n731), .A2(n730), .X(n759) );
  SEN_ND2_T_1 U366 ( .A1(n715), .A2(n714), .X(n730) );
  SEN_ND2_T_0P5 U367 ( .A1(n883), .A2(n885), .X(n954) );
  SEN_NR2B_V1DG_3 U369 ( .A(n1006), .B(n311), .X(n312) );
  SEN_ND2_T_2 U371 ( .A1(n1129), .A2(n1128), .X(n1132) );
  SEN_ND3_S_0P5 U372 ( .A1(n270), .A2(n378), .A3(n374), .X(n518) );
  SEN_NR2_T_1 U374 ( .A1(n606), .A2(n605), .X(n612) );
  SEN_ND3_T_2 U378 ( .A1(n316), .A2(n317), .A3(n374), .X(n846) );
  SEN_AO21B_1 U380 ( .A1(n1043), .A2(n1015), .B(n1045), .X(n1026) );
  SEN_INV_S_2 U388 ( .A(A[28]), .X(n267) );
  SEN_OAI211_3 U391 ( .A1(n1301), .A2(A[30]), .B1(n279), .B2(n299), .X(n1302)
         );
  SEN_MUXI2_DG_0P75 U394 ( .D0(n1037), .D1(n1029), .S(B[21]), .X(n1030) );
  SEN_AN2_S_0P5 U397 ( .A1(B[9]), .A2(A[9]), .X(n235) );
  SEN_OA21B_0P5 U398 ( .A1(n1071), .A2(n385), .B(n355), .X(n236) );
  SEN_INV_S_0P5 U399 ( .A(n865), .X(n293) );
  SEN_ND2_S_0P5 U400 ( .A1(n843), .A2(n272), .X(n237) );
  SEN_AN2_S_1 U401 ( .A1(n330), .A2(n331), .X(n238) );
  SEN_AN2_S_1 U402 ( .A1(n1011), .A2(n1010), .X(n239) );
  SEN_INV_S_2 U403 ( .A(n1190), .X(n1193) );
  SEN_ND3_T_0P8 U404 ( .A1(n1205), .A2(n1204), .A3(n1203), .X(Z[28]) );
  SEN_INV_S_0P5 U406 ( .A(n969), .X(n966) );
  SEN_ND2_S_3 U408 ( .A1(n623), .A2(n459), .X(n328) );
  SEN_INV_3 U411 ( .A(n740), .X(n738) );
  SEN_AOAI211_G_0P5 U412 ( .A1(n860), .A2(n815), .B(n293), .C(n861), .X(n837)
         );
  SEN_ND2_0P8 U413 ( .A1(n345), .A2(n419), .X(n427) );
  SEN_AOI211_G_2 U414 ( .A1(n434), .A2(n433), .B1(n432), .B2(n498), .X(n435)
         );
  SEN_MUXI2_S_1 U420 ( .D0(n1249), .D1(n1248), .S(n1247), .X(n1258) );
  SEN_ND2B_2 U426 ( .A(n915), .B(n952), .X(n918) );
  SEN_AOI211_G_1 U428 ( .A1(n1040), .A2(n1042), .B1(n431), .B2(n430), .X(n432)
         );
  SEN_ND2_2 U429 ( .A1(n427), .A2(n497), .X(n431) );
  SEN_AO21_2 U430 ( .A1(n731), .A2(n353), .B(n733), .X(n765) );
  SEN_OR3B_2 U431 ( .B1(n241), .B2(A[0]), .A(n560), .X(n561) );
  SEN_INV_S_2 U432 ( .A(A[1]), .X(n560) );
  SEN_INV_S_4 U433 ( .A(n240), .X(n241) );
  SEN_ND2_S_4 U434 ( .A1(n771), .A2(n770), .X(n740) );
  SEN_ND2_4 U435 ( .A1(n734), .A2(n289), .X(n771) );
  SEN_NR2_T_1P5 U436 ( .A1(n1214), .A2(n271), .X(n333) );
  SEN_AOAI211_G_2 U442 ( .A1(n1265), .A2(n1266), .B(n1263), .C(n1267), .X(
        n1173) );
  SEN_NR2B_V1DG_1 U450 ( .A(n715), .B(n719), .X(n402) );
  SEN_INV_S_1P5 U453 ( .A(n1294), .X(n1295) );
  SEN_ND2_S_3 U454 ( .A1(n283), .A2(n1250), .X(n1294) );
  SEN_ND3_S_2 U455 ( .A1(n313), .A2(n314), .A3(n374), .X(n904) );
  SEN_MUXI2_DG_1 U458 ( .D0(n1196), .D1(n1195), .S(n1194), .X(n1205) );
  SEN_AOI21B_1 U460 ( .A1(n1119), .A2(n1116), .B(n1115), .X(n1129) );
  SEN_ND2_T_1 U461 ( .A1(n874), .A2(n845), .X(n849) );
  SEN_AOAI211_0P75 U467 ( .A1(n403), .A2(n402), .B(n401), .C(n400), .X(n406)
         );
  SEN_ND2_S_1 U471 ( .A1(n989), .A2(n304), .X(n961) );
  SEN_ND2_0P8 U474 ( .A1(B[3]), .A2(A[3]), .X(n607) );
  SEN_OR3B_2 U476 ( .B1(A[19]), .B2(A[20]), .A(n1023), .X(n1032) );
  SEN_ND2_T_1P5 U479 ( .A1(n1176), .A2(n1175), .X(n1181) );
  SEN_OR3B_1 U480 ( .B1(n249), .B2(n298), .A(n847), .X(n848) );
  SEN_MUXI2_S_1 U481 ( .D0(n846), .D1(n1298), .S(B[15]), .X(n847) );
  SEN_INV_3 U482 ( .A(A[2]), .X(n240) );
  SEN_MUXI2_D_1 U486 ( .D0(n514), .D1(n522), .S(n503), .X(n506) );
  SEN_MUXI2_S_2 U487 ( .D0(n1139), .D1(n1298), .S(B[25]), .X(n1140) );
  SEN_ND2_T_1 U490 ( .A1(n1080), .A2(n1079), .X(n1081) );
  SEN_MUXI2_S_1 U492 ( .D0(n1075), .D1(n1078), .S(B[23]), .X(n1076) );
  SEN_AN2_S_4 U493 ( .A1(n320), .A2(n321), .X(n279) );
  SEN_AOAI211_1 U494 ( .A1(n354), .A2(n1145), .B(n1146), .C(n1144), .X(Z[25])
         );
  SEN_ND2_0P5 U495 ( .A1(B[15]), .A2(A[15]), .X(n952) );
  SEN_AO21B_2 U498 ( .A1(n617), .A2(n616), .B(n615), .X(n619) );
  SEN_ND2_2 U499 ( .A1(n266), .A2(n732), .X(n677) );
  SEN_OR4B_4 U501 ( .B1(n1127), .B2(n1126), .B3(n1125), .A(n1124), .X(n1128)
         );
  SEN_AO21B_4 U506 ( .A1(n775), .A2(n332), .B(n774), .X(n780) );
  SEN_AN2_2 U507 ( .A1(n777), .A2(n778), .X(n332) );
  SEN_AN2_S_1 U508 ( .A1(n988), .A2(n994), .X(n304) );
  SEN_ND2B_S_0P5 U509 ( .A(B[27]), .B(A[27]), .X(n1239) );
  SEN_INV_S_2 U514 ( .A(n1147), .X(n324) );
  SEN_OR2_DG_1 U517 ( .A1(n841), .A2(n377), .X(n310) );
  SEN_NR2_G_0P5 U518 ( .A1(n438), .A2(n719), .X(n442) );
  SEN_NR2B_V1_1 U520 ( .A(n266), .B(n453), .X(n457) );
  SEN_AN3B_0P5 U521 ( .B1(n865), .B2(n988), .A(n454), .X(n455) );
  SEN_AOAI211_0P5 U522 ( .A1(n395), .A2(n394), .B(n393), .C(n392), .X(n399) );
  SEN_ND2_T_1 U523 ( .A1(n861), .A2(n860), .X(n863) );
  SEN_ND2B_S_0P5 U524 ( .A(B[1]), .B(A[1]), .X(n590) );
  SEN_ND2B_S_0P5 U526 ( .A(B[4]), .B(A[4]), .X(n618) );
  SEN_ND2_T_1 U527 ( .A1(n586), .A2(n585), .X(n606) );
  SEN_ND2B_1 U529 ( .A(A[8]), .B(B[8]), .X(n714) );
  SEN_NR2_S_0P5 U530 ( .A1(A[9]), .A2(B[9]), .X(n337) );
  SEN_INV_S_1P5 U531 ( .A(n711), .X(n338) );
  SEN_ND2B_V1DG_1 U533 ( .A(n889), .B(n304), .X(n923) );
  SEN_ND2B_V1DG_1 U534 ( .A(B[15]), .B(A[15]), .X(n959) );
  SEN_INV_0P65 U535 ( .A(n274), .X(n294) );
  SEN_ND3_T_2 U536 ( .A1(n1009), .A2(n278), .A3(n239), .X(n1012) );
  SEN_OR3B_2 U538 ( .B1(A[23]), .B2(A[24]), .A(n1131), .X(n1137) );
  SEN_ND2B_S_0P5 U539 ( .A(A[0]), .B(B[0]), .X(n531) );
  SEN_AOAI211_0P75 U542 ( .A1(n835), .A2(n274), .B(n834), .C(n290), .X(n843)
         );
  SEN_NR2_G_0P8 U543 ( .A1(n961), .A2(n890), .X(n838) );
  SEN_NR2_1 U544 ( .A1(n913), .A2(n911), .X(n888) );
  SEN_INV_S_0P5 U545 ( .A(n1015), .X(n1024) );
  SEN_OAI21_0P75 U546 ( .A1(n1070), .A2(n1069), .B(n346), .X(n1074) );
  SEN_INV_2 U547 ( .A(n1132), .X(n1150) );
  SEN_MUXI2_S_0P5 U551 ( .D0(n747), .D1(n749), .S(B[11]), .X(n748) );
  SEN_MUXI2_S_0P5 U552 ( .D0(n749), .D1(n1298), .S(B[11]), .X(n750) );
  SEN_ND2_0P8 U555 ( .A1(n971), .A2(n970), .X(n977) );
  SEN_ND2B_S_1 U556 ( .A(n1034), .B(n1033), .X(n1035) );
  SEN_MUXI2_DG_0P75 U557 ( .D0(n1031), .D1(n296), .S(B[21]), .X(n1034) );
  SEN_ND2_S_2 U559 ( .A1(n336), .A2(n1215), .X(n1217) );
  SEN_OA2BB2_0P5 U560 ( .A1(n1244), .A2(n373), .B1(n377), .B2(n1245), .X(n256)
         );
  SEN_OAI21_0P75 U561 ( .A1(n529), .A2(n528), .B(n527), .X(Z[0]) );
  SEN_ND2_S_0P5 U562 ( .A1(n860), .A2(n815), .X(n242) );
  SEN_ND2_S_0P5 U563 ( .A1(n853), .A2(n852), .X(n914) );
  SEN_INV_S_0P5 U564 ( .A(B[15]), .X(n853) );
  SEN_OAI22_S_0P5 U565 ( .A1(B[15]), .A2(A[15]), .B1(A[16]), .B2(B[16]), .X(
        n253) );
  SEN_AN3B_0P5 U566 ( .B1(n989), .B2(n988), .A(n990), .X(n997) );
  SEN_ND2_S_0P5 U567 ( .A1(n604), .A2(n389), .X(n580) );
  SEN_OAI22_S_0P5 U568 ( .A1(n642), .A2(n271), .B1(n377), .B2(n1312), .X(n645)
         );
  SEN_ND2_S_0P5 U569 ( .A1(n1304), .A2(B[8]), .X(n689) );
  SEN_INV_S_0P5 U570 ( .A(n242), .X(n444) );
  SEN_OA21B_0P5 U571 ( .A1(n795), .A2(n385), .B(n355), .X(n786) );
  SEN_ND2_S_0P5 U572 ( .A1(n682), .A2(n683), .X(n687) );
  SEN_OAI22_S_0P5 U573 ( .A1(n271), .A2(n870), .B1(n378), .B2(n869), .X(n872)
         );
  SEN_OAI211_0P5 U574 ( .A1(n735), .A2(n354), .B1(n729), .B2(n728), .X(Z[10])
         );
  SEN_OA21B_0P5 U575 ( .A1(n839), .A2(n385), .B(n355), .X(n824) );
  SEN_ND2_S_0P5 U576 ( .A1(n725), .A2(n1300), .X(n243) );
  SEN_INV_S_0P5 U577 ( .A(n243), .X(n702) );
  SEN_OA2BB2_1 U578 ( .A1(n1026), .A2(n373), .B1(n377), .B2(n1028), .X(n244)
         );
  SEN_INV_S_0P5 U579 ( .A(n244), .X(n1037) );
  SEN_ND2_S_0P5 U580 ( .A1(n297), .A2(B[12]), .X(n793) );
  SEN_ND2B_S_0P5 U581 ( .A(A[15]), .B(B[15]), .X(n926) );
  SEN_NR2_S_0P5 U582 ( .A1(A[20]), .A2(B[20]), .X(n245) );
  SEN_INV_S_0P5 U583 ( .A(n245), .X(n1043) );
  SEN_OA21B_0P5 U584 ( .A1(n896), .A2(n385), .B(n355), .X(n874) );
  SEN_NR2B_V1_1 U586 ( .A(n580), .B(n298), .X(n571) );
  SEN_OAI21_S_0P5 U587 ( .A1(n378), .A2(n744), .B(n741), .X(n747) );
  SEN_ND2_S_0P5 U588 ( .A1(n786), .A2(n787), .X(n791) );
  SEN_OAI211_0P5 U589 ( .A1(n271), .A2(n937), .B1(n375), .B2(n936), .X(n939)
         );
  SEN_OAI211_0P5 U590 ( .A1(n832), .A2(n354), .B1(n830), .B2(n829), .X(Z[14])
         );
  SEN_ND2_S_0P5 U591 ( .A1(n761), .A2(n757), .X(n440) );
  SEN_ND2B_S_0P5 U592 ( .A(B[21]), .B(A[21]), .X(n1040) );
  SEN_NR2_S_0P5 U593 ( .A1(A[22]), .A2(B[22]), .X(n246) );
  SEN_INV_S_0P5 U594 ( .A(n246), .X(n1064) );
  SEN_OA21B_0P5 U595 ( .A1(n604), .A2(n386), .B(n355), .X(n578) );
  SEN_AN2_S_0P5 U596 ( .A1(n389), .A2(n795), .X(n247) );
  SEN_INV_0P5 U597 ( .A(n247), .X(n789) );
  SEN_NR2B_V1_1 U598 ( .A(n826), .B(n298), .X(n806) );
  SEN_OA2BB2_0P5 U599 ( .A1(n373), .A2(n937), .B1(n378), .B2(n935), .X(n248)
         );
  SEN_INV_S_0P5 U600 ( .A(n248), .X(n940) );
  SEN_OAI211_0P5 U601 ( .A1(n271), .A2(n1152), .B1(n375), .B2(n1151), .X(n1155) );
  SEN_ND2B_S_0P5 U602 ( .A(n315), .B(n765), .X(n767) );
  SEN_ND2B_S_0P5 U603 ( .A(B[19]), .B(A[19]), .X(n1041) );
  SEN_OAI21_S_0P5 U604 ( .A1(A[21]), .A2(B[21]), .B(n1043), .X(n1061) );
  SEN_ND2_S_0P5 U605 ( .A1(n824), .A2(n825), .X(n828) );
  SEN_MUXI2_S_0P5 U606 ( .D0(n872), .D1(n873), .S(n871), .X(n882) );
  SEN_NR2B_V1_1 U607 ( .A(n926), .B(n871), .X(n422) );
  SEN_AN2_S_0P5 U608 ( .A1(n389), .A2(n896), .X(n249) );
  SEN_INV_0P5 U609 ( .A(n249), .X(n877) );
  SEN_NR2B_V1_1 U610 ( .A(n1055), .B(n298), .X(n1033) );
  SEN_OAI22_S_0P5 U611 ( .A1(n370), .A2(n284), .B1(n377), .B2(n1074), .X(n1075) );
  SEN_AN3B_0P5 U613 ( .B1(n988), .B2(n994), .A(n890), .X(n816) );
  SEN_ND2_S_0P5 U614 ( .A1(B[21]), .A2(A[21]), .X(n1044) );
  SEN_ND2_S_0P5 U615 ( .A1(n874), .A2(n875), .X(n879) );
  SEN_ND2_S_0P5 U616 ( .A1(n901), .A2(n900), .X(n907) );
  SEN_MUXI2_S_0P5 U617 ( .D0(n1018), .D1(n1019), .S(n472), .X(n1021) );
  SEN_ND4_S_0P5 U618 ( .A1(n407), .A2(n993), .A3(n964), .A4(n930), .X(n300) );
  SEN_ND2_S_0P5 U619 ( .A1(A[12]), .A2(B[12]), .X(n885) );
  SEN_NR2_S_0P5 U620 ( .A1(B[25]), .A2(A[25]), .X(n250) );
  SEN_INV_S_0P5 U621 ( .A(n250), .X(n1234) );
  SEN_NR3_0P5 U622 ( .A1(n890), .A2(n961), .A3(n990), .X(n866) );
  SEN_INV_S_0P5 U623 ( .A(n995), .X(n890) );
  SEN_AN2_S_0P5 U624 ( .A1(n389), .A2(n1023), .X(n251) );
  SEN_INV_0P5 U625 ( .A(n251), .X(n984) );
  SEN_ND2_S_0P5 U627 ( .A1(n295), .A2(B[4]), .X(n581) );
  SEN_OA21B_0P5 U628 ( .A1(n742), .A2(n385), .B(n355), .X(n723) );
  SEN_OAI22_S_0P5 U629 ( .A1(n1186), .A2(n271), .B1(n378), .B2(n1163), .X(
        n1154) );
  SEN_NR2_S_0P5 U631 ( .A1(n293), .A2(n454), .X(n443) );
  SEN_ND2_S_0P5 U632 ( .A1(n1188), .A2(n487), .X(n252) );
  SEN_INV_S_0P5 U633 ( .A(n252), .X(n488) );
  SEN_INV_S_0P5 U634 ( .A(n253), .X(n919) );
  SEN_OA21B_0P5 U635 ( .A1(n659), .A2(n386), .B(n355), .X(n647) );
  SEN_NR2B_V1_1 U636 ( .A(n984), .B(n298), .X(n974) );
  SEN_NR2B_2 U637 ( .A(n1216), .B(n380), .X(n335) );
  SEN_MUXI2_S_0P5 U638 ( .D0(n1052), .D1(n1053), .S(n424), .X(n1059) );
  SEN_ND2_S_0P5 U639 ( .A1(n764), .A2(n266), .X(n254) );
  SEN_INV_S_0P5 U640 ( .A(n254), .X(n398) );
  SEN_INV_S_0P5 U641 ( .A(n265), .X(n266) );
  SEN_ND2B_S_0P5 U643 ( .A(A[16]), .B(B[16]), .X(n927) );
  SEN_NR2_S_0P5 U644 ( .A1(A[17]), .A2(B[17]), .X(n255) );
  SEN_INV_S_0P5 U645 ( .A(n255), .X(n916) );
  SEN_ND2_S_0P5 U646 ( .A1(B[19]), .A2(A[19]), .X(n1046) );
  SEN_NR2B_V1_1 U647 ( .A(n1239), .B(n492), .X(n495) );
  SEN_ND4_S_0P5 U648 ( .A1(n933), .A2(n960), .A3(n959), .A4(n995), .X(n962) );
  SEN_MUX2_S_0P5 U649 ( .D0(n570), .D1(n295), .S(B[3]), .X(n572) );
  SEN_ND2_S_0P5 U650 ( .A1(n901), .A2(n942), .X(n946) );
  SEN_MUXI2_S_0P5 U651 ( .D0(n1109), .D1(n1110), .S(n482), .X(n1112) );
  SEN_NR2B_V1_1 U652 ( .A(A[7]), .B(B[7]), .X(n265) );
  SEN_NR2B_V1_1 U653 ( .A(B[31]), .B(A[31]), .X(n498) );
  SEN_ND2B_S_0P5 U655 ( .A(A[17]), .B(B[17]), .X(n930) );
  SEN_NR2_S_0P5 U656 ( .A1(B[19]), .A2(A[19]), .X(n999) );
  SEN_OA21_1 U657 ( .A1(n342), .A2(n1068), .B(n1067), .X(n346) );
  SEN_AOI21_S_0P5 U658 ( .A1(A[26]), .A2(B[26]), .B(n1166), .X(n318) );
  SEN_AOAI211_0P5 U659 ( .A1(n1281), .A2(n1282), .B(n1286), .C(n1283), .X(n259) );
  SEN_OA2BB2_0P5 U660 ( .A1(n373), .A2(n796), .B1(n377), .B2(n781), .X(n257)
         );
  SEN_INV_S_0P5 U661 ( .A(n257), .X(n784) );
  SEN_ND2_S_0P5 U662 ( .A1(n1304), .A2(B[26]), .X(n1161) );
  SEN_ND2_S_0P5 U663 ( .A1(n770), .A2(n772), .X(n258) );
  SEN_INV_S_0P5 U664 ( .A(n258), .X(n275) );
  SEN_ND2_S_0P5 U665 ( .A1(n1118), .A2(n1119), .X(n1127) );
  SEN_ND2_S_0P5 U667 ( .A1(n290), .A2(n952), .X(n911) );
  SEN_INV_0P8 U668 ( .A(n269), .X(n290) );
  SEN_ND2B_S_0P5 U669 ( .A(B[17]), .B(A[17]), .X(n933) );
  SEN_ND2_S_0P5 U670 ( .A1(A[18]), .A2(B[18]), .X(n1006) );
  SEN_AOI31_0P5 U672 ( .A1(n1260), .A2(n1235), .A3(n1232), .B(n1268), .X(n1238) );
  SEN_INV_S_0P5 U673 ( .A(n259), .X(n1284) );
  SEN_ND3_S_0P5 U674 ( .A1(n374), .A2(n1048), .A3(n1047), .X(n1053) );
  SEN_OA21B_0P5 U675 ( .A1(n1131), .A2(n385), .B(n355), .X(n343) );
  SEN_ND2_S_0P5 U677 ( .A1(n1136), .A2(n1156), .X(n1159) );
  SEN_AN3B_2 U678 ( .B1(n348), .B2(n1222), .A(n298), .X(n281) );
  SEN_ND2_S_0P5 U679 ( .A1(n1304), .A2(B[28]), .X(n1204) );
  SEN_ND2_S_0P5 U680 ( .A1(B[17]), .A2(A[17]), .X(n1007) );
  SEN_ND2_S_0P5 U681 ( .A1(n862), .A2(n861), .X(n454) );
  SEN_AO2BB2_0P5 U682 ( .A1(A[16]), .A2(B[16]), .B1(n886), .B2(n952), .X(n887)
         );
  SEN_OR4B_1 U683 ( .B1(n1099), .B2(n1098), .B3(n1100), .A(n1124), .X(n1101)
         );
  SEN_AOI21B_2 U684 ( .A1(n1265), .A2(n318), .B(n1270), .X(n1275) );
  SEN_ND2_S_0P5 U685 ( .A1(n503), .A2(INST[1]), .X(n502) );
  SEN_OAI221_0P5 U686 ( .A1(n1055), .A2(A[21]), .B1(n296), .B2(n1060), .C(
        n1300), .X(n1056) );
  SEN_ND2B_S_0P5 U687 ( .A(n385), .B(A[23]), .X(n1085) );
  SEN_ND2_S_0P5 U688 ( .A1(n1298), .A2(B[28]), .X(n1199) );
  SEN_OR2_DG_1 U689 ( .A1(n1216), .A2(n378), .X(n336) );
  SEN_ND2_S_0P5 U691 ( .A1(n297), .A2(B[30]), .X(n1256) );
  SEN_NR2_S_0P5 U693 ( .A1(B[7]), .A2(A[7]), .X(n260) );
  SEN_INV_S_0P5 U694 ( .A(n260), .X(n772) );
  SEN_ND2_S_0P5 U696 ( .A1(n611), .A2(n586), .X(n261) );
  SEN_INV_S_0P5 U697 ( .A(n261), .X(n562) );
  SEN_AOI21B_0P5 U698 ( .A1(n891), .A2(n959), .B(n927), .X(n262) );
  SEN_INV_S_0P5 U699 ( .A(n262), .X(n892) );
  SEN_ND3_S_0P5 U701 ( .A1(n1120), .A2(n1122), .A3(n1097), .X(n1070) );
  SEN_MAJ3_1 U702 ( .A1(B[25]), .A2(A[25]), .A3(n1233), .X(n1152) );
  SEN_ND2_S_0P5 U703 ( .A1(n514), .A2(INST[1]), .X(n507) );
  SEN_OAI21B_0P5 U704 ( .A1(n339), .A2(n1061), .B(n1065), .X(n1049) );
  SEN_ND2_S_0P5 U705 ( .A1(n1176), .A2(n1198), .X(n1202) );
  SEN_ND2_S_0P5 U706 ( .A1(n1245), .A2(n384), .X(n327) );
  SEN_ND2B_1 U707 ( .A(n975), .B(n974), .X(n976) );
  SEN_ND2_T_1 U709 ( .A1(n980), .A2(n979), .X(Z[19]) );
  SEN_MUXI2_S_2 U710 ( .D0(n977), .D1(n976), .S(A[19]), .X(n980) );
  SEN_NR2B_V1_1 U712 ( .A(n593), .B(n450), .X(n394) );
  SEN_AOAI211_0P75 U717 ( .A1(n442), .A2(n441), .B(n440), .C(n439), .X(n445)
         );
  SEN_ND2B_V1DG_1 U719 ( .A(B[16]), .B(A[16]), .X(n960) );
  SEN_BUF_1 U721 ( .A(B[13]), .X(n263) );
  SEN_AOI211_G_2 U722 ( .A1(n467), .A2(n466), .B1(n465), .B2(n464), .X(n468)
         );
  SEN_AOAI211_0P75 U723 ( .A1(n598), .A2(n616), .B(n452), .C(n451), .X(n466)
         );
  SEN_AOAI211_0P5 U725 ( .A1(A[19]), .A2(n978), .B(n297), .C(B[19]), .X(n979)
         );
  SEN_NR2B_V1_1 U727 ( .A(n637), .B(n643), .X(n451) );
  SEN_NR2_1 U730 ( .A1(n923), .A2(n890), .X(n894) );
  SEN_OAI22_1 U731 ( .A1(n895), .A2(n270), .B1(n897), .B2(n378), .X(n899) );
  SEN_MUXI2_DG_1 U733 ( .D0(n907), .D1(n906), .S(A[17]), .X(n908) );
  SEN_INV_0P65 U738 ( .A(n376), .X(n374) );
  SEN_ND2B_V1_2 U740 ( .A(A[12]), .B(B[12]), .X(n815) );
  SEN_OAI221_2 U742 ( .A1(n969), .A2(n370), .B1(n968), .B2(n378), .C(n374), 
        .X(n972) );
  SEN_INV_S_1P5 U747 ( .A(n1031), .X(n1029) );
  SEN_INV_4 U748 ( .A(n267), .X(n268) );
  SEN_OAI211_2 U750 ( .A1(n1173), .A2(n370), .B1(n375), .B2(n1172), .X(n1178)
         );
  SEN_AOAI211_0P5 U752 ( .A1(A[21]), .A2(n1037), .B(n1304), .C(B[21]), .X(
        n1038) );
  SEN_OAI211_1 U753 ( .A1(n1190), .A2(n271), .B1(n1189), .B2(n375), .X(n1196)
         );
  SEN_ND2_2 U755 ( .A1(n927), .A2(n926), .X(n928) );
  SEN_OA21_4 U756 ( .A1(n1150), .A2(n1149), .B(n1148), .X(n341) );
  SEN_OAI211_1 U757 ( .A1(n1200), .A2(A[27]), .B1(n299), .B2(n1199), .X(n1201)
         );
  SEN_ND2B_S_0P5 U760 ( .A(B[29]), .B(A[29]), .X(n1282) );
  SEN_INV_S_0P5 U761 ( .A(n1289), .X(n376) );
  SEN_NR2_S_0P5 U762 ( .A1(n1149), .A2(n486), .X(n408) );
  SEN_ND2B_S_0P5 U764 ( .A(B[26]), .B(A[26]), .X(n1164) );
  SEN_INV_0P5 U765 ( .A(n699), .X(n700) );
  SEN_INV_S_0P5 U767 ( .A(n1087), .X(n1077) );
  SEN_ND3_S_0P5 U768 ( .A1(n615), .A2(n658), .A3(n758), .X(n460) );
  SEN_ND2_0P5 U769 ( .A1(n410), .A2(n409), .X(n349) );
  SEN_NR2B_V1_1 U771 ( .A(n1041), .B(n472), .X(n473) );
  SEN_NR2B_V1_1 U772 ( .A(n713), .B(n438), .X(n396) );
  SEN_NR2B_V1_1 U773 ( .A(n761), .B(n782), .X(n400) );
  SEN_ND2B_S_0P5 U774 ( .A(A[10]), .B(n735), .X(n770) );
  SEN_NR3_0P5 U775 ( .A1(n1004), .A2(n1003), .A3(n1002), .X(n1011) );
  SEN_ND2_S_0P5 U776 ( .A1(A[1]), .A2(B[1]), .X(n586) );
  SEN_ND2B_S_0P5 U778 ( .A(B[5]), .B(A[5]), .X(n637) );
  SEN_ND2B_S_0P5 U779 ( .A(B[6]), .B(A[6]), .X(n764) );
  SEN_ND2B_V1DG_1 U780 ( .A(B[9]), .B(A[9]), .X(n731) );
  SEN_ND2B_S_0P5 U781 ( .A(B[10]), .B(A[10]), .X(n766) );
  SEN_INV_1P5 U783 ( .A(n815), .X(n864) );
  SEN_ND2B_S_0P5 U785 ( .A(B[11]), .B(A[11]), .X(n988) );
  SEN_ND2B_S_0P5 U787 ( .A(B[20]), .B(A[20]), .X(n1042) );
  SEN_ND2B_S_0P5 U788 ( .A(A[22]), .B(B[22]), .X(n1097) );
  SEN_INV_S_0P5 U789 ( .A(n485), .X(n1149) );
  SEN_INV_1P25 U790 ( .A(n500), .X(n503) );
  SEN_INV_0P65 U791 ( .A(INST[1]), .X(n522) );
  SEN_OR2_DG_1 U794 ( .A1(n305), .A2(n379), .X(n314) );
  SEN_INV_S_0P5 U795 ( .A(n373), .X(n271) );
  SEN_AN3B_0P5 U797 ( .B1(n1007), .B2(n953), .A(n294), .X(n955) );
  SEN_OR3B_2 U798 ( .B1(A[17]), .B2(A[18]), .A(n949), .X(n950) );
  SEN_ND4_2 U800 ( .A1(n1235), .A2(n1234), .A3(n1260), .A4(n1233), .X(n1237)
         );
  SEN_BUF_S_1 U801 ( .A(n554), .X(n288) );
  SEN_OAI22_S_0P5 U803 ( .A1(n661), .A2(n270), .B1(n674), .B2(n377), .X(n664)
         );
  SEN_INV_S_0P5 U805 ( .A(n1104), .X(n1105) );
  SEN_ND2_S_0P5 U806 ( .A1(n812), .A2(n811), .X(Z[13]) );
  SEN_ND2_S_0P5 U807 ( .A1(n824), .A2(n802), .X(n809) );
  SEN_ND2_S_0P8 U809 ( .A1(n1039), .A2(n1038), .X(Z[21]) );
  SEN_ND3_S_0P5 U810 ( .A1(n1162), .A2(n1161), .A3(n1160), .X(Z[26]) );
  SEN_ND2_4 U812 ( .A1(n769), .A2(n767), .X(n994) );
  SEN_MUXI2_DG_1 U815 ( .D0(n849), .D1(n848), .S(A[15]), .X(n850) );
  SEN_AOAI211_1 U819 ( .A1(n354), .A2(n910), .B(n909), .C(n908), .X(Z[17]) );
  SEN_INV_S_0P5 U820 ( .A(n376), .X(n375) );
  SEN_NR2B_V1_1 U822 ( .A(n988), .B(n782), .X(n439) );
  SEN_AOI21B_4 U825 ( .A1(n763), .A2(n762), .B(n761), .X(n769) );
  SEN_INV_0P8 U829 ( .A(n967), .X(n968) );
  SEN_ND2_4 U831 ( .A1(n738), .A2(n737), .X(n777) );
  SEN_MUXI2_S_1 U832 ( .D0(n940), .D1(n939), .S(n938), .X(n948) );
  SEN_ND2_T_2 U834 ( .A1(n1265), .A2(n1206), .X(n1233) );
  SEN_AOI211_3 U837 ( .A1(n383), .A2(n1028), .B1(n1027), .B2(n376), .X(n1031)
         );
  SEN_OR2_5 U838 ( .A1(n333), .A2(n334), .X(n1223) );
  SEN_ND2B_S_0P5 U840 ( .A(A[30]), .B(B[30]), .X(n1278) );
  SEN_ND2B_V1_1 U842 ( .A(n270), .B(n1173), .X(n1168) );
  SEN_NR2_S_0P5 U843 ( .A1(n638), .A2(n643), .X(n392) );
  SEN_OAI21_0P75 U844 ( .A1(n958), .A2(n1000), .B(n1006), .X(n969) );
  SEN_ND2B_S_0P5 U846 ( .A(B[22]), .B(A[22]), .X(n1067) );
  SEN_INV_S_0P5 U847 ( .A(n1251), .X(n1298) );
  SEN_INV_S_0P5 U848 ( .A(n474), .X(n469) );
  SEN_NR2_S_0P5 U849 ( .A1(n449), .A2(n448), .X(n467) );
  SEN_OAI21B_0P5 U851 ( .A1(n924), .A2(n871), .B(n471), .X(n475) );
  SEN_ND2_S_0P5 U852 ( .A1(n1096), .A2(n1097), .X(n1117) );
  SEN_INV_1 U853 ( .A(n349), .X(n350) );
  SEN_ND2_S_0P5 U854 ( .A1(B[11]), .A2(A[11]), .X(n1001) );
  SEN_INV_S_0P5 U855 ( .A(n773), .X(n774) );
  SEN_ND2B_S_1 U856 ( .A(n736), .B(n289), .X(n737) );
  SEN_OR2_1 U857 ( .A1(A[12]), .A2(B[12]), .X(n854) );
  SEN_INV_S_0P5 U858 ( .A(n1097), .X(n1068) );
  SEN_ND2B_1 U859 ( .A(n268), .B(B[28]), .X(n1242) );
  SEN_BUF_S_1 U861 ( .A(n1187), .X(n301) );
  SEN_NR2_S_0P5 U863 ( .A1(n1077), .A2(n298), .X(n1080) );
  SEN_ND2_S_0P5 U864 ( .A1(n459), .A2(n615), .X(n452) );
  SEN_INV_S_0P5 U865 ( .A(n731), .X(n438) );
  SEN_NR2_S_0P5 U866 ( .A1(n411), .A2(n1279), .X(n409) );
  SEN_ND3_1 U867 ( .A1(n416), .A2(n414), .A3(n413), .X(n415) );
  SEN_ND2_S_0P5 U869 ( .A1(n952), .A2(n951), .X(n1005) );
  SEN_ND2B_S_0P5 U871 ( .A(A[19]), .B(B[19]), .X(n1121) );
  SEN_INV_S_0P5 U872 ( .A(n616), .X(n613) );
  SEN_INV_S_0P5 U875 ( .A(n459), .X(n638) );
  SEN_OR2_1 U876 ( .A1(A[8]), .A2(B[8]), .X(n711) );
  SEN_INV_S_0P5 U878 ( .A(n885), .X(n1002) );
  SEN_AOI31_1 U879 ( .A1(n778), .A2(n777), .A3(n776), .B(n780), .X(n1008) );
  SEN_INV_S_0P5 U880 ( .A(n933), .X(n991) );
  SEN_INV_S_0P5 U881 ( .A(n1122), .X(n1100) );
  SEN_ND2B_S_0P5 U882 ( .A(B[30]), .B(A[30]), .X(n1283) );
  SEN_AOI21B_0P5 U883 ( .A1(n711), .A2(n692), .B(n709), .X(n344) );
  SEN_INV_S_0P5 U884 ( .A(B[10]), .X(n735) );
  SEN_INV_S_0P5 U886 ( .A(B[14]), .X(n832) );
  SEN_INV_S_0P5 U887 ( .A(n1016), .X(n1025) );
  SEN_AOAI211_0P5 U888 ( .A1(n1046), .A2(n1045), .B(n1061), .C(n1044), .X(
        n1065) );
  SEN_ND2B_S_0P5 U889 ( .A(n1032), .B(n388), .X(n1055) );
  SEN_ND2_S_0P5 U890 ( .A1(n1283), .A2(n1278), .X(n1246) );
  SEN_AOI211_0P5 U891 ( .A1(n1263), .A2(n1267), .B1(n1262), .B2(n1261), .X(
        n1276) );
  SEN_MUXI2_S_0P5 U892 ( .D0(n664), .D1(n667), .S(B[7]), .X(n665) );
  SEN_INV_S_0P5 U894 ( .A(n868), .X(n870) );
  SEN_ND2_S_0P5 U896 ( .A1(n383), .A2(n1163), .X(n1151) );
  SEN_ND3_S_0P5 U897 ( .A1(n603), .A2(n602), .A3(n601), .X(Z[4]) );
  SEN_ND2_S_0P5 U898 ( .A1(B[4]), .A2(n297), .X(n601) );
  SEN_AOAI211_0P5 U899 ( .A1(A[9]), .A2(n706), .B(n297), .C(B[9]), .X(n707) );
  SEN_ND2_S_0P5 U900 ( .A1(A[15]), .A2(n844), .X(n851) );
  SEN_ND3_S_0P5 U901 ( .A1(n1113), .A2(n1112), .A3(n1111), .X(Z[24]) );
  SEN_INV_S_0P5 U905 ( .A(INST[3]), .X(n528) );
  SEN_ND2B_V1DG_1 U908 ( .A(A[14]), .B(B[14]), .X(n861) );
  SEN_INV_S_0P5 U909 ( .A(n623), .X(n639) );
  SEN_AOAI211_0P5 U910 ( .A1(n919), .A2(n1315), .B(n917), .C(n916), .X(n277)
         );
  SEN_AO31_2 U911 ( .A1(n778), .A2(n777), .A3(n776), .B(n780), .X(n278) );
  SEN_OR3B_2 U913 ( .B1(A[9]), .B2(A[10]), .A(n742), .X(n743) );
  SEN_AN2_S_4 U914 ( .A1(n347), .A2(n1219), .X(n283) );
  SEN_ND2_S_0P5 U917 ( .A1(n884), .A2(n290), .X(n1003) );
  SEN_INV_S_0P5 U918 ( .A(n1251), .X(n295) );
  SEN_INV_S_0P5 U919 ( .A(n295), .X(n296) );
  SEN_AN2_S_0P5 U920 ( .A1(n510), .A2(n514), .X(n351) );
  SEN_INV_S_0P5 U921 ( .A(n354), .X(n297) );
  SEN_NR2_S_0P5 U924 ( .A1(n431), .A2(n300), .X(n420) );
  SEN_ND2_2 U926 ( .A1(n1221), .A2(n389), .X(n347) );
  SEN_AN4B_1 U927 ( .B1(n1120), .B2(n469), .B3(n1122), .A(n468), .X(n480) );
  SEN_INV_1 U928 ( .A(n504), .X(n505) );
  SEN_AOA211_DG_1 U929 ( .A1(n894), .A2(n893), .B(n892), .C(n960), .X(n305) );
  SEN_AOA211_DG_1 U930 ( .A1(n1274), .A2(n1273), .B(n1272), .C(n1271), .X(n306) );
  SEN_OR2_1 U932 ( .A1(n695), .A2(n377), .X(n308) );
  SEN_INV_S_0P5 U933 ( .A(n384), .X(n377) );
  SEN_BUF_1 U934 ( .A(n1114), .X(n309) );
  SEN_MUXI2_DG_3 U935 ( .D0(n1303), .D1(n1302), .S(A[31]), .X(n1307) );
  SEN_AOAI211_1 U936 ( .A1(n838), .A2(n865), .B(n837), .C(n862), .X(n841) );
  SEN_AOAI211_1 U937 ( .A1(n888), .A2(n274), .B(n887), .C(n951), .X(n898) );
  SEN_ND2_S_0P5 U938 ( .A1(n764), .A2(n766), .X(n315) );
  SEN_OR2_DG_1 U939 ( .A1(n843), .A2(n270), .X(n316) );
  SEN_OR2_1 U940 ( .A1(n842), .A2(n379), .X(n317) );
  SEN_INV_S_0P5 U941 ( .A(n482), .X(n1108) );
  SEN_OAI21_S_0P5 U942 ( .A1(n932), .A2(n931), .B(n930), .X(n963) );
  SEN_OR2_2P5 U943 ( .A1(n335), .A2(n376), .X(n334) );
  SEN_OAI21_S_0P5 U944 ( .A1(n1107), .A2(n271), .B(n1106), .X(n1109) );
  SEN_INV_S_0P5 U945 ( .A(n1240), .X(n411) );
  SEN_ND2B_S_0P5 U947 ( .A(B[14]), .B(A[14]), .X(n862) );
  SEN_ND2_S_0P5 U948 ( .A1(n1298), .A2(B[31]), .X(n321) );
  SEN_INV_S_0P5 U949 ( .A(B[31]), .X(n319) );
  SEN_INV_S_0P5 U950 ( .A(n960), .X(n931) );
  SEN_ND2_S_0P5 U951 ( .A1(n1013), .A2(n1012), .X(n339) );
  SEN_OR3B_0P5 U952 ( .B1(A[11]), .B2(A[12]), .A(n795), .X(n323) );
  SEN_INV_S_4 U953 ( .A(n1171), .X(n1218) );
  SEN_AN3B_0P5 U954 ( .B1(n1007), .B2(n1006), .A(n1005), .X(n1010) );
  SEN_ND2B_S_0P5 U956 ( .A(n1137), .B(n388), .X(n1157) );
  SEN_ND2_S_0P5 U957 ( .A1(n1298), .A2(B[27]), .X(n331) );
  SEN_OR3B_4 U958 ( .B1(A[25]), .B2(A[26]), .A(n1170), .X(n1171) );
  SEN_OR2_DG_1 U959 ( .A1(A[5]), .A2(B[5]), .X(n329) );
  SEN_ND2_S_0P5 U960 ( .A1(n383), .A2(n1213), .X(n1192) );
  SEN_ND2_S_0P5 U961 ( .A1(A[8]), .A2(B[8]), .X(n709) );
  SEN_ND2_S_0P5 U962 ( .A1(B[25]), .A2(A[25]), .X(n1207) );
  SEN_ND2_S_0P5 U963 ( .A1(A[10]), .A2(B[10]), .X(n778) );
  SEN_ND2B_S_0P5 U964 ( .A(n380), .B(n1050), .X(n1048) );
  SEN_INV_S_0P5 U965 ( .A(n1001), .X(n1004) );
  SEN_INV_S_0P5 U966 ( .A(n1117), .X(n1118) );
  SEN_INV_S_0P5 U967 ( .A(n1282), .X(n1279) );
  SEN_AOA211_DG_1 U968 ( .A1(n1042), .A2(n1041), .B(n1066), .C(n1040), .X(n342) );
  SEN_INV_S_0P5 U969 ( .A(n1243), .X(n417) );
  SEN_ND2B_S_0P5 U970 ( .A(B[2]), .B(n241), .X(n591) );
  SEN_ND2B_S_0P5 U971 ( .A(A[5]), .B(B[5]), .X(n459) );
  SEN_ND2_S_0P5 U972 ( .A1(A[26]), .A2(B[26]), .X(n1267) );
  SEN_INV_S_0P5 U973 ( .A(n389), .X(n386) );
  SEN_ND2_S_0P5 U974 ( .A1(n383), .A2(n1150), .X(n1130) );
  SEN_AO2BB2_0P5 U975 ( .A1(n718), .A2(n379), .B1(n272), .B2(n717), .X(n721)
         );
  SEN_INV_S_0P5 U976 ( .A(n472), .X(n1017) );
  SEN_INV_S_0P5 U977 ( .A(n453), .X(n678) );
  SEN_BUF_AS_0P5 U978 ( .A(n389), .X(n388) );
  SEN_ND2_S_0P5 U979 ( .A1(n713), .A2(n714), .X(n453) );
  SEN_ND2_S_0P5 U980 ( .A1(n389), .A2(n1131), .X(n1087) );
  SEN_NR2_S_0P5 U981 ( .A1(n1100), .A2(n470), .X(n479) );
  SEN_ND2B_S_0P5 U982 ( .A(n902), .B(n388), .X(n943) );
  SEN_OAI21_S_0P5 U983 ( .A1(n1206), .A2(n250), .B(n1231), .X(n1208) );
  SEN_INV_S_0P5 U984 ( .A(n424), .X(n1051) );
  SEN_ND2_S_0P5 U985 ( .A1(n1243), .A2(n1242), .X(n1277) );
  SEN_ND2_S_0P5 U986 ( .A1(n539), .A2(n538), .X(n540) );
  SEN_MUXI2_S_0P5 U987 ( .D0(n534), .D1(n537), .S(B[1]), .X(n535) );
  SEN_NR2_S_0P5 U988 ( .A1(A[11]), .A2(B[11]), .X(n773) );
  SEN_ND2_S_0P5 U989 ( .A1(n862), .A2(n865), .X(n990) );
  SEN_ND2_S_0P5 U990 ( .A1(n1298), .A2(B[29]), .X(n348) );
  SEN_INV_S_0P5 U991 ( .A(B[7]), .X(n675) );
  SEN_INV_S_0P5 U992 ( .A(n383), .X(n380) );
  SEN_OAI21_S_0P5 U994 ( .A1(n691), .A2(n385), .B(n1219), .X(n681) );
  SEN_OAI21_S_0P5 U995 ( .A1(n814), .A2(n833), .B(n884), .X(n818) );
  SEN_AOAI211_0P5 U996 ( .A1(n816), .A2(n989), .B(n836), .C(n1310), .X(n819)
         );
  SEN_AOI221_2 U997 ( .A1(n481), .A2(n480), .B1(n479), .B2(n478), .C(n477), 
        .X(n484) );
  SEN_OAI21_S_0P5 U998 ( .A1(n1023), .A2(n385), .B(n1219), .X(n981) );
  SEN_OAI21_S_0P5 U999 ( .A1(n740), .A2(n739), .B(n332), .X(n746) );
  SEN_INV_S_0P5 U1000 ( .A(n486), .X(n1153) );
  SEN_ND2_S_0P5 U1001 ( .A1(n1051), .A2(n1120), .X(n430) );
  SEN_ND2_S_0P5 U1002 ( .A1(n930), .A2(n927), .X(n471) );
  SEN_OAI21_S_0P5 U1003 ( .A1(n1150), .A2(n1149), .B(n1148), .X(n1163) );
  SEN_ND2_S_0P5 U1004 ( .A1(n960), .A2(n959), .X(n992) );
  SEN_ND2_S_0P5 U1005 ( .A1(n1041), .A2(n993), .X(n428) );
  SEN_INV_S_0P5 U1008 ( .A(n658), .X(n449) );
  SEN_ND3_S_0P5 U1009 ( .A1(n1122), .A2(n1121), .A3(n1120), .X(n1126) );
  SEN_OR3B_0P5 U1010 ( .B1(n522), .B2(INST[3]), .A(n351), .X(n1251) );
  SEN_ND2_S_0P5 U1011 ( .A1(n1243), .A2(n1242), .X(n494) );
  SEN_AOI21B_1 U1012 ( .A1(n445), .A2(n444), .B(n443), .X(n446) );
  SEN_ND2_S_0P5 U1013 ( .A1(A[16]), .A2(B[16]), .X(n951) );
  SEN_ND2B_S_0P5 U1014 ( .A(A[7]), .B(B[7]), .X(n758) );
  SEN_ND2B_S_0P5 U1015 ( .A(A[11]), .B(B[11]), .X(n761) );
  SEN_ND2_S_0P5 U1016 ( .A1(A[6]), .A2(B[6]), .X(n776) );
  SEN_ND3_S_0P5 U1017 ( .A1(n759), .A2(n758), .A3(n757), .X(n763) );
  SEN_INV_S_0P5 U1018 ( .A(n355), .X(n1219) );
  SEN_ND2_S_0P5 U1019 ( .A1(B[24]), .A2(n297), .X(n1111) );
  SEN_INV_S_0P5 U1020 ( .A(n354), .X(n1304) );
  SEN_INV_S_0P5 U1021 ( .A(A[15]), .X(n852) );
  SEN_ND2B_S_0P5 U1022 ( .A(A[1]), .B(B[1]), .X(n458) );
  SEN_INV_S_0P5 U1023 ( .A(B[1]), .X(n551) );
  SEN_OR3B_4 U1024 ( .B1(A[5]), .B2(A[6]), .A(n659), .X(n660) );
  SEN_OAI211_0P5 U1025 ( .A1(n717), .A2(n370), .B1(n716), .B2(n374), .X(n722)
         );
  SEN_ND2B_S_0P5 U1026 ( .A(n380), .B(n718), .X(n716) );
  SEN_OAI221_0P5 U1027 ( .A1(n550), .A2(n270), .B1(n379), .B2(n533), .C(n374), 
        .X(n537) );
  SEN_INV_S_0P5 U1028 ( .A(n566), .X(n567) );
  SEN_OAI221_0P5 U1029 ( .A1(n797), .A2(n379), .B1(n796), .B2(n270), .C(n374), 
        .X(n785) );
  SEN_OAI221_0P5 U1030 ( .A1(n694), .A2(n379), .B1(n692), .B2(n270), .C(n374), 
        .X(n680) );
  SEN_ND2_S_0P5 U1031 ( .A1(n383), .A2(n1132), .X(n1133) );
  SEN_INV_S_0P5 U1032 ( .A(n801), .X(n798) );
  SEN_OAI22_S_0P5 U1033 ( .A1(n565), .A2(n270), .B1(n566), .B2(n377), .X(n575)
         );
  SEN_INV_S_0P5 U1034 ( .A(n568), .X(n565) );
  SEN_INV_S_0P5 U1035 ( .A(n898), .X(n895) );
  SEN_ND2B_S_0P5 U1036 ( .A(n380), .B(n935), .X(n936) );
  SEN_OAI211_0P5 U1037 ( .A1(n818), .A2(n271), .B1(n817), .B2(n374), .X(n823)
         );
  SEN_ND2B_S_0P5 U1038 ( .A(n379), .B(n819), .X(n817) );
  SEN_OAI211_0P5 U1039 ( .A1(n596), .A2(n270), .B1(n375), .B2(n595), .X(n600)
         );
  SEN_ND2_S_0P5 U1040 ( .A1(n383), .A2(n597), .X(n595) );
  SEN_OAI22_S_0P5 U1041 ( .A1(n271), .A2(n820), .B1(n819), .B2(n377), .X(n822)
         );
  SEN_INV_S_0P5 U1042 ( .A(n818), .X(n820) );
  SEN_OAI22_S_0P5 U1043 ( .A1(n562), .A2(n271), .B1(n563), .B2(n377), .X(n556)
         );
  SEN_OAI21_S_0P5 U1044 ( .A1(n1066), .A2(n1069), .B(n342), .X(n1050) );
  SEN_AO2BB2_0P5 U1045 ( .A1(n597), .A2(n379), .B1(n272), .B2(n596), .X(n599)
         );
  SEN_AO2BB2_0P5 U1046 ( .A1(n1050), .A2(n379), .B1(n272), .B2(n1049), .X(
        n1052) );
  SEN_AO2BB2_0P5 U1047 ( .A1(n1016), .A2(n379), .B1(n272), .B2(n1015), .X(
        n1018) );
  SEN_AO2BB2_0P5 U1048 ( .A1(n677), .A2(n379), .B1(n373), .B2(n692), .X(n679)
         );
  SEN_ND2_S_0P5 U1049 ( .A1(n272), .A2(n746), .X(n741) );
  SEN_ND2_S_0P5 U1050 ( .A1(n883), .A2(n1009), .X(n796) );
  SEN_ND2_S_0P5 U1051 ( .A1(n304), .A2(n995), .X(n781) );
  SEN_INV_S_0P5 U1052 ( .A(n676), .X(n661) );
  SEN_INV_S_0P5 U1053 ( .A(n611), .X(n587) );
  SEN_ND3_S_0P5 U1054 ( .A1(n375), .A2(n641), .A3(n640), .X(n646) );
  SEN_ND2_S_0P5 U1055 ( .A1(n272), .A2(n642), .X(n641) );
  SEN_ND2_S_0P5 U1056 ( .A1(n383), .A2(n1312), .X(n640) );
  SEN_ND2B_S_0P5 U1057 ( .A(n1049), .B(n272), .X(n1047) );
  SEN_OAI211_0P5 U1058 ( .A1(n1025), .A2(n379), .B1(n375), .B2(n1014), .X(
        n1019) );
  SEN_ND2_S_0P5 U1059 ( .A1(n373), .A2(n1024), .X(n1014) );
  SEN_INV_S_0P5 U1060 ( .A(n782), .X(n783) );
  SEN_INV_S_0P5 U1061 ( .A(n1269), .X(n1262) );
  SEN_INV_S_0P5 U1062 ( .A(n643), .X(n644) );
  SEN_OAI211_0P5 U1063 ( .A1(n663), .A2(n379), .B1(n375), .B2(n662), .X(n667)
         );
  SEN_INV_S_0P5 U1064 ( .A(n674), .X(n663) );
  SEN_ND2_S_0P5 U1065 ( .A1(n272), .A2(n661), .X(n662) );
  SEN_INV_S_0P5 U1066 ( .A(n1268), .X(n1274) );
  SEN_INV_S_0P5 U1067 ( .A(n544), .X(n536) );
  SEN_INV_S_0P5 U1068 ( .A(n981), .X(n971) );
  SEN_INV_S_0P5 U1069 ( .A(n1005), .X(n953) );
  SEN_INV_S_0P5 U1070 ( .A(n736), .X(n712) );
  SEN_ND2_S_0P5 U1071 ( .A1(n383), .A2(n1104), .X(n1103) );
  SEN_NR2B_V1_1 U1072 ( .A(n1094), .B(n482), .X(n483) );
  SEN_INV_S_0P5 U1073 ( .A(n841), .X(n842) );
  SEN_AO21B_1 U1074 ( .A1(n1231), .A2(n1229), .B(n1236), .X(n1210) );
  SEN_NR3B_1 U1075 ( .A(n993), .B1(n992), .B2(n991), .X(n996) );
  SEN_ND2_S_0P5 U1076 ( .A1(n1191), .A2(n384), .X(n1189) );
  SEN_OAI22_S_0P5 U1077 ( .A1(n622), .A2(n370), .B1(n1313), .B2(n377), .X(n632) );
  SEN_INV_S_0P5 U1078 ( .A(n325), .X(n622) );
  SEN_ND3_S_0P5 U1079 ( .A1(n459), .A2(n592), .A3(n593), .X(n461) );
  SEN_INV_S_0P5 U1080 ( .A(n288), .X(n463) );
  SEN_AN2_S_0P5 U1081 ( .A1(n528), .A2(n522), .X(n352) );
  SEN_INV_S_0P5 U1082 ( .A(n951), .X(n917) );
  SEN_AOAI211_0P5 U1083 ( .A1(n894), .A2(n893), .B(n892), .C(n960), .X(n897)
         );
  SEN_INV_S_0P5 U1084 ( .A(n921), .X(n893) );
  SEN_INV_S_0P5 U1085 ( .A(n1242), .X(n1212) );
  SEN_ND2_S_0P5 U1086 ( .A1(n1120), .A2(n1122), .X(n1066) );
  SEN_INV_S_0P5 U1087 ( .A(n714), .X(n693) );
  SEN_NR3_0P5 U1088 ( .A1(n813), .A2(n1002), .A3(n294), .X(n814) );
  SEN_AOAI211_0P5 U1089 ( .A1(n732), .A2(n353), .B(n730), .C(n731), .X(n718)
         );
  SEN_AOAI211_0P5 U1090 ( .A1(n620), .A2(n594), .B(n617), .C(n616), .X(n597)
         );
  SEN_INV_S_0P5 U1091 ( .A(n614), .X(n594) );
  SEN_OAI21_S_0P5 U1092 ( .A1(n934), .A2(n963), .B(n933), .X(n935) );
  SEN_NR3_0P5 U1093 ( .A1(n923), .A2(n922), .A3(n921), .X(n934) );
  SEN_ND2_S_0P5 U1094 ( .A1(n960), .A2(n995), .X(n922) );
  SEN_OAI22_S_0P5 U1095 ( .A1(n532), .A2(n370), .B1(n378), .B2(n531), .X(n534)
         );
  SEN_OAI21_S_0P5 U1096 ( .A1(n462), .A2(n564), .B(n591), .X(n566) );
  SEN_INV_S_0P5 U1097 ( .A(n592), .X(n564) );
  SEN_NR3_0P5 U1098 ( .A1(n954), .A2(n1003), .A3(n294), .X(n859) );
  SEN_ND2_S_0P5 U1099 ( .A1(n678), .A2(n758), .X(n397) );
  SEN_ND2_S_0P5 U1100 ( .A1(n637), .A2(n618), .X(n393) );
  SEN_INV_S_0P5 U1101 ( .A(n889), .X(n405) );
  SEN_ND2_S_0P5 U1102 ( .A1(n821), .A2(n860), .X(n404) );
  SEN_AN2_S_0P5 U1103 ( .A1(n485), .A2(n1119), .X(n490) );
  SEN_ND2_S_0P5 U1104 ( .A1(n1153), .A2(n1148), .X(n489) );
  SEN_OAI21B_0P5 U1105 ( .A1(n1308), .A2(n732), .B(n760), .X(n744) );
  SEN_ND2_S_0P5 U1106 ( .A1(n1235), .A2(n1260), .X(n1229) );
  SEN_ND2_S_0P5 U1107 ( .A1(n960), .A2(n927), .X(n871) );
  SEN_NR3_0P5 U1108 ( .A1(n913), .A2(n912), .A3(n911), .X(n920) );
  SEN_ND2_S_0P5 U1109 ( .A1(n274), .A2(n951), .X(n912) );
  SEN_INV_S_0P5 U1110 ( .A(n1003), .X(n956) );
  SEN_OAI21B_0P5 U1111 ( .A1(n386), .A2(n560), .B(n544), .X(n549) );
  SEN_INV_S_0P5 U1112 ( .A(n1096), .X(n1095) );
  SEN_OAI21_S_0P5 U1113 ( .A1(n589), .A2(n608), .B(n607), .X(n596) );
  SEN_NR2_S_0P5 U1114 ( .A1(n606), .A2(n587), .X(n589) );
  SEN_ND2_S_0P5 U1115 ( .A1(n1234), .A2(n1235), .X(n1263) );
  SEN_OAI21_S_0P5 U1116 ( .A1(n303), .A2(n562), .B(n585), .X(n568) );
  SEN_ND2_S_0P5 U1117 ( .A1(n865), .A2(n989), .X(n889) );
  SEN_NR2_S_0P5 U1118 ( .A1(n425), .A2(n430), .X(n407) );
  SEN_OAI21_S_0P5 U1119 ( .A1(n949), .A2(n385), .B(n1219), .X(n941) );
  SEN_ND4B_1 U1120 ( .A(n429), .B1(n428), .B2(n427), .B3(n426), .X(n436) );
  SEN_INV_S_0P5 U1121 ( .A(n1166), .X(n1266) );
  SEN_ND2_S_0P5 U1122 ( .A1(n1206), .A2(n1207), .X(n1166) );
  SEN_NR3B_1 U1123 ( .A(n731), .B1(n719), .B2(n782), .X(n456) );
  SEN_ND2_S_0P5 U1124 ( .A1(n1121), .A2(n964), .X(n474) );
  SEN_ND2_S_0P5 U1125 ( .A1(n383), .A2(n1105), .X(n1106) );
  SEN_INV_S_0P5 U1126 ( .A(n1241), .X(n1281) );
  SEN_ND2_S_0P5 U1127 ( .A1(n1240), .A2(n1239), .X(n1241) );
  SEN_ND2_S_0P5 U1128 ( .A1(n926), .A2(n925), .X(n891) );
  SEN_INV_S_0P5 U1129 ( .A(n656), .X(n642) );
  SEN_OAI21_S_0P5 U1130 ( .A1(n386), .A2(n545), .B(n1219), .X(n544) );
  SEN_NR2_S_0P5 U1131 ( .A1(n1279), .A2(n1246), .X(n493) );
  SEN_ND2_S_0P5 U1132 ( .A1(n915), .A2(n914), .X(n886) );
  SEN_ND2_S_0P5 U1133 ( .A1(n860), .A2(n815), .X(n836) );
  SEN_INV_S_0P5 U1134 ( .A(n1120), .X(n470) );
  SEN_ND2_S_0P5 U1135 ( .A1(n854), .A2(n855), .X(n833) );
  SEN_ND2_S_0P5 U1136 ( .A1(n1042), .A2(n1122), .X(n472) );
  SEN_ND2_S_0P5 U1137 ( .A1(n1231), .A2(n1230), .X(n1268) );
  SEN_OR4B_1 U1138 ( .B1(n412), .B2(n411), .B3(n1279), .A(n410), .X(n414) );
  SEN_ND2_S_0P5 U1139 ( .A1(n1148), .A2(n1115), .X(n412) );
  SEN_ND2_S_0P5 U1140 ( .A1(n933), .A2(n960), .X(n421) );
  SEN_INV_S_0P5 U1141 ( .A(n454), .X(n821) );
  SEN_INV_S_0P5 U1142 ( .A(n531), .X(n533) );
  SEN_ND2B_S_0P5 U1143 ( .A(n701), .B(n388), .X(n725) );
  SEN_ND2B_S_0P5 U1144 ( .A(n323), .B(n388), .X(n826) );
  SEN_ND2B_S_0P5 U1145 ( .A(n627), .B(n389), .X(n649) );
  SEN_ND2_S_0P5 U1146 ( .A1(n1017), .A2(n1121), .X(n425) );
  SEN_ND2_S_0P5 U1147 ( .A1(n1259), .A2(n1273), .X(n1269) );
  SEN_ND2_S_0P5 U1148 ( .A1(n1115), .A2(n1119), .X(n482) );
  SEN_INV_S_0P5 U1149 ( .A(n758), .X(n448) );
  SEN_OR4B_1 U1150 ( .B1(n418), .B2(n1246), .B3(n417), .A(n416), .X(n419) );
  SEN_ND2_S_0P5 U1151 ( .A1(n1108), .A2(n1096), .X(n418) );
  SEN_ND2B_S_0P5 U1152 ( .A(n301), .B(n383), .X(n1169) );
  SEN_ND2_S_0P5 U1153 ( .A1(n389), .A2(n691), .X(n685) );
  SEN_ND2_S_0P5 U1154 ( .A1(n1270), .A2(n1269), .X(n1272) );
  SEN_INV_S_0P5 U1155 ( .A(n1246), .X(n1247) );
  SEN_INV_S_0P5 U1156 ( .A(n719), .X(n720) );
  SEN_NR2_S_0P5 U1157 ( .A1(n425), .A2(n424), .X(n426) );
  SEN_ND2_S_0P5 U1158 ( .A1(n1051), .A2(n1040), .X(n477) );
  SEN_INV_S_0P5 U1159 ( .A(n1260), .X(n1261) );
  SEN_BUF_AS_0P5 U1160 ( .A(n384), .X(n383) );
  SEN_ND2_S_0P5 U1161 ( .A1(n553), .A2(n552), .X(n555) );
  SEN_ND2_S_0P5 U1162 ( .A1(n384), .A2(n563), .X(n552) );
  SEN_AOI21_S_0P5 U1163 ( .A1(n272), .A2(n562), .B(n376), .X(n553) );
  SEN_MUXI2_S_0P5 U1164 ( .D0(n1089), .D1(n1088), .S(A[24]), .X(n1113) );
  SEN_ND4_S_0P5 U1165 ( .A1(INST[3]), .A2(INST[2]), .A3(INST[1]), .A4(INST[0]), 
        .X(n216) );
  SEN_OAI221_0P5 U1166 ( .A1(n1251), .A2(n650), .B1(n649), .B2(A[5]), .C(n1300), .X(n651) );
  SEN_INV_S_0P5 U1167 ( .A(B[6]), .X(n650) );
  SEN_OAI221_0P5 U1168 ( .A1(n1251), .A2(n735), .B1(n725), .B2(A[9]), .C(n1300), .X(n726) );
  SEN_OAI221_0P5 U1169 ( .A1(n1251), .A2(n832), .B1(n826), .B2(A[13]), .C(
        n1300), .X(n827) );
  SEN_OAI221_0P5 U1170 ( .A1(n1251), .A2(n944), .B1(n943), .B2(A[17]), .C(
        n1300), .X(n945) );
  SEN_INV_S_0P5 U1171 ( .A(B[18]), .X(n944) );
  SEN_AO21B_1 U1172 ( .A1(n833), .A2(n884), .B(n856), .X(n834) );
  SEN_INV_S_0P5 U1173 ( .A(n884), .X(n831) );
  SEN_ND2_S_0P5 U1174 ( .A1(A[4]), .A2(B[4]), .X(n609) );
  SEN_ND2B_S_0P5 U1175 ( .A(B[18]), .B(A[18]), .X(n993) );
  SEN_ND2_S_0P5 U1176 ( .A1(B[23]), .A2(A[23]), .X(n1090) );
  SEN_INV_S_0P5 U1177 ( .A(A[23]), .X(n1092) );
  SEN_MUXI2_S_0P5 U1178 ( .D0(n575), .D1(n570), .S(B[3]), .X(n569) );
  SEN_MUXI2_S_0P5 U1179 ( .D0(n632), .D1(n625), .S(B[5]), .X(n624) );
  SEN_MUXI2_S_0P5 U1180 ( .D0(n810), .D1(n803), .S(B[13]), .X(n802) );
  SEN_OAI21_S_0P5 U1181 ( .A1(n1280), .A2(n1279), .B(n1278), .X(n1286) );
  SEN_INV_S_0P5 U1182 ( .A(n1277), .X(n1280) );
  SEN_MUXI2_S_0P5 U1183 ( .D0(n1057), .D1(n1056), .S(A[22]), .X(n1058) );
  SEN_OAI21_S_0P5 U1184 ( .A1(n1054), .A2(n385), .B(n236), .X(n1057) );
  SEN_INV_S_0P5 U1185 ( .A(A[21]), .X(n1054) );
  SEN_ND2_S_0P5 U1186 ( .A1(B[27]), .A2(A[27]), .X(n1231) );
  SEN_ND2_S_0P5 U1187 ( .A1(n1207), .A2(n1267), .X(n1232) );
  SEN_OAI211_0P5 U1188 ( .A1(n984), .A2(A[19]), .B1(n299), .B2(n983), .X(n985)
         );
  SEN_ND2B_S_0P5 U1189 ( .A(n1251), .B(B[20]), .X(n983) );
  SEN_OAI211_0P5 U1190 ( .A1(n877), .A2(A[15]), .B1(n299), .B2(n876), .X(n878)
         );
  SEN_ND2_S_0P5 U1191 ( .A1(B[16]), .A2(n1298), .X(n876) );
  SEN_OAI211_0P5 U1192 ( .A1(n685), .A2(A[7]), .B1(n299), .B2(n684), .X(n686)
         );
  SEN_ND2_S_0P5 U1193 ( .A1(B[8]), .A2(n1298), .X(n684) );
  SEN_OAI211_0P5 U1194 ( .A1(n789), .A2(A[11]), .B1(n299), .B2(n788), .X(n790)
         );
  SEN_ND2_S_0P5 U1195 ( .A1(B[12]), .A2(n1298), .X(n788) );
  SEN_OAI211_0P5 U1196 ( .A1(n1087), .A2(A[23]), .B1(n299), .B2(n1086), .X(
        n1088) );
  SEN_ND2B_S_0P5 U1197 ( .A(n1251), .B(B[24]), .X(n1086) );
  SEN_INV_S_0P5 U1198 ( .A(A[0]), .X(n545) );
  SEN_MUXI2_S_0P5 U1199 ( .D0(n706), .D1(n699), .S(B[9]), .X(n698) );
  SEN_ND2B_S_0P5 U1200 ( .A(A[24]), .B(B[24]), .X(n1119) );
  SEN_AO21B_1 U1201 ( .A1(n383), .A2(n1074), .B(n1073), .X(n1078) );
  SEN_MUXI2_S_0P5 U1202 ( .D0(n600), .D1(n599), .S(n598), .X(n602) );
  SEN_MUXI2_S_0P5 U1203 ( .D0(n584), .D1(n583), .S(A[4]), .X(n603) );
  SEN_AOI21_S_0P5 U1204 ( .A1(n523), .A2(n518), .B(n517), .X(n519) );
  SEN_ND2_S_0P5 U1205 ( .A1(n386), .A2(n1300), .X(n517) );
  SEN_ND2_S_0P5 U1206 ( .A1(B[29]), .A2(A[29]), .X(n1273) );
  SEN_AOAI211_0P5 U1207 ( .A1(n354), .A2(n1084), .B(n1093), .C(n1083), .X(
        Z[23]) );
  SEN_ND2_S_0P5 U1208 ( .A1(A[23]), .A2(n1075), .X(n1084) );
  SEN_MUXI2_S_0P5 U1209 ( .D0(n1082), .D1(n1081), .S(A[23]), .X(n1083) );
  SEN_AOAI211_0P5 U1210 ( .A1(n354), .A2(n756), .B(n755), .C(n754), .X(Z[11])
         );
  SEN_INV_S_0P5 U1211 ( .A(B[11]), .X(n755) );
  SEN_ND2_S_0P5 U1212 ( .A1(A[11]), .A2(n747), .X(n756) );
  SEN_ND2B_S_0P5 U1214 ( .A(A[23]), .B(B[23]), .X(n1096) );
  SEN_ND3B_0P5 U1215 ( .A(B[0]), .B1(A[0]), .B2(n458), .X(n391) );
  SEN_NR2B_V1_1 U1216 ( .A(n591), .B(n613), .X(n390) );
  SEN_ND2_S_0P5 U1217 ( .A1(n766), .A2(n988), .X(n401) );
  SEN_ND2_S_0P5 U1218 ( .A1(n959), .A2(n862), .X(n921) );
  SEN_OAI21_S_0P5 U1219 ( .A1(A[29]), .A2(B[29]), .B(n1236), .X(n1259) );
  SEN_AN2_S_0P5 U1220 ( .A1(n216), .A2(n530), .X(n354) );
  SEN_EN2_0P5 U1222 ( .A1(INST[0]), .A2(n515), .X(n516) );
  SEN_ND2B_S_0P5 U1223 ( .A(A[26]), .B(n1167), .X(n1235) );
  SEN_ND2B_S_0P5 U1224 ( .A(A[18]), .B(B[18]), .X(n964) );
  SEN_ND2_S_0P5 U1225 ( .A1(n715), .A2(n714), .X(n441) );
  SEN_ND2_S_0P5 U1226 ( .A1(A[24]), .A2(B[24]), .X(n1206) );
  SEN_ND2B_S_0P5 U1227 ( .A(B[25]), .B(A[25]), .X(n1148) );
  SEN_ND2B_S_0P5 U1228 ( .A(B[23]), .B(A[23]), .X(n1094) );
  SEN_ND2B_S_0P5 U1229 ( .A(n386), .B(A[30]), .X(n1296) );
  SEN_INV_S_0P5 U1230 ( .A(B[0]), .X(n523) );
  SEN_ND2_S_0P5 U1231 ( .A1(n1067), .A2(n1097), .X(n424) );
  SEN_INV_S_0P5 U1232 ( .A(n487), .X(n1165) );
  SEN_ND3_S_0P5 U1233 ( .A1(n1067), .A2(n1094), .A3(n345), .X(n434) );
  SEN_ND3_S_0P5 U1234 ( .A1(n299), .A2(n547), .A3(n546), .X(n548) );
  SEN_ND2_S_0P5 U1235 ( .A1(B[2]), .A2(n1298), .X(n546) );
  SEN_ND3B_0P5 U1236 ( .A(n386), .B1(n545), .B2(n560), .X(n547) );
  SEN_ND2_S_0P5 U1237 ( .A1(n1185), .A2(n1184), .X(n1260) );
  SEN_INV_S_0P5 U1238 ( .A(A[27]), .X(n1184) );
  SEN_INV_S_0P5 U1239 ( .A(B[23]), .X(n1093) );
  SEN_ND2B_S_0P5 U1240 ( .A(A[29]), .B(B[29]), .X(n1243) );
  SEN_ND2B_S_0P5 U1241 ( .A(B[24]), .B(A[24]), .X(n1115) );
  SEN_INV_S_0P5 U1242 ( .A(n471), .X(n447) );
  SEN_ND2_S_0P5 U1243 ( .A1(A[20]), .A2(B[20]), .X(n1045) );
  SEN_ND2B_S_0P5 U1244 ( .A(A[30]), .B(n1264), .X(n1270) );
  SEN_INV_S_0P5 U1245 ( .A(B[29]), .X(n1227) );
  SEN_ND2_S_0P5 U1246 ( .A1(A[25]), .A2(n1134), .X(n1145) );
  SEN_ND2_S_0P5 U1247 ( .A1(A[27]), .A2(n1174), .X(n1183) );
  SEN_AOAI211_0P5 U1248 ( .A1(n354), .A2(n673), .B(n675), .C(n672), .X(Z[7])
         );
  SEN_ND2_S_0P5 U1249 ( .A1(A[7]), .A2(n664), .X(n673) );
  SEN_MUXI2_S_0P5 U1250 ( .D0(n671), .D1(n670), .S(A[7]), .X(n672) );
  SEN_ND2_S_0P5 U1251 ( .A1(n682), .A2(n665), .X(n671) );
  SEN_AOAI211_0P5 U1252 ( .A1(n354), .A2(n543), .B(n551), .C(n542), .X(Z[1])
         );
  SEN_ND2_S_0P5 U1253 ( .A1(A[1]), .A2(n534), .X(n543) );
  SEN_MUXI2_S_0P5 U1254 ( .D0(n541), .D1(n540), .S(A[1]), .X(n542) );
  SEN_ND2_S_0P5 U1255 ( .A1(n536), .A2(n535), .X(n541) );
  SEN_INV_S_0P5 U1256 ( .A(B[17]), .X(n909) );
  SEN_ND2_S_0P5 U1257 ( .A1(A[17]), .A2(n899), .X(n910) );
  SEN_ND3B_0P5 U1258 ( .A(n582), .B1(n581), .B2(n299), .X(n583) );
  SEN_NR2_S_0P5 U1259 ( .A1(n580), .A2(A[3]), .X(n582) );
  SEN_OR3B_0P5 U1260 ( .B1(n510), .B2(INST[0]), .A(n352), .X(n1289) );
  SEN_ND2_S_0P5 U1261 ( .A1(n1102), .A2(n1101), .X(n1104) );
  SEN_INV_S_0P5 U1262 ( .A(n1116), .X(n1102) );
  SEN_ND3_S_0P5 U1263 ( .A1(n1097), .A2(n1120), .A3(n1096), .X(n1098) );
  SEN_ND2B_S_0P5 U1264 ( .A(n629), .B(n628), .X(n630) );
  SEN_INV_S_0P5 U1267 ( .A(n625), .X(n626) );
  SEN_AN3_0P5 U1268 ( .A1(INST[2]), .A2(INST[0]), .A3(n352), .X(n355) );
  SEN_OR2_DG_1 U1269 ( .A1(n268), .A2(B[28]), .X(n1236) );
  SEN_NR2_S_0P5 U1270 ( .A1(n417), .A2(n1246), .X(n413) );
  SEN_ND2_S_0P5 U1271 ( .A1(n268), .A2(B[28]), .X(n1230) );
  SEN_ND2_S_0P5 U1273 ( .A1(n1120), .A2(n497), .X(n429) );
  SEN_ND2B_S_0P5 U1274 ( .A(n386), .B(A[29]), .X(n1250) );
  SEN_ND2B_S_0P5 U1275 ( .A(A[25]), .B(B[25]), .X(n485) );
  SEN_INV_S_0P5 U1276 ( .A(INST[2]), .X(n510) );
  SEN_ND3_S_0P5 U1277 ( .A1(n794), .A2(n793), .A3(n792), .X(Z[12]) );
  SEN_MUXI2_S_0P5 U1278 ( .D0(n791), .D1(n790), .S(A[12]), .X(n792) );
  SEN_MUXI2_S_0P5 U1279 ( .D0(n785), .D1(n784), .S(n783), .X(n794) );
  SEN_ND3_S_0P5 U1280 ( .A1(n882), .A2(n881), .A3(n880), .X(Z[16]) );
  SEN_ND2_S_0P5 U1281 ( .A1(B[16]), .A2(n297), .X(n881) );
  SEN_MUXI2_S_0P5 U1282 ( .D0(n879), .D1(n878), .S(A[16]), .X(n880) );
  SEN_ND3_S_0P5 U1283 ( .A1(n690), .A2(n689), .A3(n688), .X(Z[8]) );
  SEN_MUXI2_S_0P5 U1284 ( .D0(n687), .D1(n686), .S(A[8]), .X(n688) );
  SEN_MUXI2_S_0P5 U1285 ( .D0(n680), .D1(n679), .S(n678), .X(n690) );
  SEN_ND3_S_0P5 U1286 ( .A1(n655), .A2(n654), .A3(n653), .X(Z[6]) );
  SEN_ND2_S_0P5 U1287 ( .A1(B[6]), .A2(n1304), .X(n654) );
  SEN_MUXI2_S_0P5 U1288 ( .D0(n646), .D1(n645), .S(n644), .X(n655) );
  SEN_MUXI2_S_0P5 U1289 ( .D0(n652), .D1(n651), .S(A[6]), .X(n653) );
  SEN_MUXI2_S_0P5 U1290 ( .D0(n946), .D1(n945), .S(A[18]), .X(n947) );
  SEN_INV_S_0P5 U1291 ( .A(B[25]), .X(n1146) );
  SEN_INV_S_0P5 U1292 ( .A(B[27]), .X(n1185) );
  SEN_NR2_S_0P5 U1293 ( .A1(n1251), .A2(n1264), .X(n1253) );
  SEN_OR3B_0P5 U1294 ( .B1(n528), .B2(INST[1]), .A(n351), .X(n1291) );
  SEN_OR3B_0P5 U1295 ( .B1(n514), .B2(INST[2]), .A(n352), .X(n1293) );
  SEN_ND2_S_0P5 U1296 ( .A1(n669), .A2(n668), .X(n670) );
  SEN_NR2_S_0P5 U1297 ( .A1(n666), .A2(n298), .X(n669) );
  SEN_MUXI2_S_0P5 U1298 ( .D0(n667), .D1(n1298), .S(B[7]), .X(n668) );
  SEN_INV_S_0P5 U1299 ( .A(n685), .X(n666) );
  SEN_AOI21_S_0P5 U1300 ( .A1(n545), .A2(n389), .B(n298), .X(n539) );
  SEN_MUXI2_S_0P5 U1301 ( .D0(n537), .D1(n1298), .S(B[1]), .X(n538) );
  SEN_INV_0P5 U1302 ( .A(n943), .X(n903) );
  SEN_ND2_S_0P5 U1303 ( .A1(n751), .A2(n750), .X(n752) );
  SEN_NR2_S_0P5 U1304 ( .A1(n247), .A2(n298), .X(n751) );
  SEN_NR3_0P5 U1305 ( .A1(n526), .A2(n525), .A3(n524), .X(n527) );
  SEN_NR2_S_0P5 U1306 ( .A1(n530), .A2(n523), .X(n524) );
  SEN_INV_S_0P5 U1307 ( .A(n941), .X(n901) );
  SEN_ND2_S_0P5 U1308 ( .A1(n786), .A2(n748), .X(n753) );
  SEN_ND3_S_0P5 U1309 ( .A1(n1022), .A2(n1021), .A3(n1020), .X(Z[20]) );
  SEN_ND2_S_0P5 U1310 ( .A1(B[20]), .A2(n1304), .X(n1020) );
  SEN_MUXI2_S_0P5 U1311 ( .D0(n986), .D1(n985), .S(A[20]), .X(n1022) );
  SEN_ND3_S_0P5 U1312 ( .A1(n559), .A2(n558), .A3(n557), .X(Z[2]) );
  SEN_ND2_S_0P5 U1313 ( .A1(B[2]), .A2(n1304), .X(n557) );
  SEN_MUXI2_S_0P5 U1314 ( .D0(n556), .D1(n555), .S(n288), .X(n558) );
  SEN_MUXI2_S_0P5 U1315 ( .D0(n549), .D1(n548), .S(n241), .X(n559) );
  SEN_ND2B_S_0P5 U1316 ( .A(n572), .B(n571), .X(n573) );
  SEN_ND2_S_0P5 U1317 ( .A1(n343), .A2(n1085), .X(n1089) );
  SEN_ND2_S_0P5 U1318 ( .A1(n971), .A2(n982), .X(n986) );
  SEN_ND2B_S_0P5 U1319 ( .A(n386), .B(A[19]), .X(n982) );
  SEN_ND2_S_0P5 U1320 ( .A1(n579), .A2(n578), .X(n584) );
  SEN_ND2_S_0P5 U1321 ( .A1(A[3]), .A2(n388), .X(n579) );
  SEN_ND2_S_0P5 U1322 ( .A1(n648), .A2(n647), .X(n652) );
  SEN_ND2_S_0P5 U1323 ( .A1(A[5]), .A2(n388), .X(n648) );
  SEN_ND2_S_0P5 U1324 ( .A1(n724), .A2(n723), .X(n727) );
  SEN_ND2_S_0P5 U1325 ( .A1(A[9]), .A2(n388), .X(n724) );
  SEN_ND2_S_0P5 U1326 ( .A1(A[13]), .A2(n388), .X(n825) );
  SEN_ND2_S_0P5 U1327 ( .A1(A[25]), .A2(n388), .X(n1156) );
  SEN_ND2_S_0P5 U1328 ( .A1(A[27]), .A2(n389), .X(n1198) );
  SEN_ND2_S_0P5 U1329 ( .A1(A[7]), .A2(n388), .X(n683) );
  SEN_INV_S_0P5 U1330 ( .A(n681), .X(n682) );
  SEN_ND2_S_0P5 U1331 ( .A1(A[11]), .A2(n388), .X(n787) );
  SEN_ND2_S_0P5 U1332 ( .A1(A[15]), .A2(n388), .X(n875) );
  SEN_ND2_S_0P5 U1333 ( .A1(A[17]), .A2(n388), .X(n942) );
  SEN_MUXI2_S_0P5 U1335 ( .D0(n809), .D1(n808), .S(A[13]), .X(n812) );
  SEN_ND2_S_0P5 U1336 ( .A1(n634), .A2(n633), .X(Z[5]) );
  SEN_AOAI211_0P5 U1337 ( .A1(A[5]), .A2(n632), .B(n1304), .C(B[5]), .X(n633)
         );
  SEN_MUXI2_S_0P5 U1338 ( .D0(n631), .D1(n630), .S(A[5]), .X(n634) );
  SEN_ND2_S_0P5 U1339 ( .A1(n647), .A2(n624), .X(n631) );
  SEN_ND2_S_0P5 U1340 ( .A1(n577), .A2(n576), .X(Z[3]) );
  SEN_AOAI211_0P5 U1341 ( .A1(A[3]), .A2(n575), .B(n1304), .C(B[3]), .X(n576)
         );
  SEN_MUXI2_S_0P5 U1342 ( .D0(n574), .D1(n573), .S(A[3]), .X(n577) );
  SEN_ND2_S_0P5 U1343 ( .A1(n578), .A2(n569), .X(n574) );
  SEN_MUXI2_S_0P5 U1345 ( .D0(n705), .D1(n704), .S(A[9]), .X(n708) );
  SEN_ND2_S_0P5 U1346 ( .A1(n723), .A2(n698), .X(n705) );
  SEN_INV_S_0P5 U1347 ( .A(B[30]), .X(n1264) );
  SEN_INV_S_0P5 U1348 ( .A(B[26]), .X(n1167) );
  SEN_INV_S_0P5 U1349 ( .A(B[22]), .X(n1060) );
  SEN_ND2B_S_0P5 U1350 ( .A(B[31]), .B(A[31]), .X(n497) );
  SEN_ND2B_S_0P5 U1351 ( .A(A[26]), .B(B[26]), .X(n487) );
  SEN_OAI211_0P5 U1352 ( .A1(n513), .A2(n216), .B1(n512), .B2(n511), .X(n526)
         );
  SEN_EN2_0P5 U1353 ( .A1(B[0]), .A2(SEL), .X(n513) );
  SEN_ND2B_S_0P5 U1354 ( .A(n1251), .B(n550), .X(n511) );
  SEN_ND2_S_0P5 U1355 ( .A1(n533), .A2(n518), .X(n512) );
  SEN_ND2_S_0P5 U1356 ( .A1(A[30]), .A2(B[30]), .X(n1271) );
  SEN_OAI211_0P5 U1357 ( .A1(n354), .A2(n1060), .B1(n1059), .B2(n1058), .X(
        Z[22]) );
  SEN_OR3B_0P5 U1358 ( .B1(n522), .B2(INST[3]), .A(n521), .X(n530) );
  SEN_EN2_0P5 U1359 ( .A1(INST[0]), .A2(n520), .X(n521) );
  SEN_ND2_S_0P5 U1360 ( .A1(INST[2]), .A2(SEL), .X(n520) );
  SEN_ND2B_S_0P5 U1361 ( .A(SEL), .B(INST[2]), .X(n515) );
  SEN_MUXI2_S_0P5 U1362 ( .D0(n828), .D1(n827), .S(A[14]), .X(n829) );
  SEN_MUXI2_S_0P5 U1363 ( .D0(n823), .D1(n822), .S(n821), .X(n830) );
  SEN_MUXI2_S_0P5 U1364 ( .D0(n727), .D1(n726), .S(A[10]), .X(n728) );
  SEN_MUXI2_S_0P5 U1365 ( .D0(n722), .D1(n721), .S(n720), .X(n729) );
  SEN_AOAI211_0P5 U1366 ( .A1(n739), .A2(n712), .B(n734), .C(n289), .X(n717)
         );
  SEN_INV_S_0P5 U1367 ( .A(n309), .X(n1107) );
  SEN_OAI211_0P5 U1368 ( .A1(n309), .A2(n270), .B1(n375), .B2(n1103), .X(n1110) );
  SEN_NR2_0P5 U263 ( .A1(n991), .A2(n938), .X(n476) );
  SEN_ND2_0P5 U264 ( .A1(n591), .A2(n592), .X(n554) );
  SEN_AOAI211_G_0P5 U270 ( .A1(A[13]), .A2(n810), .B(n1304), .C(n263), .X(n811) );
  SEN_OR3B_2 U271 ( .B1(A[13]), .B2(A[14]), .A(n839), .X(n840) );
  SEN_ND2_T_1 U273 ( .A1(n1188), .A2(n1187), .X(n340) );
  SEN_ND3_S_1 U274 ( .A1(n885), .A2(n884), .A3(n883), .X(n913) );
  SEN_AOAI211_1 U275 ( .A1(n354), .A2(n1228), .B(n1227), .C(n1226), .X(Z[29])
         );
  SEN_AN3B_0P5 U276 ( .B1(n955), .B2(n956), .A(n954), .X(n958) );
  SEN_NR2_S_2 U278 ( .A1(n954), .A2(n831), .X(n835) );
  SEN_OR2_1P5 U285 ( .A1(n337), .A2(n338), .X(n734) );
  SEN_OAI211_1 U286 ( .A1(n944), .A2(n354), .B1(n948), .B2(n947), .X(Z[18]) );
  SEN_BUF_1 U287 ( .A(n733), .X(n1308) );
  SEN_ND2_T_1P5 U288 ( .A1(n757), .A2(n759), .X(n733) );
  SEN_OR3B_1 U289 ( .B1(n903), .B2(n298), .A(n905), .X(n906) );
  SEN_MUXI2_DG_1 U292 ( .D0(n904), .D1(n1298), .S(B[17]), .X(n905) );
  SEN_MUXI2_D_1 U293 ( .D0(n899), .D1(n904), .S(B[17]), .X(n900) );
  SEN_ND2B_S_4 U297 ( .A(n1309), .B(n635), .X(n656) );
  SEN_AN2_DG_16 U298 ( .A1(B[5]), .A2(A[5]), .X(n1309) );
  SEN_ND3_T_0P65 U300 ( .A1(n457), .A2(n456), .A3(n455), .X(n465) );
  SEN_AOAI211_2 U301 ( .A1(n858), .A2(n884), .B(n857), .C(n290), .X(n915) );
  SEN_ND2_S_4 U303 ( .A1(n280), .A2(n281), .X(n1224) );
  SEN_INV_S_1P5 U304 ( .A(n805), .X(n839) );
  SEN_OR3B_2 U306 ( .B1(A[11]), .B2(A[12]), .A(n795), .X(n805) );
  SEN_INV_S_1P5 U308 ( .A(n950), .X(n1023) );
  SEN_MUXI2_DG_0P75 U309 ( .D0(n1294), .D1(n1255), .S(A[30]), .X(n1257) );
  SEN_MUXI2_DG_1 U310 ( .D0(n804), .D1(n296), .S(n263), .X(n807) );
  SEN_INV_0P8 U311 ( .A(n799), .X(n800) );
  SEN_ND2B_V1DG_1 U313 ( .A(n241), .B(B[2]), .X(n592) );
  SEN_INV_S_0P5 U315 ( .A(n293), .X(n1310) );
  SEN_INV_S_0P5 U320 ( .A(n657), .X(n1311) );
  SEN_INV_S_0P5 U328 ( .A(n1311), .X(n1312) );
  SEN_INV_S_0P5 U329 ( .A(n639), .X(n1313) );
  SEN_AOAI211_2 U330 ( .A1(n621), .A2(n620), .B(n619), .C(n618), .X(n623) );
  SEN_NR2_S_4 U333 ( .A1(n312), .A2(n999), .X(n1013) );
  SEN_ND2_T_1P5 U335 ( .A1(n1178), .A2(n1185), .X(n330) );
  SEN_BUF_1 U342 ( .A(n987), .X(n1314) );
  SEN_ND2_4 U348 ( .A1(n993), .A2(n987), .X(n1123) );
  SEN_AO21_2 U349 ( .A1(n560), .A2(n551), .B(n532), .X(n611) );
  SEN_ND2_S_0P5 U350 ( .A1(A[0]), .A2(B[0]), .X(n532) );
  SEN_AOAI211_G_4 U352 ( .A1(n1186), .A2(n1267), .B(n1229), .C(n1231), .X(
        n1190) );
  SEN_ND2_S_0P8 U353 ( .A1(n591), .A2(n590), .X(n614) );
  SEN_NR2_T_1P5 U355 ( .A1(n614), .A2(n613), .X(n621) );
  SEN_OAI22_S_1 U356 ( .A1(n798), .A2(n370), .B1(n799), .B2(n378), .X(n810) );
  SEN_MUX2_6 U357 ( .D0(n972), .D1(n295), .S(B[19]), .X(n975) );
  SEN_AOAI211_0P75 U359 ( .A1(n354), .A2(n851), .B(n853), .C(n850), .X(Z[15])
         );
  SEN_AOAI211_G_3 U360 ( .A1(n612), .A2(n611), .B(n610), .C(n609), .X(n325) );
  SEN_ND2_2 U361 ( .A1(n325), .A2(n329), .X(n635) );
  SEN_OR2_1 U362 ( .A1(n1244), .A2(n271), .X(n326) );
  SEN_NR3_1 U363 ( .A1(n962), .A2(n990), .A3(n961), .X(n965) );
  SEN_ND2B_V1DG_1 U368 ( .A(n807), .B(n806), .X(n808) );
  SEN_INV_0P8 U370 ( .A(n803), .X(n804) );
  SEN_OAI221_1 U373 ( .A1(n568), .A2(n370), .B1(n567), .B2(n378), .C(n374), 
        .X(n570) );
  SEN_INV_0P5 U375 ( .A(n1291), .X(n384) );
  SEN_ND2_G_4 U376 ( .A1(n1295), .A2(n282), .X(n1303) );
  SEN_MUXI2_DG_0P75 U377 ( .D0(n626), .D1(n296), .S(B[5]), .X(n629) );
  SEN_AO21B_2 U379 ( .A1(n1016), .A2(n1122), .B(n1042), .X(n1028) );
  SEN_ND2_S_1 U381 ( .A1(n1041), .A2(n1069), .X(n1016) );
  SEN_ND2_S_0P65 U382 ( .A1(n1121), .A2(n1123), .X(n1099) );
  SEN_AOAI211_3 U383 ( .A1(n865), .A2(n864), .B(n863), .C(n862), .X(n925) );
  SEN_OAI21_G_1 U384 ( .A1(n346), .A2(n1095), .B(n1094), .X(n1116) );
  SEN_AOAI211_G_3 U385 ( .A1(n1238), .A2(n1237), .B(n1259), .C(n1273), .X(
        n1244) );
  SEN_OR2_1 U386 ( .A1(A[14]), .A2(B[14]), .X(n856) );
  SEN_INV_4 U387 ( .A(n760), .X(n762) );
  SEN_ND2B_V1_1 U389 ( .A(A[9]), .B(B[9]), .X(n715) );
  SEN_OAI21_2 U390 ( .A1(n797), .A2(n864), .B(n989), .X(n799) );
  SEN_INV_0P65 U392 ( .A(n781), .X(n797) );
  SEN_ND2_S_0P65 U393 ( .A1(n989), .A2(n815), .X(n782) );
  SEN_INV_S_0P5 U395 ( .A(n1099), .X(n998) );
  SEN_ND2_T_1 U396 ( .A1(n1240), .A2(n1242), .X(n492) );
  SEN_AO21B_2 U405 ( .A1(n1239), .A2(n1164), .B(n273), .X(n410) );
  SEN_AN2_DG_1 U407 ( .A1(n1194), .A2(n1188), .X(n273) );
  SEN_AO21B_2 U409 ( .A1(n273), .A2(n408), .B(n350), .X(n416) );
  SEN_ND2B_V1DG_1 U410 ( .A(B[28]), .B(n268), .X(n1240) );
  SEN_ND2_T_2 U415 ( .A1(n1012), .A2(n1013), .X(n1062) );
  SEN_AOAI211_G_1 U416 ( .A1(n423), .A2(n422), .B(n421), .C(n420), .X(n437) );
  SEN_AOAI211_0P75 U417 ( .A1(n406), .A2(n405), .B(n404), .C(n893), .X(n423)
         );
  SEN_OAI21_T_3 U418 ( .A1(n1220), .A2(B[29]), .B(n283), .X(n1225) );
  SEN_INV_2 U419 ( .A(n1217), .X(n1220) );
  SEN_ND2_T_4 U421 ( .A1(n1187), .A2(n1188), .X(n1285) );
  SEN_OAI21_S_8 U422 ( .A1(n322), .A2(n991), .B(n964), .X(n987) );
  SEN_OA21_4 U423 ( .A1(n932), .A2(n931), .B(n930), .X(n322) );
  SEN_AO2BB2_4 U424 ( .A1(B[4]), .A2(A[4]), .B1(n608), .B2(n607), .X(n610) );
  SEN_AN2_S_1 U425 ( .A1(A[14]), .A2(B[14]), .X(n269) );
  SEN_MUXI2_S_1 U427 ( .D0(n1155), .D1(n1154), .S(n1153), .X(n1162) );
  SEN_INV_S_4 U437 ( .A(n1000), .X(n311) );
  SEN_BUF_1 U438 ( .A(n918), .X(n1315) );
  SEN_INV_S_1P5 U439 ( .A(n1265), .X(n1209) );
  SEN_AOI211_G_2 U440 ( .A1(n1209), .A2(n1234), .B1(n1208), .B2(n1232), .X(
        n1211) );
  SEN_MUXI2_DG_1 U441 ( .D0(n509), .D1(n508), .S(INST[2]), .X(n529) );
  SEN_OAI21_T_2 U443 ( .A1(n484), .A2(n1117), .B(n483), .X(n491) );
  SEN_OAI21_T_2 U444 ( .A1(n271), .A2(n1193), .B(n1192), .X(n1195) );
  SEN_INV_1 U445 ( .A(n1123), .X(n1125) );
  SEN_OAI21_0P75 U446 ( .A1(n965), .A2(n1314), .B(n993), .X(n967) );
  SEN_AOI21B_1 U447 ( .A1(n373), .A2(n284), .B(n375), .X(n1073) );
  SEN_INV_0P5 U448 ( .A(n298), .X(n299) );
  SEN_AN2_1 U449 ( .A1(n649), .A2(n299), .X(n628) );
  SEN_INV_0P5 U451 ( .A(n1300), .X(n298) );
  SEN_OAI21_S_8 U452 ( .A1(n1213), .A2(n1212), .B(n1240), .X(n1216) );
  SEN_ND2B_V1_2 U456 ( .A(A[21]), .B(B[21]), .X(n1120) );
  SEN_AN2_S_4 U457 ( .A1(n1297), .A2(n1296), .X(n282) );
  SEN_MUXI2_DG_3 U459 ( .D0(n1305), .D1(n1299), .S(B[31]), .X(n1297) );
  SEN_OAI22_T_1 U462 ( .A1(n1288), .A2(n370), .B1(n1287), .B2(n377), .X(n1305)
         );
  SEN_INV_4 U463 ( .A(n1191), .X(n1213) );
  SEN_NR2B_1 U464 ( .A(n713), .B(n265), .X(n353) );
  SEN_AOAI211_G_3 U465 ( .A1(n918), .A2(n919), .B(n917), .C(n916), .X(n957) );
  SEN_OAI21_T_6 U466 ( .A1(B[24]), .A2(A[24]), .B(n1114), .X(n1265) );
  SEN_AOAI211_6 U468 ( .A1(n1093), .A2(n1092), .B(n1091), .C(n1090), .X(n1114)
         );
  SEN_INV_S_4 U469 ( .A(n561), .X(n604) );
  SEN_INV_S_3 U470 ( .A(n743), .X(n795) );
  SEN_OA21B_1 U472 ( .A1(n1170), .A2(n385), .B(n355), .X(n1136) );
  SEN_INV_S_4 U473 ( .A(n1137), .X(n1170) );
  SEN_ND2_S_2 U475 ( .A1(n1307), .A2(n1306), .X(Z[31]) );
  SEN_ND2_0P8 U477 ( .A1(n710), .A2(n709), .X(n736) );
  SEN_ND2_S_0P8 U478 ( .A1(B[7]), .A2(A[7]), .X(n710) );
  SEN_ND2_0P5 U483 ( .A1(n710), .A2(n739), .X(n692) );
  SEN_AO21B_2 U484 ( .A1(n796), .A2(n854), .B(n885), .X(n801) );
  SEN_MUXI2_DG_1 U485 ( .D0(n978), .D1(n972), .S(B[19]), .X(n970) );
  SEN_OAI22_S_1 U488 ( .A1(n966), .A2(n270), .B1(n967), .B2(n378), .X(n978) );
  SEN_ND2_0P65 U489 ( .A1(n593), .A2(n592), .X(n617) );
  SEN_ND2B_V1DG_1 U491 ( .A(A[3]), .B(B[3]), .X(n593) );
  SEN_ND2_0P8 U496 ( .A1(n764), .A2(n768), .X(n674) );
  SEN_ND2_S_0P8 U497 ( .A1(n383), .A2(n695), .X(n696) );
  SEN_OAI21_G_0P5 U500 ( .A1(n694), .A2(n693), .B(n713), .X(n695) );
  SEN_AOAI211_3 U502 ( .A1(n496), .A2(n495), .B(n494), .C(n493), .X(n499) );
  SEN_AOAI211_3 U503 ( .A1(n491), .A2(n490), .B(n489), .C(n488), .X(n496) );
  SEN_OR2_2P5 U504 ( .A1(n302), .A2(n303), .X(n608) );
  SEN_INV_S_2 U505 ( .A(n588), .X(n303) );
  SEN_OAI21_T_2 U510 ( .A1(n1211), .A2(n1210), .B(n1230), .X(n1214) );
  SEN_MUXI2_DG_3 U511 ( .D0(n1143), .D1(n1142), .S(A[25]), .X(n1144) );
  SEN_ND2_T_1 U512 ( .A1(n1136), .A2(n1135), .X(n1143) );
  SEN_ND2_2 U513 ( .A1(n1141), .A2(n1140), .X(n1142) );
  SEN_ND3_T_2 U515 ( .A1(n326), .A2(n327), .A3(n374), .X(n1249) );
  SEN_OR2_1P5 U516 ( .A1(n780), .A2(n779), .X(n1009) );
  SEN_OAI21_3 U519 ( .A1(B[6]), .A2(A[6]), .B(n656), .X(n779) );
  SEN_OR2_1P5 U525 ( .A1(n780), .A2(n779), .X(n274) );
  SEN_ND2_S_1P5 U528 ( .A1(n776), .A2(n779), .X(n676) );
  SEN_NR3B_3 U532 ( .A(n1064), .B1(n1062), .B2(n1061), .X(n1063) );
  SEN_OAI21_G_1 U537 ( .A1(n1147), .A2(n270), .B(n1130), .X(n1134) );
  SEN_OR3B_2 U540 ( .B1(A[3]), .B2(A[4]), .A(n604), .X(n627) );
  SEN_INV_S_3 U541 ( .A(n701), .X(n742) );
  SEN_INV_S_6 U548 ( .A(n840), .X(n896) );
  SEN_OAI221_1 U549 ( .A1(n296), .A2(n1167), .B1(n1157), .B2(A[25]), .C(n299), 
        .X(n1158) );
  SEN_ND2_T_0P5 U550 ( .A1(n307), .A2(n308), .X(n706) );
  SEN_ND2_G_1 U553 ( .A1(n697), .A2(n696), .X(n699) );
  SEN_ND2_T_2 U554 ( .A1(n658), .A2(n657), .X(n768) );
  SEN_ND2_S_4 U558 ( .A1(n328), .A2(n637), .X(n657) );
  SEN_INV_S_0P5 U585 ( .A(n384), .X(n378) );
  SEN_AOAI211_0P5 U612 ( .A1(n398), .A2(n399), .B(n397), .C(n396), .X(n403) );
  SEN_INV_S_0P5 U626 ( .A(n854), .X(n858) );
  SEN_ND2_0P5 U630 ( .A1(n856), .A2(n855), .X(n857) );
  SEN_ND2_G_1 U642 ( .A1(n676), .A2(n772), .X(n739) );
  SEN_ND2_0P65 U654 ( .A1(n771), .A2(n275), .X(n775) );
  SEN_OR2_DG_1 U666 ( .A1(n898), .A2(n270), .X(n313) );
  SEN_ND3_T_0P5 U671 ( .A1(n516), .A2(n528), .A3(INST[1]), .X(n1300) );
  SEN_AOAI211_0P5 U676 ( .A1(n590), .A2(n391), .B(n288), .C(n390), .X(n395) );
  SEN_AOI211_0P75 U690 ( .A1(n463), .A2(n462), .B1(n461), .B2(n460), .X(n464)
         );
  SEN_AOAI211_0P5 U692 ( .A1(n476), .A2(n475), .B(n474), .C(n473), .X(n478) );
  SEN_INV_S_0P5 U695 ( .A(n431), .X(n433) );
  SEN_ND2_S_0P5 U700 ( .A1(n241), .A2(B[2]), .X(n585) );
  SEN_OR2_DG_1 U708 ( .A1(n241), .A2(B[2]), .X(n588) );
  SEN_ND2B_V1DG_1 U711 ( .A(B[3]), .B(A[3]), .X(n616) );
  SEN_ND2B_S_0P5 U713 ( .A(A[4]), .B(B[4]), .X(n615) );
  SEN_NR2_S_0P5 U714 ( .A1(A[3]), .A2(B[3]), .X(n302) );
  SEN_ND2B_S_0P5 U715 ( .A(A[6]), .B(B[6]), .X(n658) );
  SEN_ND2B_S_0P5 U716 ( .A(B[8]), .B(A[8]), .X(n713) );
  SEN_ND2B_S_0P5 U718 ( .A(A[10]), .B(B[10]), .X(n757) );
  SEN_ND2B_S_0P5 U720 ( .A(B[12]), .B(A[12]), .X(n989) );
  SEN_ND2B_S_2 U724 ( .A(n768), .B(n769), .X(n995) );
  SEN_INV_S_1 U726 ( .A(n1072), .X(n1131) );
  SEN_ND2B_V1DG_1 U728 ( .A(A[27]), .B(B[27]), .X(n1188) );
  SEN_INV_S_0P5 U729 ( .A(INST[0]), .X(n514) );
  SEN_INV_S_0P5 U732 ( .A(n532), .X(n550) );
  SEN_ND2_S_0P5 U734 ( .A1(n590), .A2(n620), .X(n563) );
  SEN_ND2_S_0P5 U735 ( .A1(n618), .A2(n615), .X(n450) );
  SEN_OAI221_0P5 U736 ( .A1(n325), .A2(n270), .B1(n639), .B2(n378), .C(n374), 
        .X(n625) );
  SEN_ND2_S_0P5 U737 ( .A1(n764), .A2(n658), .X(n643) );
  SEN_INV_S_0P5 U739 ( .A(n677), .X(n694) );
  SEN_ND2_0P5 U741 ( .A1(n766), .A2(n757), .X(n719) );
  SEN_INV_S_0P5 U743 ( .A(n744), .X(n745) );
  SEN_OAI21_G_0P5 U744 ( .A1(n859), .A2(n886), .B(n952), .X(n868) );
  SEN_OAI21_S_0P5 U745 ( .A1(n920), .A2(n277), .B(n1007), .X(n937) );
  SEN_ND2B_V1DG_1 U746 ( .A(A[20]), .B(B[20]), .X(n1122) );
  SEN_INV_S_1 U749 ( .A(n1032), .X(n1071) );
  SEN_INV_S_0P5 U751 ( .A(n384), .X(n379) );
  SEN_INV_0P65 U754 ( .A(n1233), .X(n1147) );
  SEN_ND2_S_0P5 U758 ( .A1(n1164), .A2(n487), .X(n486) );
  SEN_MUXI2_S_0P5 U759 ( .D0(n1219), .D1(n519), .S(A[0]), .X(n525) );
  SEN_INV_S_0P5 U763 ( .A(n450), .X(n598) );
  SEN_ND2_S_0P5 U766 ( .A1(n237), .A2(n310), .X(n844) );
  SEN_MUXI2_D_1 U770 ( .D0(n844), .D1(n846), .S(B[15]), .X(n845) );
  SEN_ND2_S_0P5 U777 ( .A1(n993), .A2(n964), .X(n938) );
  SEN_INV_S_0P5 U782 ( .A(n389), .X(n385) );
  SEN_MUXI2_S_0P5 U784 ( .D0(n1078), .D1(n1298), .S(B[23]), .X(n1079) );
  SEN_NR2_S_0P5 U786 ( .A1(n1177), .A2(n298), .X(n1179) );
  SEN_INV_0P5 U792 ( .A(n1200), .X(n1177) );
  SEN_MUXI2_S_0P5 U793 ( .D0(n1202), .D1(n1201), .S(n268), .X(n1203) );
  SEN_AOAI211_0P5 U796 ( .A1(n1305), .A2(A[31]), .B(n1304), .C(B[31]), .X(
        n1306) );
  SEN_ND2_0P8 U799 ( .A1(B[13]), .A2(A[13]), .X(n884) );
  SEN_ND2_T_2 U802 ( .A1(n1223), .A2(n1227), .X(n280) );
  SEN_ND2_S_0P65 U804 ( .A1(n708), .A2(n707), .X(Z[9]) );
  SEN_OR2_DG_1 U808 ( .A1(n344), .A2(n370), .X(n307) );
  SEN_ND3_T_3 U811 ( .A1(n995), .A2(n994), .A3(n276), .X(n1124) );
  SEN_NR2_T_2 U813 ( .A1(n929), .A2(n928), .X(n932) );
  SEN_INV_S_2 U814 ( .A(n492), .X(n1194) );
  SEN_AN4B_0P5 U816 ( .B1(n861), .B2(n926), .B3(n447), .A(n446), .X(n481) );
  SEN_AOAI211_0P75 U817 ( .A1(n1285), .A2(n1281), .B(n1277), .C(n1282), .X(
        n1245) );
  SEN_INV_1 U818 ( .A(n813), .X(n883) );
  SEN_ND2B_1 U821 ( .A(n1008), .B(n1001), .X(n813) );
  SEN_OAI21_S_8 U823 ( .A1(n341), .A2(n1165), .B(n1164), .X(n1187) );
  SEN_MUXI2_DG_0P75 U824 ( .D0(n753), .D1(n752), .S(A[11]), .X(n754) );
  SEN_MUXI2_DG_1 U826 ( .D0(n502), .D1(n501), .S(INST[0]), .X(n509) );
  SEN_MUXI2_DG_1 U827 ( .D0(n504), .D1(n500), .S(INST[1]), .X(n501) );
  SEN_OAI21_S_3 U828 ( .A1(n340), .A2(n1286), .B(n1284), .X(n1287) );
  SEN_ND2B_1 U830 ( .A(A[13]), .B(B[13]), .X(n860) );
  SEN_ND2_2 U833 ( .A1(n766), .A2(n765), .X(n760) );
  SEN_OAI221_2 U835 ( .A1(n801), .A2(n271), .B1(n800), .B2(n379), .C(n374), 
        .X(n803) );
  SEN_AN2_DG_1 U836 ( .A1(n997), .A2(n996), .X(n276) );
  SEN_MUXI2_S_1 U839 ( .D0(n1036), .D1(n1035), .S(A[21]), .X(n1039) );
  SEN_ND2_S_1 U841 ( .A1(n236), .A2(n1030), .X(n1036) );
  SEN_ND2_0P65 U845 ( .A1(n998), .A2(n1124), .X(n1069) );
  SEN_AN2_S_0P5 U850 ( .A1(B[22]), .A2(A[22]), .X(n1316) );
  SEN_AN2_S_0P5 U860 ( .A1(n1065), .A2(n1064), .X(n1317) );
  SEN_NR3_G_3 U862 ( .A1(n1316), .A2(n1317), .A3(n1063), .X(n1091) );
  SEN_BUF_S_1 U868 ( .A(n1091), .X(n284) );
  SEN_AOAI211_2 U870 ( .A1(n354), .A2(n1183), .B(n1185), .C(n1182), .X(Z[27])
         );
  SEN_MUXI2_S_3 U873 ( .D0(n1181), .D1(n1180), .S(A[27]), .X(n1182) );
  SEN_ND2_G_1 U874 ( .A1(n384), .A2(n301), .X(n1172) );
  SEN_INV_0P8 U877 ( .A(n959), .X(n924) );
  SEN_MUXI2_D_1 U885 ( .D0(n507), .D1(n506), .S(n505), .X(n508) );
  SEN_AOAI211_3 U893 ( .A1(n1278), .A2(n499), .B(n498), .C(n497), .X(n504) );
  SEN_OAI221_0P5 U895 ( .A1(n746), .A2(n370), .B1(n745), .B2(n378), .C(n374), 
        .X(n749) );
  SEN_NR2_0P8 U902 ( .A1(n1026), .A2(n370), .X(n1027) );
  SEN_INV_0P65 U903 ( .A(n272), .X(n370) );
  SEN_AN2_S_1 U904 ( .A1(n351), .A2(n352), .X(n272) );
  SEN_BUF_1P5 U906 ( .A(n272), .X(n373) );
  SEN_INV_0P65 U907 ( .A(n373), .X(n270) );
  SEN_INV_0P8 U912 ( .A(n1293), .X(n389) );
endmodule

