#
# View Description  : LEF layer-definition and P&R technology file
# Stack Description : 6LM HHV stack, M1 + 4 Mx + 0 My + 1 FSG Mz layers
# Target Process    : Common Platform 65nm LP LowK, Doc cmos10lpe.design_manual.pdf, Ver ES46E2339
# Parasitics        : Std Vt
# Pitch, Offset     : X/Y=0.20/0.20, X/Y=0/0
# Date              : 2008/11/18
# Revision          : 1.1.1.3
# Copyright         : 1997-2008 by Virage Logic Corporation
#
VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

UNITS
  DATABASE  MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;
USEMINSPACING OBS OFF ;

PROPERTYDEFINITIONS
  LAYER  LEF57_SPACING STRING ;
  LAYER  LEF57_MINSTEP STRING ;
  LAYER  LEF57_ARRAYSPACING STRING ;
  LAYER  LEF57_ANTENNAGATEPLUSDIFF STRING ;
END PROPERTYDEFINITIONS

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER  PC
  TYPE  MASTERSLICE ;
END PC

LAYER  LVT
  TYPE  implant ;
  SPACING  0.18 ;
  WIDTH  0.18 ;
END LVT

LAYER  HVT
  TYPE  implant ;
  SPACING  0.18 ;
  WIDTH  0.18 ;
END HVT

LAYER  M1
  TYPE  ROUTING ;
  OFFSET  0.00 ;
  AREA  0.042 ;
  WIDTH  0.09 ;
  PITCH  0.20 ;
  SPACINGTABLE  
  PARALLELRUNLENGTH  0.00 0.38 0.42 1.5 4.5
  WIDTH  0.00 0.09 0.09 0.09 0.09 0.09
  WIDTH  0.20 0.09 0.11 0.11 0.11 0.11
  WIDTH  0.42 0.09 0.11 0.16 0.16 0.16
  WIDTH  1.50 0.09 0.11 0.16 0.50 0.50
  WIDTH  4.50 0.09 0.11 0.16 0.50 1.50 ;
  MINIMUMCUT  2 WIDTH 0.345 ;
  MINIMUMCUT  2 WIDTH 0.30 LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT  2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.00 ;
  MINIMUMCUT  2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.00 ;
  MINIMUMCUT  4 WIDTH 0.885 ;
  MINENCLOSEDAREA  0.2 ;
  RESISTANCE  RPERSQ 0.3 ;
  CAPACITANCE  CPERSQDIST 2.0487E-04 ;
  EDGECAPACITANCE  7.0880E-05 ;
  HEIGHT  0.615 ;
  THICKNESS  0.125 ;
  MAXIMUMDENSITY  70 ;
  MINIMUMDENSITY  15 ;
  MAXWIDTH  12 ;
    PROPERTY  LEF57_MINSTEP "MINSTEP 0.09 MAXEDGES 1 ;" ;
  DENSITYCHECKWINDOW  100 100 ;
  DENSITYCHECKSTEP  50 ;
  DIRECTION  HORIZONTAL ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 1000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 300.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ACCURRENTDENSITY  PEAK 3.1650 ;
  ACCURRENTDENSITY  RMS 2.3248 ;
  DCCURRENTDENSITY  AVERAGE 0.1266 ;
  DCCURRENTDENSITY  AVERAGE
  WIDTH  0.12 0.14 0.28 0.32 0.6 0.88 1.16 1.44 2.8 ;
  TABLEENTRIES  0.596 0.613 0.664 0.671 0.692 0.699 0.703 0.706 0.710 ;
END M1

LAYER  V1
  type  CUT ;
  WIDTH  0.10 ;
  SPACING  0.10 ;
  SPACING  0.13 ADJACENTCUTS 3 WITHIN 0.13 ;
  PROPERTY  LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
  PROPERTY  LEF57_ARRAYSPACING "ARRAYSPACING CUTSPACING 0.15 ARRAYCUTS 4 SPACING 0.3 ARRAYCUTS 5 SPACING 0.7 ;" ;
  ENCLOSURE  BELOW 0.02 0.02 WIDTH 0.345 ;
  ENCLOSURE  BELOW 0.03 0.01 ;
  ENCLOSURE  BELOW 0.04 0.00 ;
  ENCLOSURE  ABOVE 0.01 0.01 ;
  ENCLOSURE  ABOVE 0.02 0.01 ;
  ENCLOSURE  ABOVE 0.03 0.00 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 1.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  DCCURRENTDENSITY  AVERAGE 0.0588 ;
END V1

LAYER  M2
  TYPE  ROUTING ;
  OFFSET 0.00 ;
  AREA  0.052 ;
  WIDTH  0.10 ;
  PITCH  0.20 ;
  SPACINGTABLE  
  PARALLELRUNLENGTH  0.00 0.38 0.42 1.5 4.5
  WIDTH  0.00 0.10 0.10 0.10 0.10 0.10
  WIDTH  0.20 0.10 0.12 0.12 0.12 0.12
  WIDTH  0.42 0.10 0.12 0.16 0.16 0.16
  WIDTH  1.50 0.10 0.12 0.16 0.50 0.50
  WIDTH  4.50 0.10 0.12 0.16 0.50 1.50 ;
  MINIMUMCUT  2 WIDTH 0.345 ;
  MINIMUMCUT  2 WIDTH 0.30 LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT  2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.00 ;
  MINIMUMCUT  2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.00 ;
  MINIMUMCUT  4 WIDTH 0.885 ;
  MINENCLOSEDAREA  0.2 ;
  RESISTANCE  RPERSQ 0.2621 ;
  CAPACITANCE  CPERSQDIST 2.2206E-04 ;
  EDGECAPACITANCE  6.4183E-05 ;
  HEIGHT  0.86 ;
  THICKNESS  0.14 ;
  MAXIMUMDENSITY  70 ;
  MINIMUMDENSITY  15 ;
  MAXWIDTH  12 ;
    PROPERTY  LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
  DENSITYCHECKWINDOW  100 100 ;
  DENSITYCHECKSTEP  50 ;
  DIRECTION  HORIZONTAL ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 1000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 300.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ACCURRENTDENSITY  PEAK 3.1650 ;
  ACCURRENTDENSITY  RMS 2.3248 ;
  DCCURRENTDENSITY  AVERAGE 0.1266 ;
  DCCURRENTDENSITY  AVERAGE
  WIDTH  0.12 0.14 0.28 0.32 0.6 0.88 1.16 1.44 2.8 ;
  TABLEENTRIES  0.596 0.613 0.664 0.671 0.692 0.699 0.703 0.706 0.710 ;
END M2

LAYER  V2
  type  CUT ;
  WIDTH  0.10 ;
  SPACING  0.10 ;
  SPACING  0.13 ADJACENTCUTS 3 WITHIN 0.13 ;
  PROPERTY  LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
  PROPERTY  LEF57_ARRAYSPACING "ARRAYSPACING CUTSPACING 0.15 ARRAYCUTS 4 SPACING 0.3 ARRAYCUTS 5 SPACING 0.7 ;" ;
  ENCLOSURE  BELOW 0.02 0.02 WIDTH 0.345 ;
  ENCLOSURE  BELOW 0.03 0.01 ;
  ENCLOSURE  BELOW 0.04 0.00 ;
  ENCLOSURE  ABOVE 0.01 0.01 ;
  ENCLOSURE  ABOVE 0.02 0.01 ;
  ENCLOSURE  ABOVE 0.03 0.00 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 1.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  DCCURRENTDENSITY  AVERAGE 0.0588 ;
END V2

LAYER  M3
  TYPE  ROUTING ;
  OFFSET  0.00 ;
  AREA  0.052 ;
  WIDTH  0.10 ;
  PITCH  0.20 ;
  SPACINGTABLE  
  PARALLELRUNLENGTH  0.00 0.38 0.42 1.5 4.5
  WIDTH  0.00 0.10 0.10 0.10 0.10 0.10
  WIDTH  0.20 0.10 0.12 0.12 0.12 0.12
  WIDTH  0.42 0.10 0.12 0.16 0.16 0.16
  WIDTH  1.50 0.10 0.12 0.16 0.50 0.50
  WIDTH  4.50 0.10 0.12 0.16 0.50 1.50 ;
  MINIMUMCUT  2 WIDTH 0.345 ;
  MINIMUMCUT  2 WIDTH 0.30 LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT  2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.00 ;
  MINIMUMCUT  2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.00 ;
  MINIMUMCUT  4 WIDTH 0.885 ;
  MINENCLOSEDAREA  0.2 ;
  RESISTANCE  RPERSQ 0.2621 ;
  CAPACITANCE  CPERSQDIST 2.2947E-04 ;
  EDGECAPACITANCE  6.4710E-05 ;
  HEIGHT  1.12 ;
  THICKNESS  0.14 ;
  MAXIMUMDENSITY  70 ;
  MINIMUMDENSITY  15 ;
  MAXWIDTH  12 ;
    PROPERTY  LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
  DENSITYCHECKWINDOW  100 100 ;
  DENSITYCHECKSTEP  50 ;
  DIRECTION  VERTICAL ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 1000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 300.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ACCURRENTDENSITY  PEAK 3.1650 ;
  ACCURRENTDENSITY  RMS 2.3248 ;
  DCCURRENTDENSITY  AVERAGE 0.1266 ;
  DCCURRENTDENSITY  AVERAGE
  WIDTH  0.12 0.14 0.28 0.32 0.6 0.88 1.16 1.44 2.8 ;
  TABLEENTRIES  0.596 0.613 0.664 0.671 0.692 0.699 0.703 0.706 0.710 ;
END M3

LAYER  V3
  type  CUT ;
  WIDTH  0.10 ;
  SPACING  0.10 ;
  SPACING  0.13 ADJACENTCUTS 3 WITHIN 0.13 ;
  PROPERTY  LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
  PROPERTY  LEF57_ARRAYSPACING "ARRAYSPACING CUTSPACING 0.15 ARRAYCUTS 4 SPACING 0.3 ARRAYCUTS 5 SPACING 0.7 ;" ;
  ENCLOSURE  BELOW 0.02 0.02 WIDTH 0.345 ;
  ENCLOSURE  BELOW 0.03 0.01 ;
  ENCLOSURE  BELOW 0.04 0.00 ;
  ENCLOSURE  ABOVE 0.01 0.01 ;
  ENCLOSURE  ABOVE 0.02 0.01 ;
  ENCLOSURE  ABOVE 0.03 0.00 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 1.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  DCCURRENTDENSITY  AVERAGE 0.0588 ;
END V3

LAYER  M4
  TYPE  ROUTING ;
  OFFSET  0.00 ;
  AREA  0.052 ;
  WIDTH  0.10 ;
  PITCH  0.20 ;
  SPACINGTABLE  
  PARALLELRUNLENGTH  0.00 0.38 0.42 1.5 4.5
  WIDTH  0.00 0.10 0.10 0.10 0.10 0.10
  WIDTH  0.20 0.10 0.12 0.12 0.12 0.12
  WIDTH  0.42 0.10 0.12 0.16 0.16 0.16
  WIDTH  1.50 0.10 0.12 0.16 0.50 0.50
  WIDTH  4.50 0.10 0.12 0.16 0.50 1.50 ;
  MINIMUMCUT  2 WIDTH 0.345 ;
  MINIMUMCUT  2 WIDTH 0.30 LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT  2 WIDTH 2.00 LENGTH 2.00 WITHIN 2.00 ;
  MINIMUMCUT  2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.00 ;
  MINIMUMCUT  4 WIDTH 0.885 ;
  MINENCLOSEDAREA  0.2 ;
  RESISTANCE  RPERSQ 0.2621 ;
  CAPACITANCE  CPERSQDIST 2.1991E-04 ;
  EDGECAPACITANCE  6.4350E-05 ;
  HEIGHT  1.64 ;
  THICKNESS  0.14 ;
  MAXIMUMDENSITY  70 ;
  MINIMUMDENSITY  15 ;
  MAXWIDTH  12 ;
    PROPERTY  LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
  DENSITYCHECKWINDOW  100 100 ;
  DENSITYCHECKSTEP  50 ;
  DIRECTION  HORIZONTAL ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 1000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 300.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ACCURRENTDENSITY  PEAK 3.1650 ;
  ACCURRENTDENSITY  RMS 2.3248 ;
  DCCURRENTDENSITY  AVERAGE 0.1266 ;
  DCCURRENTDENSITY  AVERAGE
  WIDTH  0.12 0.14 0.28 0.32 0.6 0.88 1.16 1.44 2.8 ;
  TABLEENTRIES  0.596 0.613 0.664 0.671 0.692 0.699 0.703 0.706 0.710 ;
END M4

LAYER  V4
  type  CUT ;
  WIDTH  0.10 ;
  SPACING  0.10 ;
  SPACING  0.13 ADJACENTCUTS 3 WITHIN 0.13 ;
  PROPERTY  LEF57_SPACING "SPACING 0.13 PARALLELOVERLAP ;" ;
  PROPERTY  LEF57_ARRAYSPACING "ARRAYSPACING CUTSPACING 0.15 ARRAYCUTS 4 SPACING 0.3 ARRAYCUTS 5 SPACING 0.7 ;" ;
  ENCLOSURE  BELOW 0.02 0.02 WIDTH 0.345 ;
  ENCLOSURE  BELOW 0.03 0.01 ;
  ENCLOSURE  BELOW 0.04 0.00 ;
  ENCLOSURE  ABOVE 0.01 0.01 ;
  ENCLOSURE  ABOVE 0.02 0.01 ;
  ENCLOSURE  ABOVE 0.03 0.00 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 1.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  DCCURRENTDENSITY  AVERAGE 0.0588 ;
END V4

LAYER  M5
  TYPE  ROUTING ;
  OFFSET  0.00 ;
  AREA  0.052 ;
  WIDTH  0.10 ;
  PITCH  0.20 ;
  SPACINGTABLE  
  PARALLELRUNLENGTH  0.00 0.38 0.42 1.5 4.5
  WIDTH  0.00 0.10 0.10 0.10 0.10 0.10
  WIDTH  0.20 0.10 0.12 0.12 0.12 0.12
  WIDTH  0.42 0.10 0.12 0.16 0.16 0.16
  WIDTH  1.50 0.10 0.12 0.16 0.50 0.50
  WIDTH  4.50 0.10 0.12 0.16 0.50 1.50 ;
  MINIMUMCUT  2 WIDTH 0.345 FROMBELOW ;
  MINIMUMCUT  2 WIDTH 0.30 LENGTH 0.3 WITHIN 0.8 ;
  MINIMUMCUT  2 WIDTH 2.000 LENGTH 2.00 WITHIN 2.00 ;
  MINIMUMCUT  2 WIDTH 3.000 LENGTH 10.0 WITHIN 5.00 ;
  MINIMUMCUT  4 WIDTH 0.885 FROMBELOW ;
  MINIMUMCUT 2  WIDTH 1.800 FROMABOVE ;
  MINENCLOSEDAREA  0.2 ;
  RESISTANCE  RPERSQ 0.2621 ;
  CAPACITANCE  CPERSQDIST 1.4092E-04 ;
  EDGECAPACITANCE  6.7136E-05 ;
  HEIGHT  1.9 ;
  THICKNESS  0.14 ;
  MAXIMUMDENSITY  70 ;
  MINIMUMDENSITY  15 ;
  MAXWIDTH  12 ;
    PROPERTY  LEF57_MINSTEP "MINSTEP 0.10 MAXEDGES 1 ;" ;
  DENSITYCHECKWINDOW  100 100 ;
  DENSITYCHECKSTEP  50 ;
  DIRECTION  VERTICAL ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 1000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 300.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ACCURRENTDENSITY  PEAK 3.1650 ;
  ACCURRENTDENSITY  RMS 2.3248 ;
  DCCURRENTDENSITY  AVERAGE 0.1266 ;
  DCCURRENTDENSITY  AVERAGE
  WIDTH  0.12 0.14 0.28 0.32 0.6 0.88 1.16 1.44 2.8 ;
  TABLEENTRIES  0.596 0.613 0.664 0.671 0.692 0.699 0.703 0.706 0.710 ;
END M5

LAYER  NT
  type  CUT ;
  WIDTH  0.36 ;
  SPACING  0.34 ;
  SPACING  0.54 ADJACENTCUTS 3 WITHIN 0.54 ;
  PROPERTY  LEF57_SPACING
  "SPACING  0.44 PARALLELOVERLAP ;" ;
  ENCLOSURE  0.02 0.02 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 20.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 1.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 5.0 ;" ;
  DCCURRENTDENSITY  AVERAGE 0.4513 ;
END NT

LAYER  EA
  TYPE  ROUTING ;
  OFFSET  0.00 ;
  AREA  0.565 ;
  WIDTH  0.40 ;
  PITCH  0.80 ;
  SPACINGTABLE  
  PARALLELRUNLENGTH  0.00 1.50 4.50
  WIDTH  0.00 0.40 0.40 0.40
  WIDTH  1.50 0.40 0.50 0.50
  WIDTH  4.50 0.40 0.50 1.50 ;
  MINIMUMCUT  2 WIDTH 1.80 ;
  MINIMUMCUT  2 WIDTH 3.00 LENGTH 10.0 WITHIN 5.0 ;
  MINENCLOSEDAREA  0.565 ;
  RESISTANCE  RPERSQ 0.025 ;
  CAPACITANCE  CPERSQDIST 3.2011E-05 ;
  EDGECAPACITANCE  3.9730E-05 ;
  HEIGHT  3.555 ;
  THICKNESS  0.9 ;
  MAXIMUMDENSITY  80 ;
  MINIMUMDENSITY  20 ;
  MAXWIDTH  12.25 ;
    PROPERTY  LEF57_MINSTEP "MINSTEP 0.40 MAXEDGES 1 ;" ;
  DENSITYCHECKWINDOW  100 100 ;
  DENSITYCHECKSTEP  50 ;
  DIRECTION  HORIZONTAL ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFAREARATIO 1000.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ANTENNAMODEL OXIDE2 ;
  ANTENNADIFFAREARATIO 300.0 ;
  PROPERTY LEF57_ANTENNAGATEPLUSDIFF "ANTENNAGATEPLUSDIFF 2.0 ;" ;
  ACCURRENTDENSITY  PEAK 13.01312 ;
  ACCURRENTDENSITY  RMS 3.8888 ;
  DCCURRENTDENSITY  AVERAGE
  WIDTH  0.28 0.56 0.84 1.4 5.0 12.0 ;
  TABLEENTRIES  1.489 1.546 1.565 1.580 1.597 1.601 ;
END EA

VIA  Via1  DEFAULT
  LAYER  M1 ;
  RECT  -0.050 -0.090 0.050 0.090 ;
  LAYER  V1 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M2 ;
  RECT  -0.080 -0.050 0.080 0.050 ;
  RESISTANCE  6.0 ;
END Via1

VIA  Via2  DEFAULT
  LAYER  M2 ;
  RECT  -0.090 -0.050 0.090 0.050 ;
  LAYER  V2 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M3 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via2

VIA  Via3  DEFAULT
  LAYER  M3 ;
  RECT  -0.090 -0.050 0.090 0.050 ;
  LAYER  V3 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M4 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via3

VIA  Via4  DEFAULT
  LAYER  M4 ;
  RECT  -0.090 -0.050 0.090 0.050 ;
  LAYER  V4 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M5 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via4

VIA  Via5  DEFAULT
  LAYER  M5 ;
  RECT  -0.200 -0.200 0.200 0.200 ;
  LAYER  NT ;
  RECT  -0.180 -0.180 0.180 0.180 ;
  LAYER  EA ;
  RECT  -0.200 -0.200 0.200 0.200 ;
  RESISTANCE  0.27 ;
END Via5

VIA  Via1HH  DEFAULT
  LAYER  M1 ;
  RECT  -0.090 -0.050 0.090 0.050 ;
  LAYER  V1 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M2 ;
  RECT  -0.080 -0.050 0.080 0.050 ;
  RESISTANCE  6.0 ;
END Via1HH

VIA  Via1VV  DEFAULT
  LAYER  M1 ;
  RECT  -0.050 -0.090 0.050 0.090 ;
  LAYER  V1 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M2 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via1VV

VIA  Via1HV  DEFAULT
  LAYER  M1 ;
  RECT  -0.090 -0.050 0.090 0.050 ;
  LAYER  V1 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M2 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via1HV

VIA  Via1_2cut_E_HH  DEFAULT
  LAYER  M1 ;
  RECT  -0.090 -0.050 0.290 0.050 ;
  LAYER  V1 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  RECT  0.150 -0.050 0.250 0.050 ;
  LAYER  M2 ;
  RECT  -0.080 -0.050 0.280 0.050 ;
  RESISTANCE  3.0 ;
END Via1_2cut_E_HH

VIA  Via1_2cut_W_HH  DEFAULT
  LAYER  M1 ;
  RECT  -0.290 -0.050 0.090 0.050 ;
  LAYER  V1 ;
  RECT  -0.250 -0.050 -0.150 0.050 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M2 ;
  RECT  -0.280 -0.050 0.080 0.050 ;
  RESISTANCE  3.0 ;
END Via1_2cut_W_HH

VIA  Via1_2cut_N_HH  DEFAULT
  LAYER  M1 ;
  RECT  -0.090 -0.050 0.090 0.250 ;
  LAYER  V1 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  RECT  -0.050 0.150 0.050 0.250 ;
  LAYER  M2 ;
  RECT  -0.080 -0.050 0.080 0.250 ;
  RESISTANCE  3.0 ;
END Via1_2cut_N_HH

VIA  Via1_2cut_S_HH  DEFAULT
  LAYER  M1 ;
  RECT  -0.090 -0.250 0.090 0.050 ;
  LAYER  V1 ;
  RECT  -0.050 -0.250 0.050 -0.150 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M2 ;
  RECT  -0.080 -0.250 0.080 0.050 ;
  RESISTANCE  3.0 ;
END Via1_2cut_S_HH

VIA  Via1_4cut_HH  DEFAULT
  LAYER  M1 ;
  RECT  -0.190 -0.150 0.190 0.150 ;
  LAYER  V1 ;
  RECT  -0.150 -0.150 -0.050 -0.050 ;
  RECT  0.050 -0.150 0.150 -0.050 ;
  RECT  -0.150 0.050 -0.050 0.150 ;
  RECT  0.050 0.050 0.150 0.150 ;
  LAYER  M2 ;
  RECT  -0.180 -0.150 0.180 0.150 ;
  RESISTANCE  1.5 ;
END Via1_4cut_HH

VIA  Via2_MAR_E  DEFAULT
  LAYER  M2 ;
  RECT  -0.090 -0.050 0.430 0.050 ;
  LAYER  V2 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M3 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via2_MAR_E

VIA  Via2_MAR_W  DEFAULT
  LAYER  M2 ;
  RECT  -0.430 -0.050 0.090 0.050 ;
  LAYER  V2 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M3 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via2_MAR_W

VIA  Via2_2cut_E_HV  DEFAULT
  LAYER  M2 ;
  RECT  -0.090 -0.050 0.290 0.050 ;
  LAYER  V2 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  RECT  0.150 -0.050 0.250 0.050 ;
  LAYER  M3 ;
  RECT  -0.050 -0.080 0.250 0.080 ;
  RESISTANCE  3.0 ;
END Via2_2cut_E_HV

VIA  Via2_2cut_W_HV  DEFAULT
  LAYER  M2 ;
  RECT  -0.290 -0.050 0.090 0.050 ;
  LAYER  V2 ;
  RECT  -0.250 -0.050 -0.150 0.050 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M3 ;
  RECT  -0.250 -0.080 0.050 0.080 ;
  RESISTANCE  3.0 ;
END Via2_2cut_W_HV

VIA  Via2_2cut_N_HV  DEFAULT
  LAYER  M2 ;
  RECT  -0.090 -0.050 0.090 0.250 ;
  LAYER  V2 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  RECT  -0.050 0.150 0.050 0.250 ;
  LAYER  M3 ;
  RECT  -0.050 -0.080 0.050 0.280 ;
  RESISTANCE  3.0 ;
END Via2_2cut_N_HV

VIA  Via2_2cut_S_HV  DEFAULT
  LAYER  M2 ;
  RECT  -0.090 -0.250 0.090 0.050 ;
  LAYER  V2 ;
  RECT  -0.050 -0.250 0.050 -0.150 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M3 ;
  RECT  -0.050 -0.280 0.050 0.080 ;
  RESISTANCE  3.0 ;
END Via2_2cut_S_HV

VIA  Via2_4cut_HV  DEFAULT
  LAYER  M2 ;
  RECT  -0.190 -0.150 0.190 0.150 ;
  LAYER  V2 ;
  RECT  -0.150 -0.150 -0.050 -0.050 ;
  RECT  0.050 -0.150 0.150 -0.050 ;
  RECT  -0.150 0.050 -0.050 0.150 ;
  RECT  0.050 0.050 0.150 0.150 ;
  LAYER  M3 ;
  RECT  -0.150 -0.180 0.150 0.180 ;
  RESISTANCE  1.5 ;
END Via2_4cut_HV

VIA  Via3_MAR_E  DEFAULT
  LAYER  M3 ;
  RECT  -0.050 -0.090 0.050 0.430 ;
  LAYER  V3 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M4 ;
  RECT  -0.080 -0.050 0.080 0.050 ;
  RESISTANCE  6.0 ;
END Via3_MAR_E

VIA  Via3_MAR_W  DEFAULT
  LAYER  M3 ;
  RECT  -0.050 -0.430 0.050 0.090 ;
  LAYER  V3 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M4 ;
  RECT  -0.080 -0.050 0.080 0.050 ;
  RESISTANCE  6.0 ;
END Via3_MAR_W

VIA  Via3_2cut_E_HV  DEFAULT
  LAYER  M3 ;
  RECT  -0.050 -0.090 0.050 0.290 ;
  LAYER  V3 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  RECT  -0.050 0.150 0.050 0.250 ;
  LAYER  M4 ;
  RECT  -0.080 -0.050 0.080 0.250 ;
  RESISTANCE  3.0 ;
END Via3_2cut_E_HV

VIA  Via3_2cut_W_HV  DEFAULT
  LAYER  M3 ;
  RECT  -0.050 -0.290 0.050 0.090 ;
  LAYER  V3 ;
  RECT  -0.050 -0.250 0.050 -0.150 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M4 ;
  RECT  -0.080 -0.250 0.080 0.050 ;
  RESISTANCE  3.0 ;
END Via3_2cut_W_HV

VIA  Via3_2cut_N_HV  DEFAULT
  LAYER  M3 ;
  RECT  -0.050 -0.090 0.250 0.090 ;
  LAYER  V3 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  RECT  0.150 -0.050 0.250 0.050 ;
  LAYER  M4 ;
  RECT  -0.080 -0.050 0.280 0.050 ;
  RESISTANCE  3.0 ;
END Via3_2cut_N_HV

VIA  Via3_2cut_S_HV  DEFAULT
  LAYER  M3 ;
  RECT  -0.250 -0.090 0.050 0.090 ;
  LAYER  V3 ;
  RECT  -0.250 -0.050 -0.150 0.050 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M4 ;
  RECT  -0.280 -0.050 0.080 0.050 ;
  RESISTANCE  3.0 ;
END Via3_2cut_S_HV

VIA  Via3_4cut_HV  DEFAULT
  LAYER  M3 ;
  RECT  -0.150 -0.190 0.150 0.190 ;
  LAYER  V3 ;
  RECT  -0.150 -0.150 -0.050 -0.050 ;
  RECT  -0.150 0.050 -0.050 0.150 ;
  RECT  0.050 -0.150 0.150 -0.050 ;
  RECT  0.050 0.050 0.150 0.150 ;
  LAYER  M4 ;
  RECT  -0.180 -0.150 0.180 0.150 ;
  RESISTANCE  1.5 ;
END Via3_4cut_HV

VIA  Via4_MAR_N  DEFAULT
  LAYER  M4 ;
  RECT  -0.090 -0.050 0.430 0.050 ;
  LAYER  V4 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M5 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via4_MAR_N

VIA  Via4_MAR_S  DEFAULT
  LAYER  M4 ;
  RECT  -0.430 -0.050 0.090 0.050 ;
  LAYER  V4 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M5 ;
  RECT  -0.050 -0.080 0.050 0.080 ;
  RESISTANCE  6.0 ;
END Via4_MAR_S

VIA  Via4_2cut_E_VH  DEFAULT
  LAYER  M4 ;
  RECT  -0.090 -0.050 0.090 0.250 ;
  LAYER  V4 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  RECT  -0.050 0.150 0.050 0.250 ;
  LAYER  M5 ;
  RECT  -0.050 -0.080 0.050 0.280 ;
  RESISTANCE  3.0 ;
END Via4_2cut_E_VH

VIA  Via4_2cut_W_VH  DEFAULT
  LAYER  M4 ;
  RECT  -0.090 -0.250 0.090 0.050 ;
  LAYER  V4 ;
  RECT  -0.050 -0.250 0.050 -0.150 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M5 ;
  RECT  -0.050 -0.280 0.050 0.080 ;
  RESISTANCE  3.0 ;
END Via4_2cut_W_VH

VIA  Via4_2cut_N_VH  DEFAULT
  LAYER  M4 ;
  RECT  -0.090 -0.050 0.290 0.050 ;
  LAYER  V4 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  RECT  0.150 -0.050 0.250 0.050 ;
  LAYER  M5 ;
  RECT  -0.050 -0.080 0.250 0.080 ;
  RESISTANCE  3.0 ;
END Via4_2cut_N_VH

VIA  Via4_2cut_S_VH  DEFAULT
  LAYER  M4 ;
  RECT  -0.290 -0.050 0.090 0.050 ;
  LAYER  V4 ;
  RECT  -0.250 -0.050 -0.150 0.050 ;
  RECT  -0.050 -0.050 0.050 0.050 ;
  LAYER  M5 ;
  RECT  -0.250 -0.080 0.050 0.080 ;
  RESISTANCE  3.0 ;
END Via4_2cut_S_VH

VIA  Via4_4cut_VH  DEFAULT
  LAYER  M4 ;
  RECT  -0.190 -0.150 0.190 0.150 ;
  LAYER  V4 ;
  RECT  -0.150 -0.150 -0.050 -0.050 ;
  RECT  -0.150 0.050 -0.050 0.150 ;
  RECT  0.050 -0.150 0.150 -0.050 ;
  RECT  0.050 0.050 0.150 0.150 ;
  LAYER  M5 ;
  RECT  -0.150 -0.180 0.150 0.180 ;
  RESISTANCE  1.5 ;
END Via4_4cut_VH

VIA  Via5_2cut_E_HV  DEFAULT
  LAYER  M5 ;
  RECT  -0.200 -0.200 0.200 0.900 ;
  LAYER  NT ;
  RECT  -0.180 -0.180 0.180 0.180 ;
  RECT  -0.180 0.520 0.180 0.880 ;
  LAYER  EA ;
  RECT  -0.200 -0.200 0.200 0.900 ;
  RESISTANCE  0.135 ;
END Via5_2cut_E_HV

VIA  Via5_2cut_W_HV  DEFAULT
  LAYER  M5 ;
  RECT  -0.200 -0.900 0.200 0.200 ;
  LAYER  NT ;
  RECT  -0.180 -0.880 0.180 -0.520 ;
  RECT  -0.180 -0.180 0.180 0.180 ;
  LAYER  EA ;
  RECT  -0.200 -0.900 0.200 0.200 ;
  RESISTANCE  0.135 ;
END Via5_2cut_W_HV

VIA  Via5_2cut_N_HV  DEFAULT
  LAYER  M5 ;
  RECT  -0.200 -0.200 0.900 0.200 ;
  LAYER  NT ;
  RECT  -0.180 -0.180 0.180 0.180 ;
  RECT  0.520 -0.180 0.880 0.180 ;
  LAYER  EA ;
  RECT  -0.200 -0.200 0.900 0.200 ;
  RESISTANCE  0.135 ;
END Via5_2cut_N_HV

VIA  Via5_2cut_S_HV  DEFAULT
  LAYER  M5 ;
  RECT  -0.900 -0.200 0.200 0.200 ;
  LAYER  NT ;
  RECT  -0.880 -0.180 -0.520 0.180 ;
  RECT  -0.180 -0.180 0.180 0.180 ;
  LAYER  EA ;
  RECT  -0.900 -0.200 0.200 0.200 ;
  RESISTANCE  0.135 ;
END Via5_2cut_S_HV

VIA  Via5_4cut_HV  DEFAULT
  LAYER  M5 ;
  RECT  -0.550 -0.550 0.550 0.550 ;
  LAYER  NT ;
  RECT  -0.530 -0.530 -0.170 -0.170 ;
  RECT  -0.530 0.170 -0.170 0.530 ;
  RECT  0.170 -0.530 0.530 -0.170 ;
  RECT  0.170 0.170 0.530 0.530 ;
  LAYER  EA ;
  RECT  -0.550 -0.550 0.550 0.550 ;
  RESISTANCE  0.068 ;
END Via5_4cut_HV

VIARULE  viagen_V1  GENERATE
  LAYER  M1 ;
  ENCLOSURE  0.04 0.00 ;
  WIDTH  0.09 TO 12 ;
  LAYER  M2 ;
  ENCLOSURE  0.03 0.00 ;
  WIDTH  0.10 TO 12 ;
  LAYER  V1 ;
  RECT  -0.05 -0.05 0.05 0.05 ;
  SPACING  0.20 BY 0.20 ;
END viagen_V1

VIARULE  viagen_V2  GENERATE
  LAYER  M2 ;
  ENCLOSURE  0.04 0.00 ;
  WIDTH  0.10 TO 12 ;
  LAYER  M3 ;
  ENCLOSURE  0.00 0.03 ;
  WIDTH  0.10 TO 12 ;
  LAYER  V2 ;
  RECT  -0.05 -0.05 0.05 0.05 ;
  SPACING  0.20 BY 0.20 ;
END viagen_V2

VIARULE  viagen_V3  GENERATE
  LAYER  M3 ;
  ENCLOSURE  0.00 0.04 ;
  WIDTH  0.10 TO 12 ;
  LAYER  M4 ;
  ENCLOSURE  0.03 0.00 ;
  WIDTH  0.10 TO 12 ;
  LAYER  V3 ;
  RECT  -0.05 -0.05 0.05 0.05 ;
  SPACING  0.20 BY 0.20 ;
END viagen_V3

VIARULE  viagen_V4  GENERATE
  LAYER  M4 ;
  ENCLOSURE  0.04 0.00 ;
  WIDTH  0.10 TO 12 ;
  LAYER  M5 ;
  ENCLOSURE  0.00 0.03 ;
  WIDTH  0.10 TO 12 ;
  LAYER  V4 ;
  RECT  -0.05 -0.05 0.05 0.05 ;
  SPACING  0.20 BY 0.20 ;
END viagen_V4

VIARULE  viagen_NT  GENERATE
  LAYER  M5 ;
  ENCLOSURE  0.02 0.02 ;
  WIDTH  0.20 TO 12 ;
  LAYER  EA ;
  ENCLOSURE  0.02 0.02 ;
  WIDTH  0.40 TO 12.25 ;
  LAYER  NT ;
  RECT  -0.18 -0.18 0.18 0.18 ;
  SPACING  0.70 BY 0.70 ;
END viagen_NT

SPACING
  SAMENET  V1 V2 0.00 STACK ;
  SAMENET  V2 V3 0.00 STACK ;
  SAMENET  V3 V4 0.00 STACK ;
  SAMENET  V4 NT 0.00 STACK ;
  SAMENET  V1 V1 0.10 ;
  SAMENET  V2 V2 0.10 ;
  SAMENET  V3 V3 0.10 ;
  SAMENET  V4 V4 0.10 ;
  SAMENET  NT NT 0.34 ;
END SPACING

END LIBRARY
