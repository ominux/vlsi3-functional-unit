/*
 Top level module for the functional unit of Mosaic

 Author: Corey Olson
 Date: 4/29/2010
*/
module functional_unit();

endmodule
