
module Alu ( Z, A, B, DI, DO, CI, INST, FLAGS, FirstCyc );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [31:0] DI;
  output [31:0] DO;
  input [3:0] INST;
  output [3:0] FLAGS;
  input CI, FirstCyc;
  wire   \*Logic0* , N72, net41954, net58902, net58904, net58908, net58912,
         net58913, net58914, net58915, net58917, net58919, net58921, net58923,
         net58925, net58927, net58929, net58931, net58933, net58935, net58937,
         net58939, net58941, net58943, net58945, net58947, net58949, net58951,
         net58954, net58957, net58960, net58963, net58965, net58967, net58970,
         net58984, net58985, net58986, net58987, net58988, net58989, net59200,
         net59205, net59211, net59212, net59213, net59214, net59215, net59216,
         net59217, net59219, net59221, net59223, net59231, net59232, net59233,
         net59238, net59239, net59240, net59241, net59242, net59249, net59250,
         net59251, net59252, net59255, net59256, net59257, net59258, net59261,
         net59262, net59263, net59264, net59267, net59268, net59270, net59271,
         net59272, net59273, net59274, net59276, net59277, net59278, net59279,
         net59280, net59285, net59286, net59287, net59288, net59290, net59291,
         net59298, net59299, net59300, net59304, net59305, net59306, net59307,
         net59308, net59309, net59310, net59312, net59314, net59315, net59316,
         net59320, net59321, net59322, net59325, net59326, net59327, net59328,
         net59329, net59332, net59333, net59335, net59336, net59337, net59338,
         net59341, net59342, net59343, net59345, net59346, net59347, net59350,
         net59351, net59353, net59356, net59362, net59372, net59374, net59376,
         net59377, net59378, net59380, net59381, net59382, net59385, net59386,
         net59388, net59389, net59390, net59391, net59392, net59393, net59395,
         net59396, net59397, net59398, net59400, net59401, net59402, net59405,
         net59406, net59409, net59410, net59411, net59412, net59413, net59416,
         net59418, net59419, net59421, net59422, net59425, net59426, net59427,
         net59429, net59430, net59431, net59433, net59434, net59437, net59438,
         net59440, net59444, net59454, net59455, net59456, net59457, net59459,
         net59461, net59462, net59463, net59465, net59466, net59469, net59470,
         net59473, net59474, net59482, net59486, net59488, net59490, net59494,
         net59497, net59498, net59500, net59503, net59505, net59513, net59517,
         net59522, net59523, net59530, net59531, net59535, net59536, net59537,
         net59538, net59549, net59558, net59560, net59561, net59562, net59564,
         net59575, net59584, net59593, net59594, net59595, net59596, net59597,
         net59598, net59600, net59601, net59605, net59606, net59608, net59616,
         net59624, net59630, net59631, net59635, net59636, net59637, net59638,
         net59639, net59642, net59651, net59654, net59663, net59666, net59667,
         net59671, net59675, net59677, net59679, net59680, net59686, net59687,
         net59688, net59689, net59690, net59691, net59696, net59700, net59714,
         net59715, net59717, net59725, net59727, net59729, net59730, net59731,
         net59739, net59743, net59744, net59746, net59748, net59754, net59755,
         net59758, net59759, net59760, net59767, net59768, net59769, net59770,
         net59773, net59775, net59777, net59779, net59781, net59792, net59793,
         net59794, net59795, net59798, net59799, net59819, net59849, net59870,
         net59873, net59888, net59966, net59962, net59958, net59980, net59978,
         net59976, net59992, net59990, net59988, net60205, net60219, net60218,
         net60235, net60246, net60361, net60373, net60372, net60376, net60375,
         net60378, net60377, net60381, net60380, net60411, net60418, net60464,
         net60465, net60532, net60540, net60557, net60751, net60861, net60873,
         net60983, net60989, net61215, net61241, net61240, net61246, net61245,
         net61263, net61262, net61305, net61326, net61338, net61773, net61810,
         net61884, net59282, net59237, net61348, net60495, net59633, net59629,
         net59626, net59622, net59621, net59617, net59585, net59583, net59559,
         net59550, net59544, net59543, net59542, net59541, net59533, net59349,
         net59248, net59247, net59750, net59678, net59375, net59370, net61110,
         net59776, net59311, n342, n343, n344, n345, n346, n347, n348, n349,
         \FLAGS[1] , n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n419, n420, n421, n422, n424, n425, n426, n427, n428, n430,
         n431, n432, n433, n434, n435, n436, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n453, n454,
         n455, n456, n458, n459, n460, n461, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n570, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079;
  assign FLAGS[3] = \*Logic0* ;
  assign DO[31] = DI[30];
  assign DO[30] = DI[29];
  assign DO[29] = DI[28];
  assign DO[28] = DI[27];
  assign DO[27] = DI[26];
  assign DO[26] = DI[25];
  assign DO[25] = DI[24];
  assign DO[24] = DI[23];
  assign DO[23] = DI[22];
  assign DO[22] = DI[21];
  assign DO[21] = DI[20];
  assign DO[20] = DI[19];
  assign DO[19] = DI[18];
  assign DO[18] = DI[17];
  assign DO[17] = DI[16];
  assign DO[16] = DI[15];
  assign DO[15] = DI[14];
  assign DO[14] = DI[13];
  assign DO[13] = DI[12];
  assign DO[12] = DI[11];
  assign DO[11] = DI[10];
  assign DO[10] = DI[9];
  assign DO[9] = DI[8];
  assign DO[8] = DI[7];
  assign DO[7] = DI[6];
  assign DO[6] = DI[5];
  assign DO[5] = DI[4];
  assign DO[4] = DI[3];
  assign DO[3] = DI[2];
  assign DO[2] = DI[1];
  assign DO[1] = DI[0];
  assign N72 = INST[0];
  assign FLAGS[2] = net41954;
  assign DO[0] = \FLAGS[1] ;
  assign FLAGS[1] = \FLAGS[1] ;

  SEN_BUF_1 U421 ( .A(n388), .X(n342) );
  SEN_AOI21_T_1P5 U422 ( .A1(n456), .A2(net59819), .B(n463), .X(net59773) );
  SEN_INV_5 U426 ( .A(n424), .X(net59459) );
  SEN_EO2_2 U428 ( .A1(A[10]), .A2(net59978), .X(n713) );
  SEN_AN2_24 U429 ( .A1(n344), .A2(INST[1]), .X(n343) );
  SEN_INV_32 U430 ( .A(N72), .X(n344) );
  SEN_ND3_T_4 U437 ( .A1(n476), .A2(n477), .A3(n478), .X(n345) );
  SEN_ND3_T_4 U438 ( .A1(n476), .A2(n477), .A3(n478), .X(n414) );
  SEN_NR2_S_3 U439 ( .A1(net59746), .A2(net59316), .X(n478) );
  SEN_INV_S_6 U440 ( .A(net59795), .X(net59779) );
  SEN_ND2B_16 U441 ( .A(INST[2]), .B(N72), .X(n346) );
  SEN_NR2_T_2 U442 ( .A1(net59219), .A2(n832), .X(n347) );
  SEN_NR2_4 U443 ( .A1(net59219), .A2(net59221), .X(n348) );
  SEN_INV_S_1P5 U444 ( .A(n831), .X(n349) );
  SEN_ND2_T_3 U447 ( .A1(n766), .A2(n395), .X(n832) );
  SEN_INV_S_6 U448 ( .A(net59482), .X(net59221) );
  SEN_ND2B_1 U449 ( .A(n832), .B(net59482), .X(n831) );
  SEN_INV_2 U452 ( .A(n442), .X(n749) );
  SEN_AOI211_3 U453 ( .A1(n749), .A2(n807), .B1(n747), .B2(n748), .X(n750) );
  SEN_ND2B_S_1 U454 ( .A(net59287), .B(net59291), .X(n732) );
  SEN_INV_8 U455 ( .A(n680), .X(n427) );
  SEN_INV_5 U456 ( .A(net59463), .X(net59474) );
  SEN_EN3_DG_1 U457 ( .A1(net59231), .A2(net59232), .A3(net59233), .X(net58917) );
  SEN_ND3_T_16 U459 ( .A1(n467), .A2(n465), .A3(n466), .X(n464) );
  SEN_ND2_G_3 U460 ( .A1(n406), .A2(n394), .X(n820) );
  SEN_OAI21_G_0P5 U461 ( .A1(net59290), .A2(net59291), .B(n824), .X(n825) );
  SEN_AOAI211_4 U462 ( .A1(n784), .A2(n785), .B(n783), .C(net59486), .X(n790)
         );
  SEN_INV_12 U465 ( .A(n793), .X(n575) );
  SEN_INV_1 U466 ( .A(n793), .X(n795) );
  SEN_MUXI2_S_3 U467 ( .D0(n575), .D1(n716), .S(B[12]), .X(net59715) );
  SEN_OAI21_16 U468 ( .A1(net59205), .A2(INST[1]), .B(N72), .X(n793) );
  SEN_INV_5 U469 ( .A(net59798), .X(n398) );
  SEN_ND2B_16 U474 ( .A(INST[2]), .B(N72), .X(n680) );
  SEN_ND2_G_3 U475 ( .A1(net59888), .A2(n346), .X(n652) );
  SEN_AN2_S_0P5 U476 ( .A1(net59375), .A2(net59374), .X(net60532) );
  SEN_OAI211_4 U478 ( .A1(n647), .A2(n589), .B1(n686), .B2(n649), .X(net59795)
         );
  SEN_ND2_T_4 U481 ( .A1(n361), .A2(net59770), .X(net59688) );
  SEN_AOAI211_6 U482 ( .A1(net59758), .A2(net59759), .B(net59731), .C(n474), 
        .X(net59304) );
  SEN_OR3B_0P5 U483 ( .B1(net59353), .B2(net60540), .A(n818), .X(net59278) );
  SEN_BUF_1 U485 ( .A(net59310), .X(n351) );
  SEN_ND2B_V1_4 U486 ( .A(net59730), .B(n483), .X(net59375) );
  SEN_ND2_8 U487 ( .A1(n361), .A2(n479), .X(n477) );
  SEN_INV_S_6 U488 ( .A(net59688), .X(net59769) );
  SEN_INV_AS_5 U489 ( .A(net59336), .X(net59798) );
  SEN_AOI21B_3 U491 ( .A1(net59654), .A2(n601), .B(n741), .X(n742) );
  SEN_INV_1 U494 ( .A(n809), .X(n815) );
  SEN_ND2_6 U496 ( .A1(n390), .A2(n577), .X(n578) );
  SEN_ND2B_16 U499 ( .A(FirstCyc), .B(CI), .X(n655) );
  SEN_AN2_6 U500 ( .A1(n1055), .A2(n419), .X(net60205) );
  SEN_INV_4 U502 ( .A(net59792), .X(n352) );
  SEN_ND2B_V1_3 U506 ( .A(n420), .B(n515), .X(n518) );
  SEN_INV_5 U508 ( .A(net59777), .X(net59743) );
  SEN_NR2B_12 U509 ( .A(FirstCyc), .B(N72), .X(n658) );
  SEN_AOAI211_4 U511 ( .A1(net59626), .A2(n516), .B(net59353), .C(n517), .X(
        n510) );
  SEN_INV_4 U513 ( .A(n648), .X(n686) );
  SEN_INV_S_3 U515 ( .A(net59309), .X(net59746) );
  SEN_NR2_T_1P5 U517 ( .A1(net59314), .A2(net59731), .X(n704) );
  SEN_ND2_T_6 U518 ( .A1(net60861), .A2(net59342), .X(net59314) );
  SEN_INV_0P8 U519 ( .A(net59333), .X(net59325) );
  SEN_ND2_S_4 U521 ( .A1(net59767), .A2(net59768), .X(net59316) );
  SEN_ND2_S_2 U522 ( .A1(B[4]), .A2(net59990), .X(net59767) );
  SEN_INV_S_3 U525 ( .A(n352), .X(n354) );
  SEN_EN3_3 U528 ( .A1(net59212), .A2(net59513), .A3(net59214), .X(net58915)
         );
  SEN_INV_1P25 U529 ( .A(net59213), .X(net59513) );
  SEN_ND2_T_1 U539 ( .A1(n800), .A2(net58914), .X(n801) );
  SEN_EO2_0P5 U540 ( .A1(net59242), .A2(net59241), .X(n356) );
  SEN_AN2_4 U541 ( .A1(net59462), .A2(net58914), .X(n357) );
  SEN_ND2_2 U542 ( .A1(n737), .A2(n736), .X(n442) );
  SEN_INV_5 U547 ( .A(n1053), .X(n597) );
  SEN_ND2_4 U550 ( .A1(net59310), .A2(net59311), .X(net59750) );
  SEN_INV_1 U553 ( .A(net59335), .X(net59770) );
  SEN_INV_S_0P5 U554 ( .A(n342), .X(n392) );
  SEN_BUF_S_3 U555 ( .A(n555), .X(n362) );
  SEN_ND2_S_4 U556 ( .A1(net59654), .A2(net59677), .X(net59374) );
  SEN_INV_S_0P5 U562 ( .A(n509), .X(n413) );
  SEN_INV_32 U564 ( .A(n364), .X(n363) );
  SEN_ND2B_V1DG_4 U565 ( .A(net60411), .B(net59437), .X(net61810) );
  SEN_ND2_T_8 U566 ( .A1(net60989), .A2(net61305), .X(n515) );
  SEN_INV_3 U574 ( .A(net59411), .X(net59212) );
  SEN_NR2_T_4 U577 ( .A1(net59776), .A2(net59777), .X(net61110) );
  SEN_EN2_DG_8 U579 ( .A1(net58984), .A2(net58985), .X(n364) );
  SEN_ND2_T_4 U580 ( .A1(n482), .A2(n380), .X(net61348) );
  SEN_INV_4 U581 ( .A(n470), .X(n482) );
  SEN_ND2_6 U582 ( .A1(net59651), .A2(net59675), .X(net59624) );
  SEN_INV_S_3 U583 ( .A(n751), .X(n596) );
  SEN_INV_S_6 U584 ( .A(n515), .X(net59353) );
  SEN_ND2_T_4 U586 ( .A1(B[1]), .A2(net59469), .X(n683) );
  SEN_ND2_S_2 U587 ( .A1(n543), .A2(net58945), .X(n542) );
  SEN_EO2_G_2 U588 ( .A1(net59285), .A2(net59286), .X(net58945) );
  SEN_NR2_T_2 U593 ( .A1(n699), .A2(net59739), .X(net60983) );
  SEN_EO2_0P5 U595 ( .A1(A[27]), .A2(net59978), .X(n766) );
  SEN_EO2_DG_2 U596 ( .A1(A[16]), .A2(net59976), .X(net59593) );
  SEN_ND2_T_2 U597 ( .A1(n599), .A2(net59300), .X(n807) );
  SEN_NR3_T_4 U600 ( .A1(n471), .A2(net59624), .A3(net59621), .X(n470) );
  SEN_INV_4 U601 ( .A(net59370), .X(n471) );
  SEN_AOAI211_4 U602 ( .A1(n1050), .A2(net59689), .B(net59769), .C(net59686), 
        .X(net59759) );
  SEN_INV_2P5 U603 ( .A(net59356), .X(n509) );
  SEN_AOAI211_8 U604 ( .A1(net59636), .A2(net61215), .B(net59638), .C(net59639), .X(net59356) );
  SEN_INV_3 U605 ( .A(net59727), .X(net59725) );
  SEN_ND2_T_4 U606 ( .A1(net61348), .A2(n515), .X(n512) );
  SEN_NR3_T_3 U608 ( .A1(net59624), .A2(n1053), .A3(n739), .X(net59638) );
  SEN_ND2_T_3 U609 ( .A1(n352), .A2(n389), .X(net59333) );
  SEN_ND2_T_4 U610 ( .A1(n580), .A2(net59748), .X(n702) );
  SEN_AOI21B_4 U612 ( .A1(net59654), .A2(n601), .B(net59347), .X(net59675) );
  SEN_NR2_8 U614 ( .A1(n687), .A2(n1062), .X(n397) );
  SEN_ND2B_6 U621 ( .A(net61110), .B(n1048), .X(net59311) );
  SEN_ND2_8 U622 ( .A1(n578), .A2(n684), .X(net59799) );
  SEN_ND3_T_1P5 U623 ( .A1(net59341), .A2(net59686), .A3(net59316), .X(n473)
         );
  SEN_INV_8 U626 ( .A(net59291), .X(net59717) );
  SEN_ND2_G_4 U628 ( .A1(n481), .A2(n480), .X(n476) );
  SEN_ND2_T_8 U630 ( .A1(n644), .A2(n643), .X(net59322) );
  SEN_AOAI211_6 U636 ( .A1(net59689), .A2(n1050), .B(n705), .C(n704), .X(n706)
         );
  SEN_BUF_AS_5 U637 ( .A(net59696), .X(net61305) );
  SEN_AOI221_4 U638 ( .A1(n728), .A2(n727), .B1(n726), .B2(n807), .C(n1047), 
        .X(net59696) );
  SEN_ND2_T_6 U639 ( .A1(net59781), .A2(n461), .X(net59777) );
  SEN_ND3_T_4 U641 ( .A1(n596), .A2(n597), .A3(net60873), .X(n598) );
  SEN_INV_S_8 U643 ( .A(net59305), .X(net59677) );
  SEN_ND2_T_4 U644 ( .A1(net59958), .A2(n698), .X(net59305) );
  SEN_INV_S_6 U649 ( .A(net59332), .X(n411) );
  SEN_ND2_T_1P5 U650 ( .A1(n743), .A2(n742), .X(n751) );
  SEN_INV_S_6 U656 ( .A(n665), .X(n833) );
  SEN_NR2_S_5 U659 ( .A1(net60418), .A2(net59385), .X(n495) );
  SEN_AN3B_8 U661 ( .B1(net60861), .B2(net59342), .A(net59335), .X(n479) );
  SEN_OA21_8 U662 ( .A1(net59349), .A2(net59585), .B(n501), .X(n388) );
  SEN_AOAI211_8 U663 ( .A1(n499), .A2(net59258), .B(n500), .C(n485), .X(n498)
         );
  SEN_NR2_G_2 U664 ( .A1(n520), .A2(net61338), .X(net60418) );
  SEN_OAI21_S_4 U667 ( .A1(net59372), .A2(net59374), .B(n719), .X(n729) );
  SEN_ND2_4 U669 ( .A1(n800), .A2(n357), .X(n791) );
  SEN_OAI21_T_6 U673 ( .A1(n558), .A2(n559), .B(n560), .X(n528) );
  SEN_ND3_3 U675 ( .A1(n472), .A2(n444), .A3(n473), .X(n483) );
  SEN_AOI21_T_2 U679 ( .A1(net59461), .A2(net59462), .B(net59463), .X(n573) );
  SEN_NR2_T_2 U681 ( .A1(n564), .A2(n446), .X(net59494) );
  SEN_AOAI211_8 U683 ( .A1(n509), .A2(n508), .B(n510), .C(n511), .X(net59583)
         );
  SEN_OAI211_4 U684 ( .A1(n1044), .A2(net59305), .B1(net59729), .B2(net59372), 
        .X(net59679) );
  SEN_ND2B_V1DG_2 U685 ( .A(n430), .B(net59456), .X(n776) );
  SEN_ND2B_1 U688 ( .A(net59238), .B(net59239), .X(net59500) );
  SEN_AN2_2 U689 ( .A1(net59498), .A2(net59500), .X(net59497) );
  SEN_INV_2 U690 ( .A(net59239), .X(net59503) );
  SEN_INV_S_3 U691 ( .A(net59258), .X(net59382) );
  SEN_INV_1 U693 ( .A(net59561), .X(n487) );
  SEN_ND2B_2 U694 ( .A(net59400), .B(net59409), .X(net59562) );
  SEN_ND2B_6 U695 ( .A(N72), .B(INST[2]), .X(n836) );
  SEN_OR2_1 U696 ( .A1(net60372), .A2(net60373), .X(net59584) );
  SEN_NR3_T_2 U697 ( .A1(n502), .A2(net59382), .A3(n503), .X(n500) );
  SEN_INV_S_0P5 U698 ( .A(net59392), .X(net59406) );
  SEN_ND2_G_1 U700 ( .A1(n722), .A2(n721), .X(net59300) );
  SEN_ND2_T_1P5 U701 ( .A1(net59277), .A2(net59617), .X(net59276) );
  SEN_OR2_1 U702 ( .A1(net60377), .A2(net60378), .X(net59393) );
  SEN_INV_2 U703 ( .A(net59398), .X(net59240) );
  SEN_INV_3 U704 ( .A(n590), .X(net59958) );
  SEN_INV_S_2 U705 ( .A(n787), .X(n830) );
  SEN_INV_24 U706 ( .A(INST[1]), .X(n425) );
  SEN_NR2_T_2 U707 ( .A1(net59746), .A2(net59306), .X(n701) );
  SEN_INV_S_12 U708 ( .A(INST[3]), .X(n415) );
  SEN_INV_1 U709 ( .A(n610), .X(n611) );
  SEN_INV_S_2 U710 ( .A(net59409), .X(n491) );
  SEN_NR2_T_5 U712 ( .A1(INST[2]), .A2(INST[1]), .X(n657) );
  SEN_NR2_G_8 U713 ( .A1(INST[1]), .A2(A[31]), .X(n653) );
  SEN_INV_S_0P5 U714 ( .A(net59257), .X(net59386) );
  SEN_OR2_3 U715 ( .A1(net60375), .A2(net60376), .X(net59549) );
  SEN_INV_S_2 U716 ( .A(net59418), .X(net59455) );
  SEN_ND2_S_0P5 U717 ( .A1(net59422), .A2(net59455), .X(net59438) );
  SEN_INV_24 U719 ( .A(B[2]), .X(n455) );
  SEN_ND2_T_6 U720 ( .A1(n395), .A2(n646), .X(net59321) );
  SEN_EO2_1 U721 ( .A1(A[5]), .A2(net59976), .X(net59760) );
  SEN_ND2_2 U723 ( .A1(n584), .A2(n585), .X(n715) );
  SEN_ND2_2 U724 ( .A1(A[11]), .A2(net59980), .X(n584) );
  SEN_ND2_T_1 U725 ( .A1(n583), .A2(net59444), .X(n585) );
  SEN_ND2_S_1 U726 ( .A1(net59630), .A2(net59631), .X(net59280) );
  SEN_ND2_T_1 U727 ( .A1(n395), .A2(net59691), .X(net59274) );
  SEN_OR2_1 U728 ( .A1(net60380), .A2(net60381), .X(net59277) );
  SEN_INV_2 U729 ( .A(net59584), .X(net59351) );
  SEN_ND2_2 U730 ( .A1(net59605), .A2(net59606), .X(net59258) );
  SEN_ND2_G_1 U731 ( .A1(net59584), .A2(net59350), .X(n501) );
  SEN_ND2_S_1 U732 ( .A1(n754), .A2(n753), .X(net59252) );
  SEN_ND2_S_0P5 U733 ( .A1(B[16]), .A2(net59990), .X(n754) );
  SEN_MUXI2_S_0P5 U734 ( .D0(n575), .D1(n794), .S(B[17]), .X(n753) );
  SEN_ND2_T_1 U735 ( .A1(net59600), .A2(net59601), .X(net59389) );
  SEN_OR2_1 U736 ( .A1(n603), .A2(n604), .X(net59242) );
  SEN_ND2_2 U737 ( .A1(net59564), .A2(net59242), .X(net59400) );
  SEN_ND2_T_1 U739 ( .A1(n762), .A2(n761), .X(net59239) );
  SEN_ND2_2 U740 ( .A1(n395), .A2(net59538), .X(net59238) );
  SEN_ND2_G_1 U741 ( .A1(net59536), .A2(net59537), .X(net59233) );
  SEN_ND2_2 U742 ( .A1(net59530), .A2(net59531), .X(net59410) );
  SEN_EN3_1 U743 ( .A1(net59290), .A2(net59291), .A3(net59287), .X(net58947)
         );
  SEN_EN3_0P5 U744 ( .A1(net59237), .A2(net59238), .A3(net59239), .X(net58919)
         );
  SEN_EO2_S_0P5 U745 ( .A1(n832), .A2(net59221), .X(net59412) );
  SEN_EO2_S_0P5 U746 ( .A1(n830), .A2(net60361), .X(n453) );
  SEN_EN2_0P5 U747 ( .A1(n557), .A2(net59429), .X(net60464) );
  SEN_MUXI2_S_1 U748 ( .D0(n625), .D1(n961), .S(B[31]), .X(n965) );
  SEN_AN2_1 U749 ( .A1(n994), .A2(n993), .X(n365) );
  SEN_AN2_1 U750 ( .A1(n888), .A2(n887), .X(n366) );
  SEN_AN2_1 U751 ( .A1(n984), .A2(n983), .X(n367) );
  SEN_AN2_1 U752 ( .A1(n925), .A2(n924), .X(n368) );
  SEN_AN2_1 U753 ( .A1(n898), .A2(n897), .X(n369) );
  SEN_AN2_1 U754 ( .A1(n944), .A2(n943), .X(n370) );
  SEN_AN2_1 U755 ( .A1(n955), .A2(n954), .X(n371) );
  SEN_AN2_1 U756 ( .A1(n989), .A2(n988), .X(n372) );
  SEN_OR2_DG_1 U757 ( .A1(n562), .A2(net59213), .X(n373) );
  SEN_ND2_S_3 U759 ( .A1(net59754), .A2(net59755), .X(net59306) );
  SEN_INV_1P5 U760 ( .A(net59306), .X(net59730) );
  SEN_INV_2 U761 ( .A(n792), .X(n794) );
  SEN_ND3B_1 U762 ( .A(INST[2]), .B1(N72), .B2(INST[1]), .X(n850) );
  SEN_AN2_S_0P5 U763 ( .A1(net59680), .A2(net59306), .X(n375) );
  SEN_AOAI211_G_1 U765 ( .A1(net59400), .A2(n491), .B(net59561), .C(net59562), 
        .X(net59559) );
  SEN_INV_S_1 U766 ( .A(net59559), .X(net59542) );
  SEN_AN2_1 U767 ( .A1(n920), .A2(n919), .X(n376) );
  SEN_AN2_1 U768 ( .A1(n909), .A2(n908), .X(n377) );
  SEN_AN2_1 U770 ( .A1(n1017), .A2(n1016), .X(n378) );
  SEN_AN2_1 U771 ( .A1(n847), .A2(n846), .X(n379) );
  SEN_OR2_1 U772 ( .A1(net59621), .A2(net59622), .X(n380) );
  SEN_AN2_1 U773 ( .A1(n893), .A2(n892), .X(n381) );
  SEN_AN2_1 U774 ( .A1(n999), .A2(n998), .X(n382) );
  SEN_AN2_1 U775 ( .A1(n979), .A2(n978), .X(n383) );
  SEN_AN2_1 U776 ( .A1(n933), .A2(n932), .X(n384) );
  SEN_ND3_1 U777 ( .A1(n779), .A2(n778), .A3(net59457), .X(net59488) );
  SEN_INV_S_1 U778 ( .A(net59488), .X(n439) );
  SEN_AN2_1 U779 ( .A1(n960), .A2(n959), .X(n385) );
  SEN_AN2_1 U780 ( .A1(n965), .A2(n964), .X(n386) );
  SEN_ND2_0P5 U781 ( .A1(net59888), .A2(net59200), .X(n837) );
  SEN_OAI21_S_1 U782 ( .A1(net59505), .A2(net59482), .B(net60361), .X(net59473) );
  SEN_INV_2 U783 ( .A(net59473), .X(net59462) );
  SEN_OAI21_G_1 U784 ( .A1(n836), .A2(INST[1]), .B(n614), .X(n387) );
  SEN_ND3_T_16 U785 ( .A1(INST[1]), .A2(INST[2]), .A3(N72), .X(n389) );
  SEN_INV_4 U790 ( .A(net59651), .X(net59642) );
  SEN_OAI21_S_8 U791 ( .A1(n345), .A2(net59750), .B(n475), .X(n474) );
  SEN_INV_S_0P5 U792 ( .A(n471), .X(n393) );
  SEN_INV_4 U793 ( .A(net59966), .X(n394) );
  SEN_INV_4 U794 ( .A(net59966), .X(n395) );
  SEN_INV_S_4 U796 ( .A(n389), .X(net59966) );
  SEN_INV_3 U797 ( .A(n793), .X(n396) );
  SEN_INV_S_12 U799 ( .A(net59870), .X(net59469) );
  SEN_INV_2 U800 ( .A(n720), .X(n728) );
  SEN_ND3_T_2 U801 ( .A1(net59635), .A2(n828), .A3(n809), .X(n720) );
  SEN_INV_1P25 U804 ( .A(n691), .X(n582) );
  SEN_INV_1P5 U805 ( .A(n734), .X(n726) );
  SEN_OR2_5 U806 ( .A1(n677), .A2(n676), .X(n399) );
  SEN_OR2_2 U807 ( .A1(n678), .A2(n405), .X(n400) );
  SEN_OAI21_G_1 U811 ( .A1(n656), .A2(n408), .B(n608), .X(n405) );
  SEN_ND2_G_4 U814 ( .A1(n394), .A2(n752), .X(net59251) );
  SEN_OAI31_2 U815 ( .A1(net59252), .A2(net59389), .A3(net59597), .B(net59598), 
        .X(n505) );
  SEN_EO2_0P5 U817 ( .A1(A[30]), .A2(net59444), .X(n798) );
  SEN_EO2_S_1 U818 ( .A1(n401), .A2(n410), .X(net59329) );
  SEN_ND2_3 U822 ( .A1(net59635), .A2(n828), .X(n723) );
  SEN_ND2_8 U824 ( .A1(net59958), .A2(n712), .X(net59291) );
  SEN_OA31_8 U825 ( .A1(net59287), .A2(net59717), .A3(n822), .B(n714), .X(n599) );
  SEN_ND2_S_3 U827 ( .A1(n394), .A2(net59575), .X(net59550) );
  SEN_ND2_S_0P5 U828 ( .A1(net59549), .A2(net59248), .X(n489) );
  SEN_NR3_T_3 U830 ( .A1(n541), .A2(net59282), .A3(n542), .X(n539) );
  SEN_ND2B_6 U831 ( .A(FirstCyc), .B(CI), .X(n608) );
  SEN_INV_4 U832 ( .A(n689), .X(n677) );
  SEN_ND2_6 U834 ( .A1(n587), .A2(n588), .X(n712) );
  SEN_ND2_3 U835 ( .A1(n586), .A2(net59978), .X(n588) );
  SEN_ND2_S_4 U836 ( .A1(net59287), .A2(net59717), .X(n824) );
  SEN_ND2_G_4 U837 ( .A1(n574), .A2(n642), .X(n792) );
  SEN_INV_3 U838 ( .A(n651), .X(n660) );
  SEN_AN2_DG_1 U839 ( .A1(net59635), .A2(net59276), .X(net60495) );
  SEN_ND2_S_16 U841 ( .A1(FirstCyc), .A2(N72), .X(n408) );
  SEN_NR2_S_5 U842 ( .A1(n667), .A2(n666), .X(n651) );
  SEN_ND2_T_4 U844 ( .A1(net59304), .A2(n374), .X(net59651) );
  SEN_OA21_8 U845 ( .A1(n693), .A2(n692), .B(n691), .X(n456) );
  SEN_AO21B_8 U846 ( .A1(n737), .A2(n824), .B(n599), .X(n809) );
  SEN_ND2_2 U849 ( .A1(n711), .A2(n710), .X(net59287) );
  SEN_ND2_T_2 U850 ( .A1(net59300), .A2(n732), .X(n810) );
  SEN_MUXI2_S_2 U851 ( .D0(n575), .D1(n716), .S(B[9]), .X(n710) );
  SEN_INV_S_0P5 U852 ( .A(n471), .X(n445) );
  SEN_ND2B_6 U856 ( .A(N72), .B(INST[1]), .X(n665) );
  SEN_ND2_S_4 U857 ( .A1(net59666), .A2(net59667), .X(net59622) );
  SEN_ND3_2 U858 ( .A1(n734), .A2(n733), .A3(n738), .X(net59667) );
  SEN_INV_2 U859 ( .A(n811), .X(n738) );
  SEN_ND2_G_1 U861 ( .A1(n732), .A2(net59671), .X(n811) );
  SEN_ND2_T_4 U862 ( .A1(n579), .A2(n417), .X(n580) );
  SEN_INV_2 U863 ( .A(INST[2]), .X(net59849) );
  SEN_ND3_T_4 U864 ( .A1(n416), .A2(INST[2]), .A3(B[1]), .X(n664) );
  SEN_INV_32 U865 ( .A(INST[3]), .X(n416) );
  SEN_INV_S_2 U866 ( .A(net60235), .X(net59401) );
  SEN_INV_4 U868 ( .A(n685), .X(n577) );
  SEN_EN3_0P5 U869 ( .A1(n353), .A2(net59350), .A3(net59351), .X(net58935) );
  SEN_ND2_S_0P5 U871 ( .A1(n413), .A2(net59270), .X(n818) );
  SEN_ND2_G_1 U873 ( .A1(net60495), .A2(net59633), .X(n516) );
  SEN_INV_3 U875 ( .A(n743), .X(n739) );
  SEN_INV_10 U876 ( .A(net59321), .X(net59342) );
  SEN_NR2_S_2 U877 ( .A1(n720), .A2(n740), .X(n719) );
  SEN_INV_6 U880 ( .A(n589), .X(net59962) );
  SEN_ND2B_V1_8 U881 ( .A(net59205), .B(n464), .X(net59873) );
  SEN_INV_S_0P5 U882 ( .A(net59276), .X(n420) );
  SEN_AO21B_2 U883 ( .A1(n421), .A2(n422), .B(net59583), .X(n484) );
  SEN_INV_S_0P5 U884 ( .A(net60372), .X(n421) );
  SEN_INV_S_0P5 U885 ( .A(net60373), .X(n422) );
  SEN_NR2B_V1_8 U887 ( .A(net59455), .B(net59474), .X(n424) );
  SEN_ND2_T_16 U889 ( .A1(n425), .A2(A[31]), .X(n466) );
  SEN_OAI211_8 U890 ( .A1(n426), .A2(A[31]), .B1(FirstCyc), .B2(INST[2]), .X(
        n692) );
  SEN_INV_S_32 U891 ( .A(B[31]), .X(n426) );
  SEN_AO22_8 U892 ( .A1(n343), .A2(n679), .B1(n427), .B2(n428), .X(n681) );
  SEN_INV_1 U893 ( .A(INST[1]), .X(n428) );
  SEN_AOI21_T_12 U896 ( .A1(A[31]), .A2(B[31]), .B(N72), .X(n467) );
  SEN_INV_S_3 U897 ( .A(net59346), .X(net59372) );
  SEN_INV_S_1 U898 ( .A(n772), .X(n430) );
  SEN_INV_S_1 U899 ( .A(net60411), .X(n431) );
  SEN_INV_S_0P5 U900 ( .A(n746), .X(n747) );
  SEN_INV_S_2 U902 ( .A(net59270), .X(net59635) );
  SEN_INV_2 U904 ( .A(net59550), .X(net59248) );
  SEN_INV_S_1 U906 ( .A(net59438), .X(n432) );
  SEN_INV_S_1 U907 ( .A(n557), .X(n434) );
  SEN_OR4_4 U911 ( .A1(n1053), .A2(n739), .A3(n729), .A4(net59642), .X(
        net60989) );
  SEN_INV_4 U912 ( .A(net59316), .X(net59731) );
  SEN_EO2_S_1 U913 ( .A1(net59390), .A2(net59391), .X(net58925) );
  SEN_INV_S_0P5 U915 ( .A(net59215), .X(n438) );
  SEN_BUF_1 U918 ( .A(net59304), .X(n441) );
  SEN_INV_0P8 U919 ( .A(n822), .X(n737) );
  SEN_ND2_S_8 U920 ( .A1(net59700), .A2(net59267), .X(n828) );
  SEN_ND2_S_3 U921 ( .A1(n718), .A2(n717), .X(net59267) );
  SEN_INV_S_6 U922 ( .A(net59264), .X(net59700) );
  SEN_OAI221_2 U923 ( .A1(net59212), .A2(net59213), .B1(net59212), .B2(
        net59214), .C(net59215), .X(net59211) );
  SEN_BUF_1 U924 ( .A(n1057), .X(n448) );
  SEN_INV_S_0P5 U926 ( .A(n448), .X(n454) );
  SEN_ND3_T_4 U927 ( .A1(net59461), .A2(net59455), .A3(net59462), .X(n797) );
  SEN_EO3_1 U928 ( .A1(n454), .A2(net59248), .A3(net59249), .X(net58927) );
  SEN_MUXI2_S_1 U929 ( .D0(net58935), .D1(n376), .S(INST[3]), .X(Z[15]) );
  SEN_INV_0P8 U930 ( .A(net58935), .X(net59282) );
  SEN_MUXI2_S_8 U931 ( .D0(n681), .D1(n575), .S(n455), .X(n682) );
  SEN_INV_16 U932 ( .A(INST[1]), .X(net59888) );
  SEN_ND2_T_16 U933 ( .A1(FirstCyc), .A2(N72), .X(n607) );
  SEN_OAI21_3 U934 ( .A1(n656), .A2(n408), .B(n608), .X(n610) );
  SEN_OR3B_12 U935 ( .B1(INST[3]), .B2(n836), .A(INST[1]), .X(net59870) );
  SEN_INV_S_6 U936 ( .A(net59992), .X(net59990) );
  SEN_MUXI2_DG_2 U937 ( .D0(n575), .D1(n716), .S(B[5]), .X(net59768) );
  SEN_ND2_S_4 U938 ( .A1(n459), .A2(net60751), .X(net59411) );
  SEN_ND2_2 U940 ( .A1(net59714), .A2(net59715), .X(net59270) );
  SEN_MUXI2_DG_1 U943 ( .D0(n1040), .D1(n1039), .S(INST[3]), .X(Z[26]) );
  SEN_MUXI2_S_1 U944 ( .D0(n623), .D1(n628), .S(B[31]), .X(n962) );
  SEN_AN4B_0P5 U946 ( .B1(net59311), .B2(n351), .B3(net59309), .A(net59312), 
        .X(net59308) );
  SEN_INV_2 U947 ( .A(n824), .X(n740) );
  SEN_ND3_T_4 U948 ( .A1(net59744), .A2(net59743), .A3(net59343), .X(n481) );
  SEN_OAI2111_4 U951 ( .A1(net59343), .A2(net59314), .B1(net59310), .B2(
        net59311), .B3(net59309), .X(net59690) );
  SEN_ND2B_V1_1 U953 ( .A(net59280), .B(net59276), .X(net59621) );
  SEN_OA21_2 U954 ( .A1(net59624), .A2(n471), .B(net59622), .X(net60540) );
  SEN_OAI21_S_1P5 U955 ( .A1(net60532), .A2(net59372), .B(n445), .X(net59362)
         );
  SEN_AN2_S_0P5 U956 ( .A1(n393), .A2(n1076), .X(net60557) );
  SEN_INV_S_1 U957 ( .A(net59314), .X(net59686) );
  SEN_ND2_T_8 U959 ( .A1(net59794), .A2(net59962), .X(net59335) );
  SEN_ND2_T_1 U960 ( .A1(net59958), .A2(net59760), .X(net59315) );
  SEN_AN3B_4 U961 ( .B1(n493), .B2(net59542), .A(n494), .X(net59543) );
  SEN_ND2_2 U962 ( .A1(n487), .A2(net59406), .X(n493) );
  SEN_NR3B_1 U963 ( .A(n492), .B1(n491), .B2(net59392), .X(n494) );
  SEN_ND2_S_3 U964 ( .A1(net59241), .A2(net59558), .X(n492) );
  SEN_ND2_S_0P5 U965 ( .A1(n395), .A2(net59560), .X(net59392) );
  SEN_NR3_T_2 U966 ( .A1(n490), .A2(net59402), .A3(n491), .X(n488) );
  SEN_INV_2 U967 ( .A(n492), .X(n490) );
  SEN_INV_S_3 U968 ( .A(net59393), .X(net59402) );
  SEN_BUF_1 U970 ( .A(n486), .X(net60235) );
  SEN_AOAI211_G_1 U971 ( .A1(net59380), .A2(n503), .B(n505), .C(net59595), .X(
        n507) );
  SEN_AOI311_2 U972 ( .A1(n504), .A2(net59386), .A3(net59389), .B1(n506), .B2(
        n507), .X(n497) );
  SEN_ND2_S_0P5 U973 ( .A1(net59251), .A2(net59594), .X(n504) );
  SEN_NR2_S_0P5 U974 ( .A1(net59257), .A2(n505), .X(n506) );
  SEN_ND2_S_0P5 U975 ( .A1(n394), .A2(net59593), .X(net59257) );
  SEN_INV_S_0P5 U976 ( .A(n505), .X(n499) );
  SEN_INV_1 U977 ( .A(n504), .X(n502) );
  SEN_INV_S_0P5 U978 ( .A(net59389), .X(n503) );
  SEN_INV_S_0P5 U979 ( .A(n485), .X(net59381) );
  SEN_ND2_S_0P5 U980 ( .A1(net59958), .A2(net59608), .X(net59585) );
  SEN_INV_S_6 U981 ( .A(net59583), .X(net59349) );
  SEN_INV_2 U982 ( .A(net59585), .X(net59350) );
  SEN_ND2B_S_0P5 U983 ( .A(n392), .B(n519), .X(net59255) );
  SEN_INV_0P65 U984 ( .A(net59622), .X(net59633) );
  SEN_AOI21B_1 U985 ( .A1(net59629), .A2(net59274), .B(net59280), .X(n517) );
  SEN_INV_S_0P5 U986 ( .A(net59277), .X(net59629) );
  SEN_AOAI211_6 U987 ( .A1(net59356), .A2(net59270), .B(n512), .C(n513), .X(
        n511) );
  SEN_NR2_G_1 U988 ( .A1(n514), .A2(net59279), .X(n513) );
  SEN_NR3_0P5 U989 ( .A1(net59280), .A2(net59277), .A3(net59617), .X(n514) );
  SEN_INV_S_3 U990 ( .A(net59274), .X(net59617) );
  SEN_ND2_S_0P5 U991 ( .A1(n394), .A2(net59616), .X(net59279) );
  SEN_NR2_T_1 U992 ( .A1(net59583), .A2(net59584), .X(n520) );
  SEN_EO2_2 U997 ( .A1(net59396), .A2(net59397), .X(net58921) );
  SEN_NR3_T_2 U998 ( .A1(n537), .A2(n536), .A3(n535), .X(n534) );
  SEN_INV_1 U999 ( .A(net58925), .X(n535) );
  SEN_AN4B_2 U1002 ( .B1(n539), .B2(net58937), .B3(net58941), .A(n540), .X(
        n538) );
  SEN_ND2_S_1 U1003 ( .A1(net58943), .A2(net58939), .X(n541) );
  SEN_EN3_1 U1004 ( .A1(net59263), .A2(net59264), .A3(net59267), .X(net58943)
         );
  SEN_EN3_1 U1005 ( .A1(net59273), .A2(net59274), .A3(net59277), .X(net58939)
         );
  SEN_NR2_S_1 U1006 ( .A1(n544), .A2(n545), .X(n543) );
  SEN_INV_1 U1007 ( .A(net58947), .X(n544) );
  SEN_ND2_S_1 U1008 ( .A1(n546), .A2(net58949), .X(n545) );
  SEN_NR2_S_1 U1009 ( .A1(n547), .A2(n548), .X(n546) );
  SEN_INV_1 U1010 ( .A(net58951), .X(n547) );
  SEN_EN3_0P5 U1011 ( .A1(net60532), .A2(net59345), .A3(net59346), .X(net58951) );
  SEN_ND3_S_1 U1012 ( .A1(n549), .A2(net58957), .A3(net58954), .X(n548) );
  SEN_NR2_S_1 U1013 ( .A1(n550), .A2(n551), .X(n549) );
  SEN_INV_1 U1014 ( .A(net58960), .X(n550) );
  SEN_EN2_1 U1015 ( .A1(net59337), .A2(net59338), .X(net58960) );
  SEN_ND2_S_1 U1016 ( .A1(n552), .A2(net58963), .X(n551) );
  SEN_NR2_S_1 U1017 ( .A1(n553), .A2(n554), .X(n552) );
  SEN_INV_1 U1018 ( .A(net58965), .X(n553) );
  SEN_EN3_0P5 U1019 ( .A1(net61773), .A2(net59335), .A3(n1050), .X(net58965)
         );
  SEN_ND2_S_1 U1020 ( .A1(net58967), .A2(net58970), .X(n554) );
  SEN_EN2_1 U1021 ( .A1(net59328), .A2(net59329), .X(net58967) );
  SEN_EN3_0P5 U1023 ( .A1(net59320), .A2(net59321), .A3(n1061), .X(net58963)
         );
  SEN_EO2_1 U1024 ( .A1(net59307), .A2(net59308), .X(net58957) );
  SEN_EN3_0P5 U1025 ( .A1(net59298), .A2(net59299), .A3(net59300), .X(net58949) );
  SEN_EN2_1 U1026 ( .A1(net59271), .A2(net59272), .X(net58937) );
  SEN_EN2_1 U1027 ( .A1(net59261), .A2(net59262), .X(net58941) );
  SEN_INV_1 U1028 ( .A(net58933), .X(n540) );
  SEN_EO2_1 U1029 ( .A1(net59255), .A2(net59256), .X(net58933) );
  SEN_EN3_0P5 U1030 ( .A1(net59250), .A2(net59251), .A3(net59252), .X(net58931) );
  SEN_EN2_1 U1031 ( .A1(net59240), .A2(n356), .X(net58923) );
  SEN_EN2_0P5 U1033 ( .A1(net59216), .A2(net59217), .X(n530) );
  SEN_INV_S_1 U1034 ( .A(net58913), .X(net59217) );
  SEN_ND4B_1 U1035 ( .A(net58986), .B1(net58987), .B2(net58988), .B3(net58989), 
        .X(n523) );
  SEN_INV_S_0P5 U1036 ( .A(n523), .X(n525) );
  SEN_ND2_G_1 U1037 ( .A1(INST[3]), .A2(n523), .X(n526) );
  SEN_INV_S_1 U1038 ( .A(net59433), .X(net58984) );
  SEN_INV_S_1 U1039 ( .A(net59431), .X(net58985) );
  SEN_AO31_0P5 U1040 ( .A1(net59418), .A2(net59419), .A3(n557), .B(net59429), 
        .X(net60411) );
  SEN_MUXI2_S_0P5 U1041 ( .D0(n521), .D1(n386), .S(INST[3]), .X(Z[31]) );
  SEN_AN3B_4 U1042 ( .B1(net59440), .B2(net59425), .A(n568), .X(n558) );
  SEN_AO31_2 U1043 ( .A1(net60751), .A2(n459), .A3(net59214), .B(net60246), 
        .X(net59440) );
  SEN_ND2B_1 U1044 ( .A(n557), .B(net59422), .X(n559) );
  SEN_AOI21_G_0P75 U1045 ( .A1(B[29]), .A2(net59990), .B(net59470), .X(n557)
         );
  SEN_ND2_G_1 U1046 ( .A1(net59465), .A2(net59466), .X(net59422) );
  SEN_AOI32_2 U1048 ( .A1(net59456), .A2(net59457), .A3(net59410), .B1(n449), 
        .B2(net59410), .X(n561) );
  SEN_INV_S_1 U1049 ( .A(net59232), .X(net59457) );
  SEN_ND2B_S_2 U1050 ( .A(net59454), .B(net59455), .X(n562) );
  SEN_ND2_S_0P5 U1051 ( .A1(n395), .A2(net59523), .X(net59213) );
  SEN_ND3B_V1DG_2 U1052 ( .A(net58914), .B1(net60751), .B2(n459), .X(n566) );
  SEN_ND2B_V1_4 U1056 ( .A(n666), .B(n668), .X(n689) );
  SEN_ND2_G_0P65 U1057 ( .A1(n733), .A2(n735), .X(net59666) );
  SEN_NR2_T_16 U1058 ( .A1(INST[2]), .A2(INST[1]), .X(n656) );
  SEN_INV_2 U1059 ( .A(net59362), .X(net59298) );
  SEN_MUXI2_DG_1 U1061 ( .D0(n1042), .D1(n1041), .S(INST[3]), .X(Z[30]) );
  SEN_OR4B_1 U1062 ( .B1(n817), .B2(n816), .B3(n815), .A(n814), .X(net59268)
         );
  SEN_AOI21_G_0P75 U1063 ( .A1(net59252), .A2(net59378), .B(n806), .X(net59377) );
  SEN_INV_0P8 U1064 ( .A(net59378), .X(net59250) );
  SEN_OR3B_4 U1065 ( .B1(INST[1]), .B2(INST[2]), .A(N72), .X(n1012) );
  SEN_AN3_16 U1066 ( .A1(INST[1]), .A2(INST[2]), .A3(N72), .X(n589) );
  SEN_ND3_8 U1067 ( .A1(N72), .A2(B[0]), .A3(INST[1]), .X(n650) );
  SEN_INV_32 U1070 ( .A(N72), .X(net59200) );
  SEN_OAI21_2 U1071 ( .A1(net59240), .A2(net59241), .B(net59400), .X(n804) );
  SEN_ND2B_16 U1072 ( .A(INST[3]), .B(INST[2]), .X(n574) );
  SEN_ND2B_6 U1073 ( .A(INST[3]), .B(INST[2]), .X(n679) );
  SEN_INV_S_1 U1074 ( .A(n795), .X(n576) );
  SEN_INV_S_0P5 U1075 ( .A(net59341), .X(net59320) );
  SEN_INV_S_0P5 U1076 ( .A(net59689), .X(net61773) );
  SEN_OR2_16 U1077 ( .A1(n595), .A2(n343), .X(n642) );
  SEN_ND2_3 U1078 ( .A1(n709), .A2(n708), .X(n822) );
  SEN_ND2_S_1 U1079 ( .A1(B[9]), .A2(net59988), .X(n709) );
  SEN_AOAI211_6 U1080 ( .A1(net59730), .A2(net59731), .B(n707), .C(n706), .X(
        net59727) );
  SEN_ND3B_V1DG_4 U1081 ( .A(n677), .B1(n690), .B2(net59819), .X(n694) );
  SEN_ND2_G_24 U1082 ( .A1(B[1]), .A2(INST[1]), .X(n662) );
  SEN_NR3_T_12 U1083 ( .A1(INST[1]), .A2(INST[2]), .A3(net59200), .X(n595) );
  SEN_MUXI2_DG_5 U1084 ( .D0(n576), .D1(n792), .S(B[4]), .X(n648) );
  SEN_OR3B_2 U1085 ( .B1(n822), .B2(n723), .A(n809), .X(n734) );
  SEN_BUF_S_3 U1086 ( .A(net59637), .X(net61215) );
  SEN_ND3_1 U1087 ( .A1(n442), .A2(n746), .A3(n738), .X(net59637) );
  SEN_ND2_2 U1088 ( .A1(net59958), .A2(n713), .X(n823) );
  SEN_INV_1P5 U1090 ( .A(n808), .X(n735) );
  SEN_AN3B_4 U1091 ( .B1(n702), .B2(n701), .A(n700), .X(n707) );
  SEN_ND2_2 U1092 ( .A1(n824), .A2(n810), .X(n744) );
  SEN_ND3_T_4 U1093 ( .A1(n791), .A2(n790), .A3(n789), .X(net59463) );
  SEN_OAI211_1 U1094 ( .A1(net59263), .A2(net59264), .B1(n829), .B2(n828), .X(
        net59262) );
  SEN_ND2_G_4 U1096 ( .A1(net59958), .A2(n715), .X(net59264) );
  SEN_INV_2 U1097 ( .A(n667), .X(n668) );
  SEN_ND2B_6 U1098 ( .A(INST[3]), .B(DI[31]), .X(n666) );
  SEN_ND4B_8 U1099 ( .A(INST[3]), .B1(n833), .B2(B[0]), .B3(INST[2]), .X(n684)
         );
  SEN_EO2_S_1 U1100 ( .A1(A[7]), .A2(net61246), .X(n697) );
  SEN_ND2_T_2 U1101 ( .A1(net59958), .A2(n697), .X(net59345) );
  SEN_ND2_S_0P8 U1103 ( .A1(n735), .A2(n746), .X(net59636) );
  SEN_EO2_4 U1107 ( .A1(A[12]), .A2(net61246), .X(n724) );
  SEN_EO2_3 U1108 ( .A1(A[6]), .A2(net61246), .X(n698) );
  SEN_ND2_T_2 U1109 ( .A1(net59958), .A2(n724), .X(n827) );
  SEN_EO2_2 U1110 ( .A1(A[15]), .A2(net61246), .X(net59608) );
  SEN_ND2_2 U1111 ( .A1(net59958), .A2(n731), .X(net59299) );
  SEN_EO2_1 U1112 ( .A1(A[8]), .A2(net61241), .X(n731) );
  SEN_INV_S_1 U1113 ( .A(A[11]), .X(n583) );
  SEN_INV_S_1 U1114 ( .A(A[9]), .X(n586) );
  SEN_INV_S_0P5 U1115 ( .A(net59350), .X(net61338) );
  SEN_ND2_S_3 U1116 ( .A1(n770), .A2(n769), .X(net58914) );
  SEN_INV_S_1 U1117 ( .A(net59268), .X(net59263) );
  SEN_ND2_0P5 U1118 ( .A1(net59267), .A2(net59268), .X(n829) );
  SEN_AOI21_G_0P75 U1119 ( .A1(net59287), .A2(net59288), .B(n825), .X(net59286) );
  SEN_INV_2 U1120 ( .A(net59288), .X(net59290) );
  SEN_INV_S_0P5 U1121 ( .A(n827), .X(n725) );
  SEN_MUXI2_S_1 U1122 ( .D0(net58947), .D1(n369), .S(INST[3]), .X(Z[9]) );
  SEN_MUXI2_S_0P5 U1125 ( .D0(net58945), .D1(n381), .S(INST[3]), .X(Z[10]) );
  SEN_MUXI2_S_1 U1126 ( .D0(net58917), .D1(n1038), .S(INST[3]), .X(Z[24]) );
  SEN_ND2_2 U1128 ( .A1(net59264), .A2(net59663), .X(n746) );
  SEN_ND2B_6 U1129 ( .A(B[0]), .B(net59200), .X(n669) );
  SEN_AN3_1 U1130 ( .A1(INST[1]), .A2(INST[2]), .A3(N72), .X(n590) );
  SEN_INV_1 U1131 ( .A(n792), .X(n591) );
  SEN_MUX2_S_0P5 U1132 ( .D0(n575), .D1(n794), .S(B[13]), .X(net60381) );
  SEN_MUXI2_S_1 U1133 ( .D0(n575), .D1(n794), .S(B[18]), .X(net59601) );
  SEN_INV_2 U1135 ( .A(n837), .X(n628) );
  SEN_AOI21_G_1 U1136 ( .A1(n831), .A2(n830), .B(net59473), .X(n786) );
  SEN_INV_S_0P5 U1137 ( .A(n837), .X(n627) );
  SEN_BUF_1 U1138 ( .A(n602), .X(n623) );
  SEN_NR2B_V1_1 U1139 ( .A(n821), .B(net59314), .X(net59312) );
  SEN_AN2_3 U1140 ( .A1(net59346), .A2(net59677), .X(n601) );
  SEN_ND2_0P5 U1141 ( .A1(net59513), .A2(net59410), .X(net59215) );
  SEN_OAI31_0P75 U1142 ( .A1(net59242), .A2(net59409), .A3(net59564), .B(n760), 
        .X(net59561) );
  SEN_INV_0P8 U1143 ( .A(n387), .X(n630) );
  SEN_ND2_S_0P5 U1144 ( .A1(net59213), .A2(net59214), .X(n779) );
  SEN_INV_1 U1145 ( .A(net59380), .X(net59596) );
  SEN_ND2_S_0P8 U1146 ( .A1(n832), .A2(n830), .X(net59505) );
  SEN_ND2_S_0P5 U1148 ( .A1(n631), .A2(n922), .X(n923) );
  SEN_MUXI2_S_0P5 U1149 ( .D0(n620), .D1(n628), .S(B[14]), .X(n922) );
  SEN_MUXI2_S_1 U1150 ( .D0(net58941), .D1(n1035), .S(INST[3]), .X(Z[12]) );
  SEN_ND2_S_0P5 U1151 ( .A1(net59596), .A2(net59389), .X(net59595) );
  SEN_ND2_S_1 U1152 ( .A1(n1025), .A2(n379), .X(n883) );
  SEN_OAI21_T_0P5 U1153 ( .A1(n616), .A2(A[3]), .B(n612), .X(n834) );
  SEN_ND2_S_1 U1154 ( .A1(n841), .A2(n840), .X(n842) );
  SEN_OAI21_T_0P5 U1155 ( .A1(n616), .A2(A[2]), .B(n614), .X(n843) );
  SEN_MUXI2_D_1 U1156 ( .D0(net58954), .D1(n1031), .S(INST[3]), .X(Z[6]) );
  SEN_ND2_G_1 U1157 ( .A1(net59233), .A2(n774), .X(n777) );
  SEN_ND2_2 U1158 ( .A1(n774), .A2(n773), .X(n775) );
  SEN_INV_S_1 U1159 ( .A(net59522), .X(net60246) );
  SEN_NR2_S_0P5 U1160 ( .A1(net59454), .A2(net59213), .X(net59522) );
  SEN_MUXI2_S_0P5 U1161 ( .D0(net58923), .D1(n382), .S(INST[3]), .X(Z[21]) );
  SEN_MUXI2_D_1 U1162 ( .D0(net58957), .D1(n1029), .S(INST[3]), .X(Z[5]) );
  SEN_MUXI2_S_0P5 U1163 ( .D0(n619), .D1(n628), .S(B[25]), .X(n941) );
  SEN_ND2_S_0P5 U1164 ( .A1(n395), .A2(n756), .X(net59241) );
  SEN_AOI21_T_0P5 U1165 ( .A1(net59214), .A2(net59216), .B(net59454), .X(
        net59517) );
  SEN_INV_S_1 U1166 ( .A(net59388), .X(net59598) );
  SEN_ND2_G_1 U1167 ( .A1(n832), .A2(net59221), .X(n781) );
  SEN_ND2_G_1 U1168 ( .A1(B[17]), .A2(net59988), .X(net59600) );
  SEN_MUXI2_S_1 U1169 ( .D0(net58937), .D1(n368), .S(INST[3]), .X(Z[14]) );
  SEN_MUXI2_S_1 U1170 ( .D0(net58939), .D1(n377), .S(INST[3]), .X(Z[13]) );
  SEN_INV_S_1 U1171 ( .A(n619), .X(n618) );
  SEN_INV_S_0P5 U1172 ( .A(net59300), .X(net59347) );
  SEN_NR2_S_0P5 U1173 ( .A1(n771), .A2(net59232), .X(n772) );
  SEN_MUXI2_S_1 U1174 ( .D0(n575), .D1(n716), .S(B[10]), .X(n708) );
  SEN_OAI21_T_0P5 U1175 ( .A1(n616), .A2(A[11]), .B(n613), .X(n884) );
  SEN_MUXI2_D_1 U1176 ( .D0(net58943), .D1(n366), .S(INST[3]), .X(Z[11]) );
  SEN_ND2_S_1 U1177 ( .A1(n631), .A2(n917), .X(n918) );
  SEN_ND2_S_1 U1178 ( .A1(n631), .A2(n957), .X(n958) );
  SEN_ND2_S_1 U1179 ( .A1(n631), .A2(n952), .X(n953) );
  SEN_ND2_S_1 U1180 ( .A1(n631), .A2(n930), .X(n931) );
  SEN_MUXI2_D_1 U1181 ( .D0(net58933), .D1(n365), .S(INST[3]), .X(Z[16]) );
  SEN_ND2_S_2 U1182 ( .A1(n970), .A2(n969), .X(n971) );
  SEN_INV_S_2 U1183 ( .A(n620), .X(n617) );
  SEN_BUF_1 U1184 ( .A(n602), .X(n622) );
  SEN_ND2_S_1 U1185 ( .A1(net59215), .A2(n780), .X(n785) );
  SEN_BUF_1 U1186 ( .A(n602), .X(n620) );
  SEN_INV_S_0P5 U1187 ( .A(n782), .X(n784) );
  SEN_BUF_S_1 U1188 ( .A(n602), .X(n621) );
  SEN_BUF_1 U1189 ( .A(n602), .X(n619) );
  SEN_INV_S_0P5 U1190 ( .A(n837), .X(n629) );
  SEN_INV_S_0P5 U1191 ( .A(n831), .X(n788) );
  SEN_EN2_0P5 U1192 ( .A1(net59279), .A2(net59280), .X(net59271) );
  SEN_EN2_0P5 U1195 ( .A1(n823), .A2(n822), .X(net59285) );
  SEN_AOI21_G_1 U1196 ( .A1(n788), .A2(n787), .B(n786), .X(n789) );
  SEN_INV_S_0P5 U1197 ( .A(n615), .X(n612) );
  SEN_INV_S_0P5 U1198 ( .A(n615), .X(n613) );
  SEN_NR3_1 U1199 ( .A1(n928), .A2(n927), .A3(n926), .X(net58987) );
  SEN_NR3_1 U1200 ( .A1(n1020), .A2(n1019), .A3(n1018), .X(net58989) );
  SEN_INV_4 U1201 ( .A(net59410), .X(net59214) );
  SEN_ND2_S_1 U1202 ( .A1(n779), .A2(net59233), .X(n780) );
  SEN_ND3_S_1 U1203 ( .A1(n787), .A2(net58914), .A3(n781), .X(n782) );
  SEN_ND2_S_0P5 U1204 ( .A1(net59597), .A2(net59252), .X(net59380) );
  SEN_ND4_S_1 U1205 ( .A1(n366), .A2(n381), .A3(n369), .A4(n1034), .X(n928) );
  SEN_ND4_S_1 U1206 ( .A1(n383), .A2(n367), .A3(n372), .A4(n365), .X(n1020) );
  SEN_ND3_1 U1207 ( .A1(net59238), .A2(net59498), .A3(net59503), .X(n778) );
  SEN_INV_S_0P5 U1208 ( .A(net59422), .X(net59419) );
  SEN_INV_S_0P5 U1209 ( .A(n387), .X(n632) );
  SEN_NR2_S_1 U1210 ( .A1(n1021), .A2(n1023), .X(n882) );
  SEN_OR3B_0P5 U1211 ( .B1(n830), .B2(net58913), .A(n781), .X(net59454) );
  SEN_NR2_S_1 U1212 ( .A1(n1026), .A2(n1028), .X(n880) );
  SEN_NR2_S_1 U1213 ( .A1(n1030), .A2(n1032), .X(n881) );
  SEN_ND2_S_1 U1214 ( .A1(n376), .A2(n368), .X(n926) );
  SEN_ND2_S_1 U1215 ( .A1(n1037), .A2(n378), .X(n1018) );
  SEN_ND2_S_1 U1216 ( .A1(n377), .A2(n1035), .X(n927) );
  SEN_ND2_S_1 U1217 ( .A1(n382), .A2(n1036), .X(n1019) );
  SEN_MUXI2_S_0P5 U1218 ( .D0(net58919), .D1(n1037), .S(INST[3]), .X(Z[23]) );
  SEN_MUXI2_S_0P5 U1220 ( .D0(n575), .D1(n716), .S(B[11]), .X(n717) );
  SEN_MUXI2_S_0P5 U1221 ( .D0(net58921), .D1(n378), .S(INST[3]), .X(Z[22]) );
  SEN_MUXI2_S_0P5 U1223 ( .D0(net58925), .D1(n1036), .S(INST[3]), .X(Z[20]) );
  SEN_EO2_S_0P5 U1224 ( .A1(A[13]), .A2(net61263), .X(net59691) );
  SEN_MUXI2_D_1 U1225 ( .D0(net58951), .D1(n1033), .S(INST[3]), .X(Z[7]) );
  SEN_INV_S_0P5 U1226 ( .A(n1032), .X(n1033) );
  SEN_INV_S_0P5 U1227 ( .A(n1021), .X(n1022) );
  SEN_MUXI2_D_1 U1228 ( .D0(net58963), .D1(n1025), .S(INST[3]), .X(Z[3]) );
  SEN_MUXI2_S_0P5 U1229 ( .D0(net58927), .D1(n383), .S(INST[3]), .X(Z[19]) );
  SEN_ND2_S_1 U1230 ( .A1(n631), .A2(n986), .X(n987) );
  SEN_MUXI2_S_0P5 U1231 ( .D0(n623), .D1(n628), .S(B[17]), .X(n986) );
  SEN_ND2_S_1 U1232 ( .A1(n631), .A2(n981), .X(n982) );
  SEN_MUXI2_S_0P5 U1233 ( .D0(n623), .D1(n628), .S(B[18]), .X(n981) );
  SEN_MUXI2_S_0P5 U1234 ( .D0(n621), .D1(n628), .S(B[15]), .X(n917) );
  SEN_ND2_S_1 U1235 ( .A1(n631), .A2(n941), .X(n942) );
  SEN_ND2_S_1 U1236 ( .A1(n630), .A2(n851), .X(n852) );
  SEN_ND2_T_0P5 U1237 ( .A1(n630), .A2(n911), .X(n912) );
  SEN_MUXI2_S_0P5 U1238 ( .D0(n621), .D1(n627), .S(B[12]), .X(n911) );
  SEN_ND2_S_0P65 U1239 ( .A1(n630), .A2(n906), .X(n907) );
  SEN_MUXI2_S_0P5 U1240 ( .D0(n621), .D1(n627), .S(B[13]), .X(n906) );
  SEN_ND2_S_1 U1241 ( .A1(n859), .A2(n858), .X(n1023) );
  SEN_OAI21_T_0P5 U1242 ( .A1(n616), .A2(A[1]), .B(n614), .X(n855) );
  SEN_MUXI2_D_1 U1243 ( .D0(n850), .D1(n849), .S(B[0]), .X(n854) );
  SEN_NR3_1 U1244 ( .A1(n974), .A2(n973), .A3(n972), .X(net58988) );
  SEN_ND2_S_1 U1245 ( .A1(n371), .A2(n385), .X(n973) );
  SEN_ND4_S_1 U1246 ( .A1(n384), .A2(n1039), .A3(n370), .A4(n1038), .X(n974)
         );
  SEN_ND2_S_1 U1247 ( .A1(n874), .A2(n873), .X(n1026) );
  SEN_OAI21_T_0P5 U1248 ( .A1(n616), .A2(A[4]), .B(n613), .X(n870) );
  SEN_OAI21_T_0P5 U1249 ( .A1(n616), .A2(A[8]), .B(n613), .X(n899) );
  SEN_OAI21_T_0P5 U1250 ( .A1(n616), .A2(A[9]), .B(n613), .X(n894) );
  SEN_OAI21_T_0P5 U1251 ( .A1(n616), .A2(A[10]), .B(n613), .X(n889) );
  SEN_OAI21_T_0P5 U1252 ( .A1(n616), .A2(A[12]), .B(n613), .X(n910) );
  SEN_OAI21_T_0P5 U1253 ( .A1(n616), .A2(A[13]), .B(n613), .X(n905) );
  SEN_ND2_2 U1254 ( .A1(n768), .A2(n767), .X(net59482) );
  SEN_INV_S_0P5 U1255 ( .A(n1030), .X(n1031) );
  SEN_MUXI2_D_1 U1256 ( .D0(net58960), .D1(n1027), .S(INST[3]), .X(Z[4]) );
  SEN_INV_S_0P5 U1257 ( .A(n1026), .X(n1027) );
  SEN_INV_S_0P5 U1258 ( .A(n1023), .X(n1024) );
  SEN_INV_S_0P5 U1259 ( .A(n1028), .X(n1029) );
  SEN_OAI21_T_0P5 U1260 ( .A1(n617), .A2(A[30]), .B(n612), .X(n966) );
  SEN_OAI21_T_0P5 U1261 ( .A1(n617), .A2(A[17]), .B(n612), .X(n985) );
  SEN_OAI21_0P5 U1262 ( .A1(n617), .A2(A[24]), .B(n612), .X(n945) );
  SEN_OAI21_T_0P5 U1263 ( .A1(n617), .A2(A[18]), .B(n612), .X(n980) );
  SEN_OAI21_T_0P5 U1264 ( .A1(n617), .A2(A[25]), .B(n612), .X(n940) );
  SEN_OAI21_S_0P5 U1265 ( .A1(n617), .A2(A[26]), .B(n613), .X(n934) );
  SEN_OAI21_T_0P5 U1266 ( .A1(n617), .A2(A[19]), .B(n612), .X(n975) );
  SEN_OAI21_T_0P5 U1267 ( .A1(n617), .A2(A[27]), .B(n613), .X(n929) );
  SEN_OAI21_T_0P5 U1268 ( .A1(n617), .A2(A[14]), .B(n613), .X(n921) );
  SEN_OAI21_T_0P5 U1269 ( .A1(n617), .A2(A[15]), .B(n613), .X(n916) );
  SEN_OAI21_S_0P5 U1270 ( .A1(n617), .A2(A[28]), .B(n612), .X(n956) );
  SEN_OAI21_S_0P5 U1271 ( .A1(n617), .A2(A[29]), .B(n612), .X(n951) );
  SEN_OAI21_T_0P5 U1272 ( .A1(n618), .A2(A[22]), .B(n613), .X(n1013) );
  SEN_OAI21_T_0P5 U1273 ( .A1(n618), .A2(A[20]), .B(n612), .X(n1000) );
  SEN_OAI21_T_0P5 U1274 ( .A1(n618), .A2(A[21]), .B(n612), .X(n995) );
  SEN_OAI21_T_0P5 U1275 ( .A1(n618), .A2(A[23]), .B(n612), .X(n1006) );
  SEN_ND2_T_1 U1276 ( .A1(n631), .A2(n967), .X(n968) );
  SEN_MUXI2_S_0P5 U1277 ( .D0(n623), .D1(n628), .S(B[28]), .X(n957) );
  SEN_MUXI2_S_0P5 U1278 ( .D0(n623), .D1(n628), .S(B[29]), .X(n952) );
  SEN_ND2_S_0P65 U1279 ( .A1(n631), .A2(n935), .X(n936) );
  SEN_MUXI2_S_0P5 U1280 ( .D0(n620), .D1(n628), .S(B[26]), .X(n935) );
  SEN_ND2_S_1 U1281 ( .A1(n631), .A2(n962), .X(n963) );
  SEN_ND2_S_1 U1282 ( .A1(n631), .A2(n991), .X(n992) );
  SEN_MUXI2_S_0P5 U1283 ( .D0(n623), .D1(n628), .S(B[16]), .X(n991) );
  SEN_ND2_S_1 U1284 ( .A1(n630), .A2(n895), .X(n896) );
  SEN_MUXI2_S_0P5 U1285 ( .D0(n622), .D1(n627), .S(B[9]), .X(n895) );
  SEN_ND2_S_1 U1286 ( .A1(n630), .A2(n890), .X(n891) );
  SEN_MUXI2_S_0P5 U1287 ( .D0(n622), .D1(n627), .S(B[10]), .X(n890) );
  SEN_ND2_S_1 U1288 ( .A1(n630), .A2(n885), .X(n886) );
  SEN_MUXI2_S_0P5 U1289 ( .D0(n622), .D1(n627), .S(B[11]), .X(n885) );
  SEN_ND2_S_1 U1290 ( .A1(n631), .A2(n946), .X(n947) );
  SEN_MUXI2_S_0P5 U1291 ( .D0(n623), .D1(n628), .S(B[24]), .X(n946) );
  SEN_ND2_S_1 U1292 ( .A1(n630), .A2(n838), .X(n839) );
  SEN_MUXI2_S_0P5 U1293 ( .D0(n622), .D1(n627), .S(B[3]), .X(n838) );
  SEN_ND2_S_1 U1294 ( .A1(n630), .A2(n876), .X(n877) );
  SEN_MUXI2_S_0P5 U1295 ( .D0(n622), .D1(n627), .S(B[5]), .X(n876) );
  SEN_ND2_S_1 U1296 ( .A1(n630), .A2(n866), .X(n867) );
  SEN_MUXI2_S_0P5 U1297 ( .D0(n622), .D1(n627), .S(B[7]), .X(n866) );
  SEN_ND2_S_1 U1298 ( .A1(n631), .A2(n976), .X(n977) );
  SEN_MUXI2_S_0P5 U1299 ( .D0(n623), .D1(n628), .S(B[19]), .X(n976) );
  SEN_ND2_S_1 U1300 ( .A1(n630), .A2(n856), .X(n857) );
  SEN_MUXI2_S_0P5 U1301 ( .D0(n622), .D1(n627), .S(B[1]), .X(n856) );
  SEN_ND2_S_1 U1302 ( .A1(n630), .A2(n871), .X(n872) );
  SEN_MUXI2_S_0P5 U1303 ( .D0(n622), .D1(n627), .S(B[4]), .X(n871) );
  SEN_ND2_S_1 U1304 ( .A1(n630), .A2(n861), .X(n862) );
  SEN_MUXI2_S_0P5 U1305 ( .D0(n622), .D1(n627), .S(B[6]), .X(n861) );
  SEN_ND2_S_1 U1306 ( .A1(n630), .A2(n900), .X(n901) );
  SEN_MUXI2_S_0P5 U1307 ( .D0(n621), .D1(n627), .S(B[8]), .X(n900) );
  SEN_MUXI2_S_0P5 U1308 ( .D0(n620), .D1(n628), .S(B[27]), .X(n930) );
  SEN_ND2_T_0P5 U1309 ( .A1(n630), .A2(n844), .X(n845) );
  SEN_MUXI2_S_0P5 U1310 ( .D0(n619), .D1(n627), .S(B[2]), .X(n844) );
  SEN_ND2_S_1 U1311 ( .A1(n879), .A2(n878), .X(n1028) );
  SEN_OAI21_T_0P5 U1312 ( .A1(n616), .A2(A[5]), .B(n613), .X(n875) );
  SEN_ND2_S_1 U1313 ( .A1(n869), .A2(n868), .X(n1032) );
  SEN_OAI21_T_0P5 U1314 ( .A1(n616), .A2(A[7]), .B(n613), .X(n865) );
  SEN_ND2_S_1 U1315 ( .A1(n864), .A2(n863), .X(n1030) );
  SEN_OAI21_T_0P5 U1316 ( .A1(n616), .A2(A[6]), .B(n614), .X(n860) );
  SEN_ND2_S_1 U1317 ( .A1(n914), .A2(n913), .X(n915) );
  SEN_MUXI2_S_0P5 U1318 ( .D0(net58931), .D1(n372), .S(INST[3]), .X(Z[17]) );
  SEN_ND2_S_1 U1319 ( .A1(n1004), .A2(n1003), .X(n1005) );
  SEN_ND2_S_1 U1320 ( .A1(n903), .A2(n902), .X(n904) );
  SEN_ND2_S_1 U1321 ( .A1(n949), .A2(n948), .X(n950) );
  SEN_ND2_S_1 U1322 ( .A1(n632), .A2(n1014), .X(n1015) );
  SEN_ND2_S_1 U1323 ( .A1(n632), .A2(n996), .X(n997) );
  SEN_ND2_S_1 U1324 ( .A1(n632), .A2(n1001), .X(n1002) );
  SEN_ND2_S_1 U1325 ( .A1(n632), .A2(n1007), .X(n1008) );
  SEN_MUXI2_S_0P5 U1326 ( .D0(n622), .D1(n629), .S(B[23]), .X(n1007) );
  SEN_INV_S_2 U1327 ( .A(n939), .X(n1039) );
  SEN_ND2_S_2 U1328 ( .A1(n938), .A2(n937), .X(n939) );
  SEN_ND2_S_1 U1329 ( .A1(n1010), .A2(n1009), .X(n1011) );
  SEN_INV_S_2 U1330 ( .A(n971), .X(n1041) );
  SEN_INV_S_1 U1331 ( .A(n621), .X(n616) );
  SEN_INV_2 U1332 ( .A(n744), .X(n727) );
  SEN_OAI21_G_1 U1333 ( .A1(net59381), .A2(net59382), .B(n805), .X(net59378)
         );
  SEN_INV_S_1 U1334 ( .A(n771), .X(n774) );
  SEN_ND2_S_0P5 U1336 ( .A1(net59343), .A2(net59320), .X(n821) );
  SEN_ND2_S_0P5 U1337 ( .A1(net59215), .A2(net59216), .X(n773) );
  SEN_NR2_S_0P5 U1338 ( .A1(net59298), .A2(n807), .X(n817) );
  SEN_INV_S_0P5 U1339 ( .A(n810), .X(n813) );
  SEN_INV_S_1 U1340 ( .A(n850), .X(n625) );
  SEN_INV_S_1 U1341 ( .A(n850), .X(n624) );
  SEN_INV_S_1 U1342 ( .A(n850), .X(n626) );
  SEN_EO2_S_0P5 U1343 ( .A1(net59392), .A2(net59393), .X(net59391) );
  SEN_EO2_S_0P5 U1344 ( .A1(net59257), .A2(net59258), .X(net59256) );
  SEN_INV_S_1 U1345 ( .A(n802), .X(n760) );
  SEN_ND4B_1 U1346 ( .A(n883), .B1(n882), .B2(n881), .B3(n880), .X(net58986)
         );
  SEN_OAI31_1 U1347 ( .A1(net59410), .A2(net58914), .A3(net59513), .B(net59217), .X(n771) );
  SEN_EN2_0P5 U1348 ( .A1(n827), .A2(net59270), .X(net59261) );
  SEN_EN2_0P5 U1350 ( .A1(net59418), .A2(net59419), .X(net60465) );
  SEN_EN2_0P5 U1351 ( .A1(net59388), .A2(net59389), .X(net59376) );
  SEN_OAI21_G_1 U1352 ( .A1(net59250), .A2(net59251), .B(net59380), .X(n806)
         );
  SEN_EN2_0P5 U1353 ( .A1(n802), .A2(net59409), .X(net59396) );
  SEN_OAI22_S_1 U1354 ( .A1(net59298), .A2(net59347), .B1(net60557), .B2(
        net59299), .X(net59288) );
  SEN_EN2_0P5 U1355 ( .A1(net59315), .A2(net59316), .X(net59307) );
  SEN_INV_2 U1356 ( .A(net59241), .X(net59564) );
  SEN_INV_2 U1357 ( .A(net59251), .X(net59597) );
  SEN_INV_1 U1358 ( .A(net59267), .X(net59663) );
  SEN_ND2_G_1 U1359 ( .A1(net59433), .A2(net58985), .X(n799) );
  SEN_NR2_S_0P5 U1360 ( .A1(net60557), .A2(n808), .X(n816) );
  SEN_INV_S_0P5 U1361 ( .A(net59252), .X(net59594) );
  SEN_INV_2 U1362 ( .A(net59242), .X(net59558) );
  SEN_INV_S_2 U1363 ( .A(n823), .X(n714) );
  SEN_AN2_S_0P5 U1364 ( .A1(net59205), .A2(n833), .X(n602) );
  SEN_INV_S_1 U1365 ( .A(n387), .X(n631) );
  SEN_INV_S_1 U1366 ( .A(n835), .X(n633) );
  SEN_INV_S_1 U1367 ( .A(n835), .X(n634) );
  SEN_INV_S_1 U1368 ( .A(n615), .X(n614) );
  SEN_INV_S_1 U1369 ( .A(n835), .X(n635) );
  SEN_INV_2 U1370 ( .A(n1012), .X(n615) );
  SEN_ND2_S_0P5 U1371 ( .A1(B[24]), .A2(net59990), .X(net59530) );
  SEN_MUXI2_S_0P5 U1372 ( .D0(n396), .D1(n794), .S(B[25]), .X(net59531) );
  SEN_MUXI2_S_0P5 U1373 ( .D0(n793), .D1(n792), .S(B[30]), .X(net59470) );
  SEN_ND2_S_0P5 U1374 ( .A1(B[25]), .A2(net59990), .X(n770) );
  SEN_MUXI2_S_0P5 U1375 ( .D0(n396), .D1(n591), .S(B[26]), .X(n769) );
  SEN_ND2_S_0P5 U1376 ( .A1(B[8]), .A2(net59469), .X(n711) );
  SEN_EO2_S_0P5 U1377 ( .A1(A[23]), .A2(net59978), .X(net59538) );
  SEN_MUXI2_S_2 U1379 ( .D0(n575), .D1(n716), .S(B[6]), .X(net59755) );
  SEN_EO2_S_0P5 U1380 ( .A1(A[25]), .A2(net59976), .X(net59523) );
  SEN_AN2_S_0P5 U1381 ( .A1(B[20]), .A2(net59988), .X(n603) );
  SEN_MUX2_DG_1 U1382 ( .D0(n575), .D1(n794), .S(B[21]), .X(n604) );
  SEN_AN2_S_0P5 U1384 ( .A1(B[12]), .A2(net59988), .X(net60380) );
  SEN_ND2_S_0P5 U1385 ( .A1(B[11]), .A2(net59990), .X(net59714) );
  SEN_ND2_S_0P5 U1386 ( .A1(B[23]), .A2(net59988), .X(net59536) );
  SEN_MUXI2_S_0P5 U1387 ( .D0(n396), .D1(n591), .S(B[24]), .X(net59537) );
  SEN_ND2_S_0P5 U1388 ( .A1(B[21]), .A2(net59990), .X(n758) );
  SEN_MUXI2_S_0P5 U1389 ( .D0(n396), .D1(n794), .S(B[22]), .X(n757) );
  SEN_ND2_S_0P5 U1390 ( .A1(n394), .A2(n640), .X(net59431) );
  SEN_EO2_S_0P5 U1391 ( .A1(A[31]), .A2(net59978), .X(n640) );
  SEN_ND2_S_0P5 U1392 ( .A1(B[15]), .A2(net59990), .X(net59605) );
  SEN_MUXI2_S_0P5 U1393 ( .D0(n396), .D1(n794), .S(B[16]), .X(net59606) );
  SEN_ND2_S_0P5 U1394 ( .A1(B[6]), .A2(net59988), .X(n696) );
  SEN_MUXI2_S_0P5 U1395 ( .D0(n575), .D1(n794), .S(B[7]), .X(n695) );
  SEN_ND2_S_0P5 U1396 ( .A1(net59958), .A2(n765), .X(net58913) );
  SEN_EO2_S_0P5 U1397 ( .A1(A[26]), .A2(net59976), .X(n765) );
  SEN_ND2_S_0P5 U1398 ( .A1(B[28]), .A2(net59988), .X(net59465) );
  SEN_MUXI2_S_0P5 U1399 ( .D0(n396), .D1(n591), .S(B[29]), .X(net59466) );
  SEN_MUXI2_D_1 U1400 ( .D0(net58949), .D1(n1034), .S(INST[3]), .X(Z[8]) );
  SEN_AN2_S_0P5 U1401 ( .A1(B[19]), .A2(net59988), .X(net60377) );
  SEN_MUX2_DG_1 U1402 ( .D0(n396), .D1(n794), .S(B[20]), .X(net60378) );
  SEN_AN2_S_0P5 U1403 ( .A1(B[18]), .A2(net59988), .X(net60375) );
  SEN_MUX2_DG_1 U1404 ( .D0(n396), .D1(n794), .S(B[19]), .X(net60376) );
  SEN_MUXI2_S_1 U1405 ( .D0(n624), .D1(n875), .S(B[5]), .X(n879) );
  SEN_MUXI2_S_1 U1406 ( .D0(n633), .D1(n877), .S(A[5]), .X(n878) );
  SEN_MUXI2_S_1 U1407 ( .D0(n624), .D1(n870), .S(B[4]), .X(n874) );
  SEN_MUXI2_S_1 U1408 ( .D0(n633), .D1(n872), .S(A[4]), .X(n873) );
  SEN_MUXI2_S_1 U1409 ( .D0(n624), .D1(n865), .S(B[7]), .X(n869) );
  SEN_MUXI2_S_1 U1410 ( .D0(n633), .D1(n867), .S(A[7]), .X(n868) );
  SEN_MUXI2_S_1 U1411 ( .D0(n624), .D1(n860), .S(B[6]), .X(n864) );
  SEN_MUXI2_S_1 U1412 ( .D0(n633), .D1(n862), .S(A[6]), .X(n863) );
  SEN_MUXI2_S_1 U1413 ( .D0(n624), .D1(n855), .S(B[1]), .X(n859) );
  SEN_MUXI2_S_1 U1414 ( .D0(n633), .D1(n857), .S(A[1]), .X(n858) );
  SEN_MUXI2_S_0P5 U1415 ( .D0(net58970), .D1(n1022), .S(INST[3]), .X(Z[0]) );
  SEN_AN2_S_0P5 U1416 ( .A1(B[14]), .A2(net59990), .X(net60372) );
  SEN_MUX2_DG_1 U1417 ( .D0(n396), .D1(n794), .S(B[15]), .X(net60373) );
  SEN_ND2_S_0P5 U1418 ( .A1(B[7]), .A2(net59990), .X(n722) );
  SEN_MUXI2_S_0P5 U1419 ( .D0(n575), .D1(n794), .S(B[8]), .X(n721) );
  SEN_ND2_S_0P5 U1421 ( .A1(n394), .A2(n641), .X(net59232) );
  SEN_EO2_S_0P5 U1422 ( .A1(A[24]), .A2(net61241), .X(n641) );
  SEN_ND2_S_0P5 U1423 ( .A1(B[22]), .A2(net59990), .X(n762) );
  SEN_MUXI2_S_0P5 U1424 ( .D0(n396), .D1(n794), .S(B[23]), .X(n761) );
  SEN_ND2_S_0P5 U1425 ( .A1(B[13]), .A2(net59990), .X(net59630) );
  SEN_MUXI2_S_0P5 U1426 ( .D0(n575), .D1(n794), .S(B[14]), .X(net59631) );
  SEN_MUXI2_S_0P5 U1427 ( .D0(net58967), .D1(n1024), .S(INST[3]), .X(Z[1]) );
  SEN_ND2_S_0P5 U1428 ( .A1(n395), .A2(n796), .X(net59418) );
  SEN_EO2_S_0P5 U1429 ( .A1(A[29]), .A2(net59978), .X(n796) );
  SEN_EO2_S_0P5 U1430 ( .A1(A[20]), .A2(net61246), .X(net59560) );
  SEN_ND2_S_0P5 U1431 ( .A1(B[26]), .A2(net59988), .X(n768) );
  SEN_MUXI2_S_0P5 U1432 ( .D0(n396), .D1(n591), .S(B[27]), .X(n767) );
  SEN_MUXI2_S_0P5 U1433 ( .D0(net58965), .D1(n379), .S(INST[3]), .X(Z[2]) );
  SEN_ND2_G_1 U1434 ( .A1(n764), .A2(n763), .X(n787) );
  SEN_ND2_S_0P5 U1435 ( .A1(B[27]), .A2(net59988), .X(n764) );
  SEN_MUXI2_S_0P5 U1436 ( .D0(n396), .D1(n591), .S(B[28]), .X(n763) );
  SEN_ND2_S_0P5 U1437 ( .A1(n395), .A2(n798), .X(net59429) );
  SEN_EO2_S_0P5 U1438 ( .A1(A[14]), .A2(net61263), .X(net59616) );
  SEN_ND2_G_1 U1439 ( .A1(n639), .A2(n638), .X(net59433) );
  SEN_ND3_S_0P5 U1440 ( .A1(n637), .A2(n606), .A3(n663), .X(n639) );
  SEN_EN2_0P5 U1441 ( .A1(N72), .A2(n636), .X(n637) );
  SEN_EO2_S_0P5 U1442 ( .A1(A[19]), .A2(net61263), .X(net59575) );
  SEN_ND3B_1 U1443 ( .A(INST[1]), .B1(N72), .B2(INST[2]), .X(n835) );
  SEN_NR2B_V1DG_1 U1444 ( .A(n394), .B(n605), .X(net60361) );
  SEN_EN2_0P5 U1445 ( .A1(A[28]), .A2(net59444), .X(n605) );
  SEN_ND2_S_0P5 U1446 ( .A1(n394), .A2(n759), .X(n802) );
  SEN_EO2_S_0P5 U1447 ( .A1(A[22]), .A2(net61263), .X(n759) );
  SEN_ND2_S_0P5 U1448 ( .A1(n395), .A2(n755), .X(net59388) );
  SEN_ND3_S_0P5 U1450 ( .A1(INST[3]), .A2(n386), .A3(n1041), .X(n972) );
  SEN_OR3B_0P5 U1451 ( .B1(n590), .B2(n854), .A(n853), .X(n1021) );
  SEN_MUXI2_S_1 U1452 ( .D0(n633), .D1(n852), .S(A[0]), .X(n853) );
  SEN_AOI21B_1 U1453 ( .A1(n848), .A2(n619), .B(n614), .X(n849) );
  SEN_OAI21_G_1 U1454 ( .A1(n618), .A2(A[16]), .B(n612), .X(n990) );
  SEN_OR2_DG_1 U1455 ( .A1(n667), .A2(INST[3]), .X(n606) );
  SEN_INV_S_1 U1456 ( .A(n950), .X(n1038) );
  SEN_MUXI2_S_1 U1457 ( .D0(n625), .D1(n945), .S(B[24]), .X(n949) );
  SEN_MUXI2_S_1 U1458 ( .D0(n634), .D1(n947), .S(A[24]), .X(n948) );
  SEN_MUXI2_S_1 U1459 ( .D0(n625), .D1(n990), .S(B[16]), .X(n994) );
  SEN_MUXI2_S_1 U1460 ( .D0(n634), .D1(n992), .S(A[16]), .X(n993) );
  SEN_INV_S_1 U1461 ( .A(n904), .X(n1034) );
  SEN_MUXI2_S_1 U1462 ( .D0(n624), .D1(n899), .S(B[8]), .X(n903) );
  SEN_MUXI2_S_1 U1463 ( .D0(n633), .D1(n901), .S(A[8]), .X(n902) );
  SEN_MUXI2_S_1 U1464 ( .D0(n624), .D1(n843), .S(B[2]), .X(n847) );
  SEN_MUXI2_S_1 U1465 ( .D0(n633), .D1(n845), .S(A[2]), .X(n846) );
  SEN_MUXI2_S_1 U1466 ( .D0(n626), .D1(n1013), .S(B[22]), .X(n1017) );
  SEN_MUXI2_S_1 U1467 ( .D0(n635), .D1(n1015), .S(A[22]), .X(n1016) );
  SEN_INV_S_1 U1468 ( .A(n1005), .X(n1036) );
  SEN_MUXI2_S_1 U1469 ( .D0(n626), .D1(n1000), .S(B[20]), .X(n1004) );
  SEN_MUXI2_S_1 U1470 ( .D0(n635), .D1(n1002), .S(A[20]), .X(n1003) );
  SEN_MUXI2_S_1 U1471 ( .D0(n625), .D1(n921), .S(B[14]), .X(n925) );
  SEN_MUXI2_S_1 U1472 ( .D0(n634), .D1(n923), .S(A[14]), .X(n924) );
  SEN_INV_S_1 U1473 ( .A(n915), .X(n1035) );
  SEN_MUXI2_S_1 U1474 ( .D0(n624), .D1(n910), .S(B[12]), .X(n914) );
  SEN_MUXI2_S_1 U1475 ( .D0(n633), .D1(n912), .S(A[12]), .X(n913) );
  SEN_INV_S_1 U1476 ( .A(n842), .X(n1025) );
  SEN_MUXI2_S_1 U1477 ( .D0(n624), .D1(n834), .S(B[3]), .X(n841) );
  SEN_MUXI2_S_1 U1478 ( .D0(n633), .D1(n839), .S(A[3]), .X(n840) );
  SEN_INV_S_1 U1479 ( .A(n1011), .X(n1037) );
  SEN_MUXI2_S_1 U1480 ( .D0(n626), .D1(n1006), .S(B[23]), .X(n1010) );
  SEN_MUXI2_S_1 U1481 ( .D0(n635), .D1(n1008), .S(A[23]), .X(n1009) );
  SEN_MUXI2_S_1 U1482 ( .D0(n625), .D1(n995), .S(B[21]), .X(n999) );
  SEN_MUXI2_S_1 U1483 ( .D0(n635), .D1(n997), .S(A[21]), .X(n998) );
  SEN_MUXI2_S_1 U1484 ( .D0(n624), .D1(n916), .S(B[15]), .X(n920) );
  SEN_MUXI2_S_1 U1485 ( .D0(n634), .D1(n918), .S(A[15]), .X(n919) );
  SEN_MUXI2_S_1 U1486 ( .D0(n624), .D1(n905), .S(B[13]), .X(n909) );
  SEN_MUXI2_S_1 U1487 ( .D0(n633), .D1(n907), .S(A[13]), .X(n908) );
  SEN_MUXI2_S_1 U1488 ( .D0(n625), .D1(n934), .S(B[26]), .X(n938) );
  SEN_MUXI2_S_1 U1489 ( .D0(n634), .D1(n936), .S(A[26]), .X(n937) );
  SEN_MUXI2_S_1 U1490 ( .D0(n625), .D1(n980), .S(B[18]), .X(n984) );
  SEN_MUXI2_S_1 U1491 ( .D0(n634), .D1(n982), .S(A[18]), .X(n983) );
  SEN_MUXI2_S_1 U1492 ( .D0(n624), .D1(n889), .S(B[10]), .X(n893) );
  SEN_MUXI2_S_1 U1493 ( .D0(n633), .D1(n891), .S(A[10]), .X(n892) );
  SEN_MUXI2_S_1 U1494 ( .D0(n623), .D1(n628), .S(B[30]), .X(n967) );
  SEN_MUXI2_S_1 U1495 ( .D0(n620), .D1(n629), .S(B[22]), .X(n1014) );
  SEN_MUXI2_S_1 U1496 ( .D0(n622), .D1(n629), .S(B[21]), .X(n996) );
  SEN_MUXI2_S_1 U1497 ( .D0(n622), .D1(n629), .S(B[20]), .X(n1001) );
  SEN_MUXI2_S_1 U1498 ( .D0(n619), .D1(n627), .S(B[0]), .X(n851) );
  SEN_ND2_G_1 U1499 ( .A1(B[31]), .A2(INST[1]), .X(n636) );
  SEN_MUXI2_S_1 U1500 ( .D0(n625), .D1(n940), .S(B[25]), .X(n944) );
  SEN_MUXI2_S_1 U1501 ( .D0(n634), .D1(n942), .S(A[25]), .X(n943) );
  SEN_MUXI2_S_1 U1502 ( .D0(n625), .D1(n929), .S(B[27]), .X(n933) );
  SEN_MUXI2_S_1 U1503 ( .D0(n634), .D1(n931), .S(A[27]), .X(n932) );
  SEN_MUXI2_S_1 U1504 ( .D0(n625), .D1(n985), .S(B[17]), .X(n989) );
  SEN_MUXI2_S_1 U1505 ( .D0(n634), .D1(n987), .S(A[17]), .X(n988) );
  SEN_MUXI2_S_1 U1506 ( .D0(n625), .D1(n975), .S(B[19]), .X(n979) );
  SEN_MUXI2_S_1 U1507 ( .D0(n634), .D1(n977), .S(A[19]), .X(n978) );
  SEN_MUXI2_S_1 U1508 ( .D0(n624), .D1(n894), .S(B[9]), .X(n898) );
  SEN_MUXI2_S_1 U1509 ( .D0(n633), .D1(n896), .S(A[9]), .X(n897) );
  SEN_MUXI2_S_1 U1510 ( .D0(n624), .D1(n884), .S(B[11]), .X(n888) );
  SEN_MUXI2_S_1 U1511 ( .D0(n633), .D1(n886), .S(A[11]), .X(n887) );
  SEN_MUXI2_S_1 U1512 ( .D0(n625), .D1(n966), .S(B[30]), .X(n970) );
  SEN_MUXI2_S_1 U1513 ( .D0(n634), .D1(n968), .S(A[30]), .X(n969) );
  SEN_MUXI2_S_1 U1514 ( .D0(n625), .D1(n956), .S(B[28]), .X(n960) );
  SEN_MUXI2_S_1 U1515 ( .D0(n634), .D1(n958), .S(A[28]), .X(n959) );
  SEN_MUXI2_S_1 U1516 ( .D0(n625), .D1(n951), .S(B[29]), .X(n955) );
  SEN_MUXI2_S_1 U1517 ( .D0(n634), .D1(n953), .S(A[29]), .X(n954) );
  SEN_INV_S_1 U1518 ( .A(A[0]), .X(n848) );
  SEN_TIE0_1 U1519 ( .X(\*Logic0* ) );
  SEN_ND2B_S_0P5 U1520 ( .A(n447), .B(net59395), .X(net59390) );
  SEN_MUXI2_S_1 U1521 ( .D0(n634), .D1(n963), .S(A[31]), .X(n964) );
  SEN_OAI21_G_1 U1522 ( .A1(n617), .A2(A[31]), .B(n612), .X(n961) );
  SEN_EN2_S_1 U1524 ( .A1(net59430), .A2(\FLAGS[1] ), .X(FLAGS[0]) );
  SEN_ND2B_S_0P5 U1525 ( .A(net59870), .B(B[30]), .X(n638) );
  SEN_OAI211_8 U1526 ( .A1(net59231), .A2(n777), .B1(n776), .B2(n775), .X(
        net59461) );
  SEN_ND2_4 U1527 ( .A1(B[3]), .A2(net59469), .X(n649) );
  SEN_ND2_4 U1528 ( .A1(n669), .A2(n650), .X(n661) );
  SEN_INV_S_3 U1529 ( .A(net59299), .X(net59671) );
  SEN_EO2_3 U1530 ( .A1(A[17]), .A2(net61246), .X(n752) );
  SEN_EO2_3 U1531 ( .A1(A[21]), .A2(net61241), .X(n756) );
  SEN_ND2_4 U1532 ( .A1(n758), .A2(n757), .X(net59409) );
  SEN_ND2_T_4 U419 ( .A1(net59727), .A2(net59677), .X(net59729) );
  SEN_AO21B_4 U420 ( .A1(net59689), .A2(n1050), .B(net59688), .X(net59341) );
  SEN_INV_S_4 U423 ( .A(n528), .X(n435) );
  SEN_AOAI211_1 U424 ( .A1(n813), .A2(net59362), .B(n812), .C(n822), .X(n814)
         );
  SEN_OAI21_S_0P5 U425 ( .A1(net60557), .A2(n811), .B(n824), .X(n812) );
  SEN_OAI21_G_4 U427 ( .A1(n414), .A2(net59750), .B(n475), .X(n1044) );
  SEN_OAI21_S_3 U431 ( .A1(n414), .A2(net59750), .B(n475), .X(n444) );
  SEN_INV_2 U432 ( .A(net59315), .X(n475) );
  SEN_INV_1P25 U433 ( .A(net59343), .X(n1045) );
  SEN_BUF_1 U434 ( .A(net59322), .X(n1061) );
  SEN_INV_3 U435 ( .A(net60983), .X(n1077) );
  SEN_INV_S_4 U436 ( .A(net59690), .X(net59758) );
  SEN_INV_S_3 U445 ( .A(net59873), .X(n1058) );
  SEN_OAI21_G_4 U446 ( .A1(n647), .A2(n589), .B(n649), .X(n440) );
  SEN_ND2B_V1_8 U450 ( .A(n354), .B(n409), .X(n412) );
  SEN_ND2_6 U451 ( .A1(n417), .A2(n1060), .X(n361) );
  SEN_AOI21_3 U458 ( .A1(n567), .A2(n450), .B(n1068), .X(n449) );
  SEN_OR2_10 U463 ( .A1(net59343), .A2(net59687), .X(net60219) );
  SEN_ND2_2 U464 ( .A1(net59690), .A2(net59316), .X(n472) );
  SEN_ND3_T_4 U470 ( .A1(n1046), .A2(A[31]), .A3(INST[1]), .X(n654) );
  SEN_INV_32 U471 ( .A(B[31]), .X(n1046) );
  SEN_EN2_5 U472 ( .A1(A[3]), .A2(net59980), .X(n646) );
  SEN_INV_16 U473 ( .A(net59980), .X(net59978) );
  SEN_ND2_T_3 U477 ( .A1(n412), .A2(n673), .X(n699) );
  SEN_AN2_S_1P5 U479 ( .A1(net59687), .A2(net59343), .X(n407) );
  SEN_INV_12 U480 ( .A(net59322), .X(net59343) );
  SEN_OR3_4 U484 ( .A1(net59333), .A2(n460), .A3(n411), .X(n391) );
  SEN_AN2_S_16 U490 ( .A1(n464), .A2(INST[2]), .X(n468) );
  SEN_INV_0P65 U492 ( .A(n733), .X(n1047) );
  SEN_INV_3 U493 ( .A(n730), .X(n733) );
  SEN_OAI31_2 U495 ( .A1(net59267), .A2(net59700), .A3(net59270), .B(n725), 
        .X(n730) );
  SEN_ND2_6 U497 ( .A1(n1077), .A2(net59748), .X(net59310) );
  SEN_AOI21B_3 U498 ( .A1(net59744), .A2(net59743), .B(net60218), .X(n700) );
  SEN_AOAI211_4 U501 ( .A1(n660), .A2(n661), .B(n659), .C(n456), .X(n443) );
  SEN_INV_S_6 U503 ( .A(net59819), .X(n1056) );
  SEN_NR2_T_2 U504 ( .A1(net59779), .A2(net60219), .X(n1048) );
  SEN_NR2_T_2 U505 ( .A1(net59779), .A2(net60219), .X(net60218) );
  SEN_NR2_G_4 U507 ( .A1(net59779), .A2(n594), .X(net59748) );
  SEN_ND2_3 U510 ( .A1(net59304), .A2(n375), .X(n743) );
  SEN_OAI21_T_4 U512 ( .A1(n521), .A2(n525), .B(n526), .X(n524) );
  SEN_ND2_T_4 U514 ( .A1(n412), .A2(net59793), .X(net59776) );
  SEN_EO2_8 U516 ( .A1(n1054), .A2(n1059), .X(n647) );
  SEN_OR2_3 U520 ( .A1(n581), .A2(n582), .X(net59326) );
  SEN_INV_S_0P5 U523 ( .A(net59336), .X(n1049) );
  SEN_INV_2 U524 ( .A(n1049), .X(n1050) );
  SEN_ND2_T_6 U526 ( .A1(n683), .A2(n682), .X(net59336) );
  SEN_OAOI211_3 U527 ( .A1(n572), .A2(n522), .B(n523), .C(n524), .X(net41954)
         );
  SEN_MUXI2_DG_0P75 U530 ( .D0(net58915), .D1(n370), .S(INST[3]), .X(Z[25]) );
  SEN_EO2_8 U531 ( .A1(n1051), .A2(n527), .X(n521) );
  SEN_INV_32 U532 ( .A(n363), .X(n1051) );
  SEN_OR2_2 U533 ( .A1(n1052), .A2(net59992), .X(n718) );
  SEN_INV_32 U534 ( .A(B[10]), .X(n1052) );
  SEN_INV_5 U535 ( .A(net59992), .X(net59988) );
  SEN_INV_S_4 U536 ( .A(net59469), .X(net59992) );
  SEN_INV_4 U537 ( .A(net59375), .X(net59678) );
  SEN_AN2_DG_2 U538 ( .A1(net59346), .A2(net59306), .X(n374) );
  SEN_ND2_2 U543 ( .A1(n696), .A2(n695), .X(net59346) );
  SEN_ND2_T_1P5 U544 ( .A1(B[2]), .A2(net59469), .X(n644) );
  SEN_EN3_DG_2 U545 ( .A1(net59325), .A2(net59326), .A3(net59327), .X(net58970) );
  SEN_AOI22_0P5 U546 ( .A1(net59326), .A2(net59327), .B1(net59325), .B2(
        net59332), .X(net59328) );
  SEN_ND2_T_2 U548 ( .A1(n690), .A2(n689), .X(net59327) );
  SEN_INV_2 U549 ( .A(net59624), .X(n1076) );
  SEN_AN2_5 U551 ( .A1(net59679), .A2(net59680), .X(n1053) );
  SEN_INV_2 U552 ( .A(net59336), .X(net59687) );
  SEN_INV_32 U557 ( .A(A[4]), .X(n1054) );
  SEN_ND2_T_4 U558 ( .A1(n1058), .A2(A[0]), .X(n592) );
  SEN_ND2_S_2 U559 ( .A1(n611), .A2(n693), .X(n675) );
  SEN_ND2B_V1_6 U560 ( .A(n653), .B(n654), .X(n693) );
  SEN_INV_16 U561 ( .A(n645), .X(n716) );
  SEN_INV_S_3 U563 ( .A(n699), .X(n579) );
  SEN_EO2_8 U567 ( .A1(A[1]), .A2(n468), .X(n1055) );
  SEN_BUF_D_1 U568 ( .A(n460), .X(n410) );
  SEN_NR2_G_4 U569 ( .A1(n460), .A2(n411), .X(n409) );
  SEN_OR4_4 U570 ( .A1(net59427), .A2(n432), .A3(n433), .A4(n434), .X(net59437) );
  SEN_ND3_6 U571 ( .A1(n402), .A2(INST[2]), .A3(INST[1]), .X(n667) );
  SEN_INV_24 U572 ( .A(N72), .X(n402) );
  SEN_ND2_16 U573 ( .A1(n574), .A2(n642), .X(n645) );
  SEN_NR2_6 U575 ( .A1(n518), .A2(net60540), .X(n508) );
  SEN_ND2_T_5 U576 ( .A1(n598), .A2(n750), .X(net59639) );
  SEN_EO2_5 U578 ( .A1(net61884), .A2(net60465), .X(net58902) );
  SEN_ND2_4 U585 ( .A1(net59426), .A2(net59425), .X(net61884) );
  SEN_INV_10 U589 ( .A(net59799), .X(net59819) );
  SEN_INV_12 U590 ( .A(B[31]), .X(n458) );
  SEN_AOI22_4 U591 ( .A1(n703), .A2(n1060), .B1(net59335), .B2(net59343), .X(
        n705) );
  SEN_INV_S_32 U592 ( .A(A[31]), .X(n469) );
  SEN_EO3_2 U594 ( .A1(n441), .A2(net59305), .A3(net59306), .X(net58954) );
  SEN_INV_AS_3 U598 ( .A(net59642), .X(net60873) );
  SEN_AOI21_T_1 U599 ( .A1(net59242), .A2(net59398), .B(n804), .X(net59397) );
  SEN_BUF_D_1 U607 ( .A(net59349), .X(n353) );
  SEN_OAI21_S_2 U611 ( .A1(net59401), .A2(net59402), .B(n803), .X(net59398) );
  SEN_BUF_S_2 U613 ( .A(net59247), .X(n1057) );
  SEN_AOAI211_4 U615 ( .A1(net59216), .A2(n561), .B(n562), .C(n563), .X(n556)
         );
  SEN_INV_5 U616 ( .A(net59434), .X(net59430) );
  SEN_ND2_T_2 U617 ( .A1(net59237), .A2(net59497), .X(net59490) );
  SEN_OAI21_4 U618 ( .A1(net59349), .A2(net59351), .B(net59382), .X(net59385)
         );
  SEN_AOAI211_8 U619 ( .A1(net59541), .A2(net59542), .B(net59543), .C(net59544), .X(net59533) );
  SEN_NR2_T_5 U620 ( .A1(n451), .A2(net59405), .X(net59541) );
  SEN_AOAI211_6 U624 ( .A1(n487), .A2(net59393), .B(n488), .C(n486), .X(
        net59544) );
  SEN_ND2B_V1DG_4 U625 ( .A(n648), .B(n436), .X(net60861) );
  SEN_ND2B_S_4 U627 ( .A(n820), .B(n819), .X(net59309) );
  SEN_ND2_G_3 U629 ( .A1(n649), .A2(n686), .X(n819) );
  SEN_EO2_S_1 U631 ( .A1(n820), .A2(n819), .X(net59338) );
  SEN_INV_S_3 U632 ( .A(net59873), .X(n1059) );
  SEN_INV_4 U633 ( .A(net59873), .X(net59444) );
  SEN_INV_S_6 U634 ( .A(net61240), .X(net61241) );
  SEN_INV_4 U635 ( .A(net61245), .X(net59976) );
  SEN_INV_3 U640 ( .A(net61262), .X(net61263) );
  SEN_INV_3 U642 ( .A(net59978), .X(net61240) );
  SEN_AN2_6 U645 ( .A1(n391), .A2(n673), .X(n1060) );
  SEN_ND2_4 U646 ( .A1(n435), .A2(net61810), .X(net59434) );
  SEN_INV_4 U647 ( .A(n440), .X(n436) );
  SEN_EN2_5 U648 ( .A1(n662), .A2(N72), .X(n390) );
  SEN_ND2_T_8 U651 ( .A1(net59725), .A2(n474), .X(net59654) );
  SEN_ND2B_3 U652 ( .A(net59427), .B(net59425), .X(net59416) );
  SEN_AOAI211_4 U653 ( .A1(net59237), .A2(net59503), .B(net59238), .C(net59535), .X(net59456) );
  SEN_EN2_S_3 U654 ( .A1(net59412), .A2(net59223), .X(net58908) );
  SEN_MUXI2_DG_1 U655 ( .D0(net58908), .D1(n384), .S(INST[3]), .X(Z[27]) );
  SEN_EN2_S_3 U657 ( .A1(n453), .A2(n1063), .X(net58904) );
  SEN_NR3_T_6 U658 ( .A1(n347), .A2(n348), .A3(n349), .X(n1063) );
  SEN_AOI21B_3 U660 ( .A1(net59490), .A2(n439), .B(net59215), .X(n355) );
  SEN_ND2_T_4 U665 ( .A1(n573), .A2(net59440), .X(net59427) );
  SEN_EN3_1 U666 ( .A1(net58912), .A2(net58913), .A3(net58914), .X(n1040) );
  SEN_INV_0P8 U668 ( .A(net59211), .X(net58912) );
  SEN_ND2_T_6 U670 ( .A1(n1055), .A2(n389), .X(n460) );
  SEN_AOAI211_6 U671 ( .A1(net58984), .A2(net59431), .B(net59430), .C(n799), 
        .X(\FLAGS[1] ) );
  SEN_AOAI211_6 U672 ( .A1(net59205), .A2(N72), .B(INST[1]), .C(n671), .X(n672) );
  SEN_INV_32 U674 ( .A(INST[2]), .X(net59205) );
  SEN_ND3_T_8 U676 ( .A1(n402), .A2(n415), .A3(INST[2]), .X(n671) );
  SEN_ND2_G_4 U677 ( .A1(n676), .A2(n674), .X(n690) );
  SEN_AOI31_T_8 U678 ( .A1(N72), .A2(B[0]), .A3(INST[1]), .B(n670), .X(n674)
         );
  SEN_INV_4 U680 ( .A(n672), .X(n676) );
  SEN_AOI21_T_8 U682 ( .A1(n658), .A2(n657), .B(n609), .X(n691) );
  SEN_OAI21_T_8 U686 ( .A1(n656), .A2(n607), .B(n655), .X(n609) );
  SEN_ND2_6 U687 ( .A1(n664), .A2(n663), .X(n685) );
  SEN_ND2B_S_12 U692 ( .A(INST[1]), .B(INST[2]), .X(n663) );
  SEN_ND2_T_6 U699 ( .A1(A[9]), .A2(net59980), .X(n587) );
  SEN_NR2_G_2 U711 ( .A1(n745), .A2(n744), .X(n748) );
  SEN_INV_1P5 U718 ( .A(n745), .X(n736) );
  SEN_ND2_T_8 U722 ( .A1(n809), .A2(n828), .X(n745) );
  SEN_ND2_4 U738 ( .A1(net59773), .A2(n694), .X(n673) );
  SEN_NR2_S_3 U758 ( .A1(net59739), .A2(n1045), .X(n703) );
  SEN_AOAI211_6 U764 ( .A1(n661), .A2(n660), .B(n659), .C(n456), .X(net59332)
         );
  SEN_OAI31_4 U769 ( .A1(net59849), .A2(DI[31]), .A3(INST[3]), .B(n652), .X(
        n659) );
  SEN_INV_S_8 U786 ( .A(net61245), .X(net61246) );
  SEN_AN2_4 U787 ( .A1(net59799), .A2(net59962), .X(n419) );
  SEN_AOI22_0P5 U788 ( .A1(n1061), .A2(net59341), .B1(net59342), .B2(n821), 
        .X(net59337) );
  SEN_NR2_2 U789 ( .A1(n693), .A2(n692), .X(n581) );
  SEN_INV_4 U795 ( .A(n692), .X(n678) );
  SEN_EO2_3 U798 ( .A1(A[2]), .A2(n1059), .X(net59794) );
  SEN_EO2_0P5 U802 ( .A1(A[18]), .A2(net59976), .X(n755) );
  SEN_INV_6 U803 ( .A(net59978), .X(net61245) );
  SEN_INV_S_3 U808 ( .A(net59978), .X(net61262) );
  SEN_EO2_3 U809 ( .A1(A[4]), .A2(net59444), .X(n406) );
  SEN_NR2_T_8 U810 ( .A1(net60205), .A2(n397), .X(net59781) );
  SEN_INV_S_6 U812 ( .A(net59739), .X(n417) );
  SEN_ND2_8 U813 ( .A1(net61326), .A2(net59793), .X(net59739) );
  SEN_NR2_S_4 U816 ( .A1(n745), .A2(n740), .X(n741) );
  SEN_ND2_T_2 U819 ( .A1(net59799), .A2(n674), .X(n1062) );
  SEN_BUF_S_2 U820 ( .A(n1056), .X(n401) );
  SEN_ND2_G_3 U821 ( .A1(net59456), .A2(net59457), .X(net60751) );
  SEN_EN2_1 U823 ( .A1(net60464), .A2(net59421), .X(n1042) );
  SEN_EO2_2 U826 ( .A1(net60464), .A2(net59421), .X(n572) );
  SEN_ND4_S_6 U829 ( .A1(net58904), .A2(net58902), .A3(n359), .A4(n529), .X(
        n522) );
  SEN_INV_3 U833 ( .A(net59425), .X(n433) );
  SEN_ND2_4 U840 ( .A1(n566), .A2(net59517), .X(net59425) );
  SEN_ND4_8 U843 ( .A1(net59775), .A2(n443), .A3(n389), .A4(n1056), .X(
        net59793) );
  SEN_OR4_4 U847 ( .A1(n564), .A2(n446), .A3(n438), .A4(n439), .X(net59486) );
  SEN_NR2_T_4 U848 ( .A1(net59237), .A2(net59503), .X(n446) );
  SEN_AOAI211_1 U853 ( .A1(n561), .A2(net59216), .B(n562), .C(n563), .X(n360)
         );
  SEN_INV_5 U854 ( .A(n564), .X(n567) );
  SEN_OAI21B_8 U855 ( .A1(n555), .A2(n556), .B(n557), .X(n560) );
  SEN_INV_4 U860 ( .A(net59223), .X(net59219) );
  SEN_ND2_T_4 U867 ( .A1(net59413), .A2(n801), .X(net59223) );
  SEN_OAI21_S_4 U870 ( .A1(net59413), .A2(net59473), .B(net59474), .X(n568) );
  SEN_INV_3 U872 ( .A(net59461), .X(net59413) );
  SEN_MUXI2_S_1 U874 ( .D0(net58904), .D1(n385), .S(INST[3]), .X(Z[28]) );
  SEN_INV_2 U878 ( .A(net59427), .X(net59426) );
  SEN_MUXI2_S_1 U879 ( .D0(net58902), .D1(n371), .S(INST[3]), .X(Z[29]) );
  SEN_ND3_T_2 U886 ( .A1(net59962), .A2(net59794), .A3(net59322), .X(n594) );
  SEN_INV_10 U888 ( .A(net59444), .X(net59980) );
  SEN_INV_S_3 U894 ( .A(net59792), .X(net59775) );
  SEN_NR2_T_8 U895 ( .A1(n397), .A2(n398), .X(net61326) );
  SEN_ND2_T_2 U901 ( .A1(n599), .A2(net59671), .X(n808) );
  SEN_AOI211_6 U903 ( .A1(net59416), .A2(net59422), .B1(n362), .B2(n360), .X(
        net59421) );
  SEN_OAI21_S_0P5 U905 ( .A1(n451), .A2(net59405), .B(net59406), .X(n803) );
  SEN_OAI21B_6 U908 ( .A1(net59411), .A2(net59410), .B(n373), .X(n563) );
  SEN_AOI21B_0P5 U909 ( .A1(net59249), .A2(net59247), .B(net59248), .X(n447)
         );
  SEN_INV_0P65 U910 ( .A(net58929), .X(n536) );
  SEN_MUXI2_S_1 U914 ( .D0(net58929), .D1(n367), .S(INST[3]), .X(Z[18]) );
  SEN_EO2_G_2 U916 ( .A1(net59376), .A2(net59377), .X(net58929) );
  SEN_ND3_S_1 U917 ( .A1(n534), .A2(net58923), .A3(net58919), .X(n533) );
  SEN_ND2_4 U925 ( .A1(n565), .A2(net59233), .X(n459) );
  SEN_ND2_6 U939 ( .A1(n567), .A2(n450), .X(n565) );
  SEN_INV_AS_10 U941 ( .A(n1070), .X(net59247) );
  SEN_ND3_T_2 U942 ( .A1(net59490), .A2(n1071), .A3(n1072), .X(n1073) );
  SEN_ND3_S_8 U945 ( .A1(n399), .A2(n400), .A3(n675), .X(n687) );
  SEN_ND2_8 U949 ( .A1(n358), .A2(net59459), .X(n555) );
  SEN_AOAI211_4 U950 ( .A1(n1069), .A2(net59550), .B(net59247), .C(n489), .X(
        n486) );
  SEN_AOI21B_3 U952 ( .A1(net59533), .A2(net59239), .B(net59498), .X(net59535)
         );
  SEN_INV_S_6 U958 ( .A(n1075), .X(n358) );
  SEN_OAI21_S_0P5 U969 ( .A1(net60418), .A2(net59385), .B(net59386), .X(n805)
         );
  SEN_OAI21_5 U993 ( .A1(net59247), .A2(net59249), .B(net59402), .X(net59405)
         );
  SEN_AOI21B_3 U994 ( .A1(net59247), .A2(net59249), .B(net59248), .X(n451) );
  SEN_ND2B_S_0P5 U995 ( .A(n1057), .B(net59549), .X(net59395) );
  SEN_MUXI2_DG_12 U996 ( .D0(n575), .D1(n716), .S(B[3]), .X(n643) );
  SEN_EN2_S_8 U1000 ( .A1(A[1]), .A2(n468), .X(n463) );
  SEN_ND2_4 U1001 ( .A1(n592), .A2(n593), .X(net59792) );
  SEN_BUF_S_3 U1022 ( .A(n484), .X(n519) );
  SEN_INV_4 U1032 ( .A(n565), .X(net59231) );
  SEN_INV_4 U1047 ( .A(net59549), .X(net59249) );
  SEN_EO2_3 U1053 ( .A1(n530), .A2(net59211), .X(n1064) );
  SEN_INV_4 U1054 ( .A(n1064), .X(n529) );
  SEN_INV_S_4 U1055 ( .A(n669), .X(n670) );
  SEN_NR2_G_4 U1060 ( .A1(net59314), .A2(n407), .X(n480) );
  SEN_AN4_S_4 U1068 ( .A1(net58908), .A2(n531), .A3(net58917), .A4(net58915), 
        .X(n359) );
  SEN_NR2_S_2 U1069 ( .A1(n532), .A2(n533), .X(n531) );
  SEN_INV_1 U1089 ( .A(net58921), .X(n532) );
  SEN_OAI21_S_4 U1095 ( .A1(net59494), .A2(n780), .B(n355), .X(n800) );
  SEN_AN5_6 U1102 ( .A1(n1065), .A2(n1066), .A3(B[5]), .A4(INST[2]), .A5(
        INST[1]), .X(n1067) );
  SEN_INV_4 U1104 ( .A(INST[3]), .X(n1065) );
  SEN_INV_10 U1105 ( .A(N72), .X(n1066) );
  SEN_INV_S_3 U1106 ( .A(n1067), .X(net59754) );
  SEN_ND2B_V1_2 U1123 ( .A(A[0]), .B(net59873), .X(n593) );
  SEN_ND3_T_2 U1124 ( .A1(net58927), .A2(net58931), .A3(n538), .X(n537) );
  SEN_INV_S_0P5 U1127 ( .A(net59233), .X(n1068) );
  SEN_INV_0P5 U1134 ( .A(net59549), .X(n1069) );
  SEN_ND4_S_6 U1147 ( .A1(n1055), .A2(net59326), .A3(net59327), .A4(n389), .X(
        n461) );
  SEN_AOAI211_8 U1193 ( .A1(n495), .A2(n496), .B(n497), .C(n498), .X(n1070) );
  SEN_INV_S_2 U1194 ( .A(n507), .X(n496) );
  SEN_INV_4 U1219 ( .A(n446), .X(n450) );
  SEN_INV_S_0P5 U1222 ( .A(net59488), .X(n1071) );
  SEN_INV_S_0P5 U1335 ( .A(n782), .X(n1072) );
  SEN_INV_2 U1349 ( .A(n1073), .X(n783) );
  SEN_INV_S_3 U1378 ( .A(net59233), .X(net59498) );
  SEN_ND2B_V1_4 U1383 ( .A(n1074), .B(n797), .X(n1075) );
  SEN_INV_S_0P5 U1420 ( .A(net59438), .X(n1074) );
  SEN_ND3_T_16 U1449 ( .A1(n458), .A2(n469), .A3(INST[1]), .X(n465) );
  SEN_ND2_T_8 U1523 ( .A1(n388), .A2(n484), .X(n485) );
  SEN_ND3_1 U1533 ( .A1(n1076), .A2(net59370), .A3(net60495), .X(net59626) );
  SEN_ND2_T_5 U1534 ( .A1(net59744), .A2(net59743), .X(net59689) );
  SEN_INV_5 U1535 ( .A(net59776), .X(net59744) );
  SEN_AOAI211_1 U1536 ( .A1(n1078), .A2(net59274), .B(net59273), .C(net59276), 
        .X(net59272) );
  SEN_INV_S_0P5 U1537 ( .A(net59277), .X(n1078) );
  SEN_INV_S_2 U1538 ( .A(net59278), .X(net59273) );
  SEN_AOI21_S_8 U1539 ( .A1(n431), .A2(net59437), .B(n528), .X(n527) );
  SEN_INV_2 U1540 ( .A(net58914), .X(net59216) );
  SEN_AOI21B_8 U1541 ( .A1(net59237), .A2(n1079), .B(n570), .X(n564) );
  SEN_INV_S_0P5 U1542 ( .A(net59239), .X(n1079) );
  SEN_INV_8 U1543 ( .A(net59533), .X(net59237) );
  SEN_INV_S_0P5 U1544 ( .A(net59238), .X(n570) );
  SEN_OAI21_S_4 U1545 ( .A1(net59678), .A2(net59679), .B(net59680), .X(
        net59370) );
  SEN_INV_2 U1546 ( .A(net59345), .X(net59680) );
endmodule

