module ShiftLR (
	Z, 
	X, 
	S, 
	LEFT, 
	LOG);
   output [31:0] Z;
   input [31:0] X;
   input [4:0] S;
   input LEFT;
   input LOG;

   // Internal wires
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n10;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n89;
   wire n90;
   wire n92;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;

   SEN_OAI222_1 U289 (.X(n131), 
	.C2(n123), 
	.C1(n36), 
	.B2(n281), 
	.B1(n150), 
	.A2(n261), 
	.A1(n38));
   SEN_EO2_DG_4 U290 (.X(n123), 
	.A2(n256), 
	.A1(S[2]));
   SEN_NR2B_V1DG_2 U291 (.X(n256), 
	.B(n294), 
	.A(n342));
   SEN_BUF_S_1 U292 (.X(n281), 
	.A(n104));
   SEN_INV_2 U293 (.X(n78), 
	.A(n137));
   SEN_BUF_S_1 U294 (.X(n275), 
	.A(n99));
   SEN_ND2_0P5 U295 (.X(n333), 
	.A2(n167), 
	.A1(n349));
   SEN_NR3_G_1 U296 (.X(n190), 
	.A3(n152), 
	.A2(n269), 
	.A1(n268));
   SEN_BUF_S_1 U297 (.X(n280), 
	.A(n104));
   SEN_INV_S_1 U298 (.X(n23), 
	.A(n207));
   SEN_OAI211_1 U299 (.X(n151), 
	.B2(n172), 
	.B1(n39), 
	.A2(n158), 
	.A1(n66));
   SEN_AOI22_1 U300 (.X(n172), 
	.B2(n37), 
	.B1(n173), 
	.A2(n344), 
	.A1(n160));
   SEN_AO222_1 U301 (.X(n321), 
	.C2(n84), 
	.C1(n200), 
	.B2(n83), 
	.B1(n50), 
	.A2(n81), 
	.A1(n115));
   SEN_AOI221_1 U302 (.X(n213), 
	.C(n226), 
	.B2(n81), 
	.B1(n170), 
	.A2(n79), 
	.A1(n115));
   SEN_AOI221_1 U303 (.X(n209), 
	.C(n223), 
	.B2(n81), 
	.B1(n164), 
	.A2(n79), 
	.A1(n24));
   SEN_AOI221_1 U304 (.X(n201), 
	.C(n215), 
	.B2(n81), 
	.B1(n178), 
	.A2(n79), 
	.A1(n17));
   SEN_OR3_1 U305 (.X(n167), 
	.A3(n259), 
	.A2(n286), 
	.A1(n285));
   SEN_INV_S_1 U306 (.X(n34), 
	.A(n148));
   SEN_INV_S_1 U307 (.X(n81), 
	.A(n279));
   SEN_BUF_S_1 U308 (.X(n279), 
	.A(n104));
   SEN_INV_2 U309 (.X(n84), 
	.A(n123));
   SEN_INV_S_1 U310 (.X(n83), 
	.A(n108));
   SEN_AOI222_1 U311 (.X(n184), 
	.C2(n22), 
	.C1(n347), 
	.B2(n183), 
	.B1(n350), 
	.A2(n179), 
	.A1(n355));
   SEN_ND3_1 U312 (.X(Z[29]), 
	.A3(n149), 
	.A2(n267), 
	.A1(n266));
   SEN_AN3_1 U313 (.X(n149), 
	.A3(n320), 
	.A2(n319), 
	.A1(n318));
   SEN_OAI221_1 U314 (.X(n94), 
	.C(n237), 
	.B2(n280), 
	.B1(n188), 
	.A2(n317), 
	.A1(n116));
   SEN_AN2_S_1 U315 (.X(n257), 
	.A2(n258), 
	.A1(n79));
   SEN_INV_S_0P5 U316 (.X(n352), 
	.A(n257));
   SEN_INV_S_0P5 U317 (.X(n351), 
	.A(n257));
   SEN_AN3_0P5 U318 (.X(n258), 
	.A3(n86), 
	.A2(n212), 
	.A1(n130));
   SEN_OAI221_1 U319 (.X(n195), 
	.C(n211), 
	.B2(n280), 
	.B1(n190), 
	.A2(n317), 
	.A1(n113));
   SEN_INV_2 U320 (.X(n355), 
	.A(n238));
   SEN_INV_1 U321 (.X(n39), 
	.A(n152));
   SEN_INV_S_1 U322 (.X(n349), 
	.A(n338));
   SEN_AO22_1 U323 (.X(n259), 
	.B2(n133), 
	.B1(n81), 
	.A2(n28), 
	.A1(n79));
   SEN_INV_1 U324 (.X(n32), 
	.A(n216));
   SEN_INV_S_1 U325 (.X(n284), 
	.A(n195));
   SEN_ND2_G_1 U326 (.X(n137), 
	.A2(n342), 
	.A1(n212));
   SEN_AOI222_1 U327 (.X(n132), 
	.C2(n84), 
	.C1(n135), 
	.B2(n81), 
	.B1(n134), 
	.A2(n83), 
	.A1(n133));
   SEN_OA2BB2_0P5 U328 (.X(n129), 
	.B2(n132), 
	.B1(n130), 
	.A2(n131), 
	.A1(n130));
   SEN_AOI221_1 U329 (.X(n103), 
	.C(n32), 
	.B2(X[5]), 
	.B1(n337), 
	.A2(X[21]), 
	.A1(n345));
   SEN_INV_2 U330 (.X(n337), 
	.A(n331));
   SEN_OA2BB2_DG_1 U331 (.X(n235), 
	.B2(n103), 
	.B1(n106), 
	.A2(n24), 
	.A1(n83));
   SEN_AN2_DG_1 U332 (.X(n340), 
	.A2(n130), 
	.A1(n197));
   SEN_ND2_G_1 U333 (.X(n261), 
	.A2(n123), 
	.A1(n173));
   SEN_INV_S_1 U334 (.X(n260), 
	.A(n80));
   SEN_OAI22_S_0P5 U335 (.X(n215), 
	.B2(n175), 
	.B1(n106), 
	.A2(n193), 
	.A1(n261));
   SEN_AO2BB2_0P5 U336 (.X(n185), 
	.B2(n164), 
	.B1(n83), 
	.A2(n166), 
	.A1(n106));
   SEN_ND2_G_1 U337 (.X(n106), 
	.A2(n82), 
	.A1(n84));
   SEN_ND2_G_0P65 U338 (.X(n108), 
	.A2(n123), 
	.A1(n173));
   SEN_OAI211_0P5 U339 (.X(n135), 
	.B2(n159), 
	.B1(n39), 
	.A2(n158), 
	.A1(n64));
   SEN_ND2_T_0P5 U340 (.X(n158), 
	.A2(n82), 
	.A1(n78));
   SEN_AOI221_1 U341 (.X(n175), 
	.C(n32), 
	.B2(X[11]), 
	.B1(n337), 
	.A2(X[27]), 
	.A1(n346));
   SEN_ND2_G_1 U342 (.X(n262), 
	.A2(X[22]), 
	.A1(n345));
   SEN_ND2_G_1 U343 (.X(n263), 
	.A2(X[6]), 
	.A1(n336));
   SEN_AN3_1 U344 (.X(n203), 
	.A3(n297), 
	.A2(n263), 
	.A1(n262));
   SEN_INV_2 U345 (.X(n336), 
	.A(n331));
   SEN_AN2_S_1 U346 (.X(n264), 
	.A2(X[19]), 
	.A1(n346));
   SEN_AN2_S_0P5 U347 (.X(n265), 
	.A2(X[3]), 
	.A1(n337));
   SEN_NR3_0P8 U348 (.X(n120), 
	.A3(n32), 
	.A2(n265), 
	.A1(n264));
   SEN_INV_1 U349 (.X(n346), 
	.A(n341));
   SEN_OA22_DG_1 U350 (.X(n236), 
	.B2(n229), 
	.B1(n261), 
	.A2(n120), 
	.A1(n106));
   SEN_OR2_1 U351 (.X(n266), 
	.A2(n354), 
	.A1(n148));
   SEN_OR2_1 U352 (.X(n267), 
	.A2(n351), 
	.A1(n44));
   SEN_NR3_T_1 U353 (.X(n148), 
	.A3(n302), 
	.A2(n301), 
	.A1(n300));
   SEN_INV_S_1 U354 (.X(n354), 
	.A(n340));
   SEN_AN2_S_0P5 U355 (.X(n268), 
	.A2(n78), 
	.A1(X[0]));
   SEN_AN2_S_0P5 U356 (.X(n269), 
	.A2(X[16]), 
	.A1(n337));
   SEN_NR3_0P8 U357 (.X(n152), 
	.A3(n40), 
	.A2(n342), 
	.A1(LOG));
   SEN_AN2_S_0P5 U358 (.X(n270), 
	.A2(n117), 
	.A1(n316));
   SEN_AN2_S_0P5 U359 (.X(n271), 
	.A2(n321), 
	.A1(n349));
   SEN_AN2_S_1 U360 (.X(n272), 
	.A2(n110), 
	.A1(n347));
   SEN_NR3_T_2 U361 (.X(n124), 
	.A3(n272), 
	.A2(n271), 
	.A1(n270));
   SEN_OAI222_0P75 U362 (.X(n117), 
	.C2(n123), 
	.C1(n147), 
	.B2(n261), 
	.B1(n101), 
	.A2(n280), 
	.A1(n107));
   SEN_OAI222_1 U363 (.X(n110), 
	.C2(n123), 
	.C1(n127), 
	.B2(n261), 
	.B1(n126), 
	.A2(n280), 
	.A1(n125));
   SEN_OAI221_0P5 U364 (.X(Z[3]), 
	.C(n124), 
	.B2(n351), 
	.B1(n71), 
	.A2(n354), 
	.A1(n41));
   SEN_AN2_S_0P5 U365 (.X(n273), 
	.A2(X[13]), 
	.A1(n346));
   SEN_AN2_S_0P5 U366 (.X(n274), 
	.A2(X[29]), 
	.A1(n246));
   SEN_NR2_1 U367 (.X(n109), 
	.A2(n274), 
	.A1(n273));
   SEN_NR2_T_0P5 U368 (.X(n246), 
	.A2(n342), 
	.A1(n212));
   SEN_OA222_1 U369 (.X(n147), 
	.C2(n173), 
	.C1(n109), 
	.B2(n248), 
	.B1(n53), 
	.A2(n247), 
	.A1(n69));
   SEN_EO2_5 U370 (.X(n212), 
	.A2(S[4]), 
	.A1(n254));
   SEN_OAI21_4 U371 (.X(n254), 
	.B(n342), 
	.A2(n253), 
	.A1(S[3]));
   SEN_NR2_S_0P5 U372 (.X(n276), 
	.A2(n317), 
	.A1(n193));
   SEN_NR2_S_0P5 U373 (.X(n277), 
	.A2(n280), 
	.A1(n155));
   SEN_INV_S_1 U374 (.X(n278), 
	.A(n194));
   SEN_OR3_1 U375 (.X(n183), 
	.A3(n278), 
	.A2(n277), 
	.A1(n276));
   SEN_OA2BB2_0P5 U376 (.X(n194), 
	.B2(n175), 
	.B1(n261), 
	.A2(n178), 
	.A1(n80));
   SEN_OA22_1 U377 (.X(n230), 
	.B2(n193), 
	.B1(n106), 
	.A2(n120), 
	.A1(n261));
   SEN_ND2_S_0P5 U378 (.X(n104), 
	.A2(n82), 
	.A1(n123));
   SEN_OR2_DG_1 U379 (.X(n282), 
	.A2(n106), 
	.A1(n121));
   SEN_OR2_DG_1 U380 (.X(n283), 
	.A2(n84), 
	.A1(n122));
   SEN_ND3_1 U381 (.X(n146), 
	.A3(n249), 
	.A2(n283), 
	.A1(n282));
   SEN_NR2_S_0P5 U382 (.X(n285), 
	.A2(n261), 
	.A1(n181));
   SEN_NR2_S_0P5 U383 (.X(n286), 
	.A2(n260), 
	.A1(n161));
   SEN_AOI221_1 U384 (.X(n161), 
	.C(n152), 
	.B2(n74), 
	.B1(X[18]), 
	.A2(n78), 
	.A1(X[2]));
   SEN_OAI221_0P5 U385 (.X(n208), 
	.C(n218), 
	.B2(n281), 
	.B1(n181), 
	.A2(n317), 
	.A1(n125));
   SEN_OAI221_0P5 U386 (.X(n92), 
	.C(n239), 
	.B2(n280), 
	.B1(n203), 
	.A2(n317), 
	.A1(n126));
   SEN_OAI221_0P5 U387 (.X(n95), 
	.C(n105), 
	.B2(n280), 
	.B1(n103), 
	.A2(n317), 
	.A1(n101));
   SEN_OAI221_0P5 U388 (.X(n221), 
	.C(n230), 
	.B2(n280), 
	.B1(n175), 
	.A2(n317), 
	.A1(n229));
   SEN_OAI221_0P5 U389 (.X(n97), 
	.C(n114), 
	.B2(n280), 
	.B1(n113), 
	.A2(n317), 
	.A1(n112));
   SEN_OAI222_0P5 U390 (.X(n99), 
	.C2(n123), 
	.C1(n122), 
	.B2(n261), 
	.B1(n121), 
	.A2(n281), 
	.A1(n120));
   SEN_OAI221_1 U391 (.X(n227), 
	.C(n235), 
	.B2(n280), 
	.B1(n207), 
	.A2(n317), 
	.A1(n109));
   SEN_NR2_S_0P5 U392 (.X(n287), 
	.A2(n40), 
	.A1(n73));
   SEN_NR2_S_0P5 U393 (.X(n288), 
	.A2(n59), 
	.A1(n136));
   SEN_OR3_2 U394 (.X(n178), 
	.A3(n32), 
	.A2(n288), 
	.A1(n287));
   SEN_INV_S_2 U395 (.X(n73), 
	.A(n345));
   SEN_INV_1 U396 (.X(n40), 
	.A(X[31]));
   SEN_ND2_G_1 U397 (.X(n136), 
	.A2(n342), 
	.A1(n75));
   SEN_ND2_G_1 U398 (.X(n216), 
	.A2(n75), 
	.A1(n152));
   SEN_AOI22_0P75 U399 (.X(n177), 
	.B2(n178), 
	.B1(n173), 
	.A2(X[23]), 
	.A1(n160));
   SEN_ND2_G_1 U400 (.X(n289), 
	.A2(X[18]), 
	.A1(n346));
   SEN_ND2_S_0P5 U401 (.X(n290), 
	.A2(X[2]), 
	.A1(n336));
   SEN_INV_S_0P5 U402 (.X(n291), 
	.A(n32));
   SEN_AN3_1 U403 (.X(n125), 
	.A3(n291), 
	.A2(n290), 
	.A1(n289));
   SEN_OA22_DG_1 U404 (.X(n233), 
	.B2(n125), 
	.B1(n261), 
	.A2(n203), 
	.A1(n106));
   SEN_ND2_S_0P5 U405 (.X(n292), 
	.A2(X[25]), 
	.A1(n346));
   SEN_ND2_S_0P5 U406 (.X(n293), 
	.A2(X[9]), 
	.A1(n337));
   SEN_AN3_1 U407 (.X(n207), 
	.A3(n291), 
	.A2(n293), 
	.A1(n292));
   SEN_OAI22_0P5 U408 (.X(n223), 
	.B2(n207), 
	.B1(n106), 
	.A2(n103), 
	.A1(n261));
   SEN_BUF_2 U409 (.X(n316), 
	.A(n355));
   SEN_ND2_0P5 U410 (.X(n102), 
	.A2(n173), 
	.A1(n84));
   SEN_ND2_0P5 U411 (.X(n317), 
	.A2(n173), 
	.A1(n84));
   SEN_NR2_S_0P5 U412 (.X(n294), 
	.A2(S[0]), 
	.A1(S[1]));
   SEN_ND2_S_0P5 U413 (.X(n295), 
	.A2(X[20]), 
	.A1(n345));
   SEN_ND2_S_0P5 U414 (.X(n296), 
	.A2(X[4]), 
	.A1(n336));
   SEN_INV_S_0P5 U415 (.X(n297), 
	.A(n32));
   SEN_AN3_1 U416 (.X(n113), 
	.A3(n297), 
	.A2(n296), 
	.A1(n295));
   SEN_OAI22_S_0P5 U417 (.X(n226), 
	.B2(n188), 
	.B1(n106), 
	.A2(n113), 
	.A1(n261));
   SEN_OA2BB2_DG_1 U418 (.X(n237), 
	.B2(n113), 
	.B1(n106), 
	.A2(n115), 
	.A1(n83));
   SEN_NR2_G_0P5 U419 (.X(n326), 
	.A2(n317), 
	.A1(n175));
   SEN_OA2BB2_0P5 U420 (.X(n165), 
	.B2(n166), 
	.B1(n82), 
	.A2(X[25]), 
	.A1(n160));
   SEN_ND2_2 U421 (.X(n173), 
	.A2(n325), 
	.A1(n324));
   SEN_ND2_0P65 U422 (.X(n309), 
	.A2(n33), 
	.A1(n349));
   SEN_ND2_G_1 U423 (.X(n334), 
	.A2(n33), 
	.A1(n348));
   SEN_OAI221_1 U424 (.X(Z[25]), 
	.C(n169), 
	.B2(n351), 
	.B1(n48), 
	.A2(n354), 
	.A1(n168));
   SEN_ND2_S_0P5 U425 (.X(n303), 
	.A2(n78), 
	.A1(X[1]));
   SEN_ND2_S_0P5 U426 (.X(n304), 
	.A2(X[17]), 
	.A1(n74));
   SEN_AN3_1 U427 (.X(n166), 
	.A3(n39), 
	.A2(n304), 
	.A1(n303));
   SEN_NR2_T_2 U428 (.X(n255), 
	.A2(S[0]), 
	.A1(S[1]));
   SEN_INV_1 U429 (.X(n79), 
	.A(n102));
   SEN_INV_2 U430 (.X(n74), 
	.A(n136));
   SEN_AN3_S_1 U431 (.X(n153), 
	.A3(n307), 
	.A2(n306), 
	.A1(n305));
   SEN_INV_4 U432 (.X(n75), 
	.A(n212));
   SEN_INV_S_0P5 U433 (.X(n322), 
	.A(n252));
   SEN_AN3_1 U434 (.X(n157), 
	.A3(n310), 
	.A2(n309), 
	.A1(n308));
   SEN_AN3_1 U435 (.X(n169), 
	.A3(n334), 
	.A2(n333), 
	.A1(n332));
   SEN_ND2_S_0P5 U436 (.X(n298), 
	.A2(n344), 
	.A1(n346));
   SEN_ND2_S_0P5 U437 (.X(n299), 
	.A2(X[8]), 
	.A1(n336));
   SEN_AN3_1 U438 (.X(n188), 
	.A3(n291), 
	.A2(n299), 
	.A1(n298));
   SEN_OA2BB2_0P5 U439 (.X(n211), 
	.B2(n188), 
	.B1(n108), 
	.A2(n170), 
	.A1(n80));
   SEN_AN2_S_0P5 U440 (.X(n300), 
	.A2(n79), 
	.A1(n164));
   SEN_AN2_S_1 U441 (.X(n301), 
	.A2(n80), 
	.A1(n144));
   SEN_AN2_DG_1 U442 (.X(n302), 
	.A2(n123), 
	.A1(n142));
   SEN_OAI221_0P5 U443 (.X(n144), 
	.C(n39), 
	.B2(n53), 
	.B1(n331), 
	.A2(n137), 
	.A1(n69));
   SEN_INV_1 U444 (.X(n80), 
	.A(n106));
   SEN_INV_2 U445 (.X(n345), 
	.A(n341));
   SEN_INV_1 U446 (.X(n33), 
	.A(n153));
   SEN_OAI221_1 U447 (.X(Z[28]), 
	.C(n154), 
	.B2(n351), 
	.B1(n45), 
	.A2(n354), 
	.A1(n153));
   SEN_ND2_S_0P5 U448 (.X(n307), 
	.A2(n123), 
	.A1(n151));
   SEN_AOI221_0P5 U449 (.X(n155), 
	.C(n152), 
	.B2(X[19]), 
	.B1(n337), 
	.A2(n78), 
	.A1(X[3]));
   SEN_ND2_S_0P5 U450 (.X(n305), 
	.A2(n79), 
	.A1(n170));
   SEN_ND2_S_0P5 U451 (.X(n306), 
	.A2(n80), 
	.A1(n171));
   SEN_OAI221_0P5 U452 (.X(n170), 
	.C(n216), 
	.B2(n62), 
	.B1(n331), 
	.A2(n45), 
	.A1(n73));
   SEN_NR2B_V1DG_1 U453 (.X(n244), 
	.B(n102), 
	.A(n246));
   SEN_INV_S_1 U454 (.X(n347), 
	.A(n339));
   SEN_INV_S_0P5 U455 (.X(n323), 
	.A(S[3]));
   SEN_ND2B_V1_3 U456 (.X(n253), 
	.B(n255), 
	.A(S[2]));
   SEN_ND2_S_0P5 U457 (.X(n308), 
	.A2(n34), 
	.A1(n316));
   SEN_ND2_S_0P5 U458 (.X(n310), 
	.A2(n335), 
	.A1(n347));
   SEN_ND2_S_0P5 U459 (.X(n311), 
	.A2(n208), 
	.A1(n355));
   SEN_ND2_S_0P5 U460 (.X(n312), 
	.A2(n20), 
	.A1(n350));
   SEN_ND2_S_0P5 U461 (.X(n313), 
	.A2(n15), 
	.A1(n347));
   SEN_AN3_S_1 U462 (.X(n214), 
	.A3(n313), 
	.A2(n312), 
	.A1(n311));
   SEN_ND2_S_0P5 U463 (.X(n314), 
	.A2(X[23]), 
	.A1(n345));
   SEN_ND2_S_0P5 U464 (.X(n315), 
	.A2(X[7]), 
	.A1(n336));
   SEN_AN3_1 U465 (.X(n193), 
	.A3(n297), 
	.A2(n315), 
	.A1(n314));
   SEN_OAI221_1 U466 (.X(n90), 
	.C(n236), 
	.B2(n280), 
	.B1(n193), 
	.A2(n317), 
	.A1(n121));
   SEN_OA2BB2_DG_1 U467 (.X(n128), 
	.B2(n130), 
	.B1(n141), 
	.A2(n130), 
	.A1(n140));
   SEN_NR2_S_0P5 U468 (.X(n328), 
	.A2(n84), 
	.A1(n35));
   SEN_ND2_S_0P5 U469 (.X(n324), 
	.A2(n323), 
	.A1(n252));
   SEN_AOI222_1 U470 (.X(n174), 
	.C2(n162), 
	.C1(n347), 
	.B2(n22), 
	.B1(n350), 
	.A2(n167), 
	.A1(n355));
   SEN_ND3_S_1 U471 (.X(n186), 
	.A3(n204), 
	.A2(n330), 
	.A1(n329));
   SEN_ND2_S_0P5 U472 (.X(n248), 
	.A2(n173), 
	.A1(n246));
   SEN_ND2_S_0P5 U473 (.X(n247), 
	.A2(n173), 
	.A1(n345));
   SEN_OAI222_0P5 U474 (.X(n200), 
	.C2(n173), 
	.C1(n116), 
	.B2(n248), 
	.B1(n54), 
	.A2(n247), 
	.A1(n70));
   SEN_ND2_S_0P5 U475 (.X(n318), 
	.A2(n140), 
	.A1(n355));
   SEN_ND2_G_1 U476 (.X(n320), 
	.A2(n131), 
	.A1(n348));
   SEN_OA222_0P5 U477 (.X(n122), 
	.C2(n173), 
	.C1(n229), 
	.B2(n248), 
	.B1(n51), 
	.A2(n247), 
	.A1(n67));
   SEN_INV_S_0P5 U478 (.X(n82), 
	.A(n173));
   SEN_AOI221_0P5 U479 (.X(n181), 
	.C(n32), 
	.B2(n337), 
	.B1(X[14]), 
	.A2(n346), 
	.A1(X[30]));
   SEN_ND2_S_0P5 U480 (.X(n332), 
	.A2(n162), 
	.A1(n316));
   SEN_ND2_S_0P5 U481 (.X(n319), 
	.A2(n335), 
	.A1(n349));
   SEN_ND2_2 U482 (.X(n325), 
	.A2(S[3]), 
	.A1(n322));
   SEN_OA222_0P5 U483 (.X(n127), 
	.C2(n173), 
	.C1(n232), 
	.B2(n248), 
	.B1(n52), 
	.A2(n247), 
	.A1(n68));
   SEN_INV_S_1 U484 (.X(n353), 
	.A(n340));
   SEN_OA22_DG_1 U485 (.X(n105), 
	.B2(n109), 
	.B1(n108), 
	.A2(n107), 
	.A1(n106));
   SEN_OA22_DG_1 U486 (.X(n239), 
	.B2(n232), 
	.B1(n108), 
	.A2(n125), 
	.A1(n106));
   SEN_AOI22_0P5 U487 (.X(n189), 
	.B2(n37), 
	.B1(n80), 
	.A2(n170), 
	.A1(n83));
   SEN_AOI222_0P5 U488 (.X(n118), 
	.C2(n84), 
	.C1(n200), 
	.B2(n83), 
	.B1(n50), 
	.A2(n81), 
	.A1(n115));
   SEN_NR2_G_1 U489 (.X(n197), 
	.A2(n343), 
	.A1(n257));
   SEN_AOI222_1 U490 (.X(n111), 
	.C2(n97), 
	.C1(n348), 
	.B2(n110), 
	.B1(n349), 
	.A2(n275), 
	.A1(n316));
   SEN_AOI22_0P5 U491 (.X(n204), 
	.B2(n31), 
	.B1(n80), 
	.A2(n28), 
	.A1(n83));
   SEN_OR3_1 U492 (.X(n162), 
	.A3(n328), 
	.A2(n327), 
	.A1(n326));
   SEN_OAI22_S_0P5 U493 (.X(n245), 
	.B2(n106), 
	.B1(n101), 
	.A2(n84), 
	.A1(n147));
   SEN_AOI221_0P5 U494 (.X(n219), 
	.C(n32), 
	.B2(X[10]), 
	.B1(n336), 
	.A2(X[26]), 
	.A1(n346));
   SEN_AOI22_0P5 U495 (.X(n241), 
	.B2(X[0]), 
	.B1(n257), 
	.A2(n196), 
	.A1(n343));
   SEN_OAI221_0P5 U496 (.X(Z[0]), 
	.C(n241), 
	.B2(n238), 
	.B1(n43), 
	.A2(n353), 
	.A1(n240));
   SEN_INV_1 U497 (.X(n35), 
	.A(n176));
   SEN_EO2_S_0P5 U498 (.X(n130), 
	.A2(S[1]), 
	.A1(n251));
   SEN_AO221_0P5 U499 (.X(Z[1]), 
	.C(n199), 
	.B2(n350), 
	.B1(n198), 
	.A2(n197), 
	.A1(n196));
   SEN_AO22_DG_1 U500 (.X(n199), 
	.B2(X[1]), 
	.B1(n257), 
	.A2(n321), 
	.A1(n348));
   SEN_NR2_S_0P5 U501 (.X(n327), 
	.A2(n106), 
	.A1(n155));
   SEN_INV_1 U502 (.X(n29), 
	.A(n162));
   SEN_AOI222_1 U503 (.X(n187), 
	.C2(n179), 
	.C1(n347), 
	.B2(n186), 
	.B1(n350), 
	.A2(n183), 
	.A1(n355));
   SEN_AOI22_0P5 U504 (.X(n206), 
	.B2(n164), 
	.B1(n80), 
	.A2(n23), 
	.A1(n83));
   SEN_INV_S_0P5 U505 (.X(n85), 
	.A(n130));
   SEN_INV_S_0P5 U506 (.X(n5), 
	.A(n186));
   SEN_AOI222_0P5 U507 (.X(n138), 
	.C2(n123), 
	.C1(n135), 
	.B2(n80), 
	.B1(n133), 
	.A2(n79), 
	.A1(n31));
   SEN_INV_S_0P5 U508 (.X(n17), 
	.A(n120));
   SEN_AOI222_0P5 U509 (.X(n141), 
	.C2(n144), 
	.C1(n83), 
	.B2(n143), 
	.B1(n81), 
	.A2(n142), 
	.A1(n84));
   SEN_OAI221_0P5 U510 (.X(n143), 
	.C(n39), 
	.B2(n44), 
	.B1(n331), 
	.A2(n137), 
	.A1(n61));
   SEN_INV_1 U511 (.X(n24), 
	.A(n107));
   SEN_INV_1 U512 (.X(n50), 
	.A(n112));
   SEN_OR2_DG_1 U513 (.X(n339), 
	.A2(n130), 
	.A1(n86));
   SEN_AO222_1 U514 (.X(n335), 
	.C2(n123), 
	.C1(n135), 
	.B2(n80), 
	.B1(n133), 
	.A2(n79), 
	.A1(n31));
   SEN_AOI22_0P5 U515 (.X(n229), 
	.B2(X[31]), 
	.B1(n246), 
	.A2(X[15]), 
	.A1(n346));
   SEN_OR2_DG_1 U516 (.X(n329), 
	.A2(n317), 
	.A1(n203));
   SEN_OR2_DG_1 U517 (.X(n330), 
	.A2(n281), 
	.A1(n161));
   SEN_INV_S_6 U518 (.X(n331), 
	.A(n74));
   SEN_NR2_S_0P5 U519 (.X(n243), 
	.A2(n73), 
	.A1(n102));
   SEN_INV_1 U520 (.X(n22), 
	.A(n168));
   SEN_INV_2 U521 (.X(n20), 
	.A(n209));
   SEN_INV_2 U522 (.X(n15), 
	.A(n201));
   SEN_INV_2 U523 (.X(n8), 
	.A(n213));
   SEN_NR2_S_0P5 U524 (.X(n160), 
	.A2(n173), 
	.A1(n331));
   SEN_OAI221_0P5 U525 (.X(n164), 
	.C(n216), 
	.B2(n61), 
	.B1(n331), 
	.A2(n44), 
	.A1(n73));
   SEN_OAI221_0P5 U526 (.X(n171), 
	.C(n39), 
	.B2(n54), 
	.B1(n331), 
	.A2(n137), 
	.A1(n70));
   SEN_AOI221_1 U527 (.X(n168), 
	.C(n185), 
	.B2(n81), 
	.B1(n144), 
	.A2(n79), 
	.A1(n23));
   SEN_INV_S_0P5 U528 (.X(n21), 
	.A(n191));
   SEN_INV_S_0P5 U529 (.X(n2), 
	.A(n92));
   SEN_INV_S_0P5 U530 (.X(n16), 
	.A(n183));
   SEN_INV_S_0P5 U531 (.X(n7), 
	.A(n94));
   SEN_INV_S_0P5 U532 (.X(n14), 
	.A(n221));
   SEN_INV_S_0P5 U533 (.X(n6), 
	.A(n110));
   SEN_INV_S_0P5 U534 (.X(n10), 
	.A(n179));
   SEN_INV_S_0P5 U535 (.X(n25), 
	.A(n117));
   SEN_INV_S_0P5 U536 (.X(n19), 
	.A(n227));
   SEN_INV_S_0P5 U537 (.X(n3), 
	.A(n224));
   SEN_INV_S_0P5 U538 (.X(n26), 
	.A(n95));
   SEN_INV_S_0P5 U539 (.X(n12), 
	.A(n97));
   SEN_INV_1 U540 (.X(n41), 
	.A(n146));
   SEN_INV_1 U541 (.X(n37), 
	.A(n190));
   SEN_OR2_DG_1 U542 (.X(n341), 
	.A2(n342), 
	.A1(n75));
   SEN_AOI221_0P5 U543 (.X(n150), 
	.C(n152), 
	.B2(X[12]), 
	.B1(n78), 
	.A2(n337), 
	.A1(X[28]));
   SEN_INV_S_0P5 U544 (.X(n36), 
	.A(n151));
   SEN_OAI222_0P5 U545 (.X(n140), 
	.C2(n123), 
	.C1(n35), 
	.B2(n281), 
	.B1(n156), 
	.A2(n261), 
	.A1(n155));
   SEN_AOI221_0P5 U546 (.X(n156), 
	.C(n152), 
	.B2(X[11]), 
	.B1(n78), 
	.A2(n336), 
	.A1(X[27]));
   SEN_ND2_S_0P5 U547 (.X(n251), 
	.A2(n342), 
	.A1(n343));
   SEN_INV_S_0P5 U548 (.X(n27), 
	.A(n167));
   SEN_AOI22_0P5 U549 (.X(n116), 
	.B2(X[28]), 
	.B1(n246), 
	.A2(X[12]), 
	.A1(n345));
   SEN_OAI221_0P5 U550 (.X(n198), 
	.C(n250), 
	.B2(n84), 
	.B1(n127), 
	.A2(n260), 
	.A1(n126));
   SEN_AOI22_0P5 U551 (.X(n232), 
	.B2(X[30]), 
	.B1(n246), 
	.A2(X[14]), 
	.A1(n345));
   SEN_AOI22_0P5 U552 (.X(n121), 
	.B2(X[27]), 
	.B1(n246), 
	.A2(X[11]), 
	.A1(n345));
   SEN_AOI22_0P5 U553 (.X(n126), 
	.B2(X[26]), 
	.B1(n246), 
	.A2(X[10]), 
	.A1(n346));
   SEN_AOI22_0P5 U554 (.X(n101), 
	.B2(X[25]), 
	.B1(n246), 
	.A2(X[9]), 
	.A1(n345));
   SEN_AOI22_0P5 U555 (.X(n112), 
	.B2(n344), 
	.B1(n246), 
	.A2(X[8]), 
	.A1(n346));
   SEN_AO221_0P5 U556 (.X(n115), 
	.C(n32), 
	.B2(X[0]), 
	.B1(n337), 
	.A2(X[16]), 
	.A1(n345));
   SEN_INV_S_0P5 U557 (.X(n4), 
	.A(n208));
   SEN_AOI222_0P5 U558 (.X(n240), 
	.C2(n50), 
	.C1(n80), 
	.B2(X[16]), 
	.B1(n244), 
	.A2(n200), 
	.A1(n123));
   SEN_BUF_6 U559 (.X(n342), 
	.A(LEFT));
   SEN_OAI211_1 U560 (.X(n142), 
	.B2(n165), 
	.B1(n39), 
	.A2(n158), 
	.A1(n65));
   SEN_BUF_1 U561 (.X(n343), 
	.A(S[0]));
   SEN_INV_1 U562 (.X(n31), 
	.A(n181));
   SEN_INV_S_1 U563 (.X(n350), 
	.A(n338));
   SEN_INV_S_1 U564 (.X(n38), 
	.A(n171));
   SEN_OR2_1 U565 (.X(n338), 
	.A2(n86), 
	.A1(n85));
   SEN_ND2_G_1 U566 (.X(n238), 
	.A2(n85), 
	.A1(n197));
   SEN_INV_S_1 U567 (.X(n348), 
	.A(n339));
   SEN_OAI221_1 U568 (.X(n179), 
	.C(n189), 
	.B2(n281), 
	.B1(n38), 
	.A2(n317), 
	.A1(n188));
   SEN_OA2BB2_1 U569 (.X(n218), 
	.B2(n203), 
	.B1(n261), 
	.A2(n28), 
	.A1(n80));
   SEN_OAI221_1 U570 (.X(n191), 
	.C(n206), 
	.B2(n281), 
	.B1(n166), 
	.A2(n317), 
	.A1(n103));
   SEN_OAI221_1 U571 (.X(n224), 
	.C(n233), 
	.B2(n280), 
	.B1(n219), 
	.A2(n317), 
	.A1(n232));
   SEN_OA2BB2_1 U572 (.X(n114), 
	.B2(n116), 
	.B1(n108), 
	.A2(n115), 
	.A1(n80));
   SEN_OAI221_1 U573 (.X(n133), 
	.C(n39), 
	.B2(n52), 
	.B1(n331), 
	.A2(n137), 
	.A1(n68));
   SEN_OAI222_1 U574 (.X(Z[31]), 
	.C2(n351), 
	.C1(n40), 
	.B2(n86), 
	.B1(n129), 
	.A2(n128), 
	.A1(n343));
   SEN_OAI221_0P5 U575 (.X(n134), 
	.C(n39), 
	.B2(n60), 
	.B1(n137), 
	.A2(n42), 
	.A1(n331));
   SEN_OAI221_1 U576 (.X(Z[4]), 
	.C(n119), 
	.B2(n351), 
	.B1(n70), 
	.A2(n354), 
	.A1(n118));
   SEN_AOI222_1 U577 (.X(n119), 
	.C2(n275), 
	.C1(n348), 
	.B2(n117), 
	.B1(n349), 
	.A2(n110), 
	.A1(n316));
   SEN_OAI221_1 U578 (.X(Z[30]), 
	.C(n139), 
	.B2(n351), 
	.B1(n42), 
	.A2(n354), 
	.A1(n138));
   SEN_OA2BB2_1 U579 (.X(n139), 
	.B2(n128), 
	.B1(n86), 
	.A2(n131), 
	.A1(n316));
   SEN_AOI222_1 U580 (.X(n154), 
	.C2(n140), 
	.C1(n348), 
	.B2(n34), 
	.B1(n349), 
	.A2(n335), 
	.A1(n316));
   SEN_OAI221_1 U581 (.X(Z[6]), 
	.C(n100), 
	.B2(n351), 
	.B1(n68), 
	.A2(n354), 
	.A1(n6));
   SEN_AOI222_1 U582 (.X(n100), 
	.C2(n95), 
	.C1(n348), 
	.B2(n275), 
	.B1(n349), 
	.A2(n97), 
	.A1(n316));
   SEN_OAI221_1 U583 (.X(Z[7]), 
	.C(n98), 
	.B2(n351), 
	.B1(n67), 
	.A2(n354), 
	.A1(n18));
   SEN_INV_S_1 U584 (.X(n18), 
	.A(n275));
   SEN_AOI222_1 U585 (.X(n98), 
	.C2(n92), 
	.C1(n348), 
	.B2(n97), 
	.B1(n349), 
	.A2(n95), 
	.A1(n316));
   SEN_OAI221_1 U586 (.X(Z[5]), 
	.C(n111), 
	.B2(n351), 
	.B1(n69), 
	.A2(n354), 
	.A1(n25));
   SEN_INV_1 U587 (.X(n28), 
	.A(n219));
   SEN_OAI221_1 U588 (.X(Z[24]), 
	.C(n174), 
	.B2(n352), 
	.B1(n49), 
	.A2(n354), 
	.A1(n10));
   SEN_INV_S_1 U589 (.X(n49), 
	.A(n344));
   SEN_OAI221_1 U590 (.X(Z[9]), 
	.C(n89), 
	.B2(n352), 
	.B1(n65), 
	.A2(n353), 
	.A1(n26));
   SEN_AOI222_1 U591 (.X(n89), 
	.C2(n94), 
	.C1(n347), 
	.B2(n92), 
	.B1(n350), 
	.A2(n90), 
	.A1(n355));
   SEN_OAI221_1 U592 (.X(Z[10]), 
	.C(n234), 
	.B2(n351), 
	.B1(n64), 
	.A2(n353), 
	.A1(n2));
   SEN_AOI222_1 U593 (.X(n234), 
	.C2(n227), 
	.C1(n348), 
	.B2(n90), 
	.B1(n349), 
	.A2(n94), 
	.A1(n316));
   SEN_OAI221_1 U594 (.X(Z[20]), 
	.C(n192), 
	.B2(n352), 
	.B1(n54), 
	.A2(n353), 
	.A1(n284));
   SEN_AOI222_1 U595 (.X(n192), 
	.C2(n183), 
	.C1(n347), 
	.B2(n191), 
	.B1(n350), 
	.A2(n186), 
	.A1(n355));
   SEN_OAI221_1 U596 (.X(Z[21]), 
	.C(n187), 
	.B2(n352), 
	.B1(n53), 
	.A2(n353), 
	.A1(n21));
   SEN_OAI221_1 U597 (.X(Z[23]), 
	.C(n180), 
	.B2(n352), 
	.B1(n51), 
	.A2(n354), 
	.A1(n16));
   SEN_AOI222_1 U598 (.X(n180), 
	.C2(n167), 
	.C1(n347), 
	.B2(n179), 
	.B1(n350), 
	.A2(n22), 
	.A1(n355));
   SEN_OAI221_1 U599 (.X(Z[12]), 
	.C(n228), 
	.B2(n352), 
	.B1(n62), 
	.A2(n353), 
	.A1(n7));
   SEN_AOI222_1 U600 (.X(n228), 
	.C2(n221), 
	.C1(n348), 
	.B2(n227), 
	.B1(n349), 
	.A2(n224), 
	.A1(n316));
   SEN_OAI221_1 U601 (.X(Z[13]), 
	.C(n225), 
	.B2(n352), 
	.B1(n61), 
	.A2(n353), 
	.A1(n19));
   SEN_AOI222_1 U602 (.X(n225), 
	.C2(n8), 
	.C1(n347), 
	.B2(n224), 
	.B1(n350), 
	.A2(n221), 
	.A1(n355));
   SEN_OAI221_1 U603 (.X(Z[14]), 
	.C(n222), 
	.B2(n352), 
	.B1(n60), 
	.A2(n353), 
	.A1(n3));
   SEN_AOI222_1 U604 (.X(n222), 
	.C2(n20), 
	.C1(n347), 
	.B2(n221), 
	.B1(n350), 
	.A2(n8), 
	.A1(n355));
   SEN_OAI221_1 U605 (.X(Z[15]), 
	.C(n217), 
	.B2(n352), 
	.B1(n59), 
	.A2(n353), 
	.A1(n14));
   SEN_AOI222_1 U606 (.X(n217), 
	.C2(n208), 
	.C1(n347), 
	.B2(n8), 
	.B1(n350), 
	.A2(n20), 
	.A1(n355));
   SEN_OAI221_1 U607 (.X(Z[22]), 
	.C(n184), 
	.B2(n352), 
	.B1(n52), 
	.A2(n353), 
	.A1(n5));
   SEN_OAI221_1 U608 (.X(Z[8]), 
	.C(n96), 
	.B2(n351), 
	.B1(n66), 
	.A2(n354), 
	.A1(n12));
   SEN_AOI222_1 U609 (.X(n96), 
	.C2(n90), 
	.C1(n348), 
	.B2(n95), 
	.B1(n349), 
	.A2(n92), 
	.A1(n316));
   SEN_INV_S_1 U610 (.X(n86), 
	.A(n343));
   SEN_INV_S_1 U611 (.X(n43), 
	.A(n198));
   SEN_AOI221_1 U612 (.X(n107), 
	.C(n32), 
	.B2(X[1]), 
	.B1(n336), 
	.A2(X[17]), 
	.A1(n345));
   SEN_AOI22_1 U613 (.X(n249), 
	.B2(X[19]), 
	.B1(n244), 
	.A2(X[3]), 
	.A1(n243));
   SEN_OA2BB2_1 U614 (.X(n159), 
	.B2(n161), 
	.B1(n82), 
	.A2(X[26]), 
	.A1(n160));
   SEN_AOI22_1 U615 (.X(n250), 
	.B2(X[18]), 
	.B1(n244), 
	.A2(X[2]), 
	.A1(n243));
   SEN_ND2_S_0P5 U616 (.X(n252), 
	.A2(n253), 
	.A1(n342));
   SEN_OAI221_1 U617 (.X(Z[16]), 
	.C(n214), 
	.B2(n352), 
	.B1(n58), 
	.A2(n353), 
	.A1(n213));
   SEN_INV_S_1 U618 (.X(n58), 
	.A(X[16]));
   SEN_OAI221_1 U619 (.X(Z[17]), 
	.C(n210), 
	.B2(n352), 
	.B1(n57), 
	.A2(n353), 
	.A1(n209));
   SEN_INV_S_1 U620 (.X(n57), 
	.A(X[17]));
   SEN_AOI222_1 U621 (.X(n210), 
	.C2(n195), 
	.C1(n347), 
	.B2(n208), 
	.B1(n350), 
	.A2(n15), 
	.A1(n355));
   SEN_OAI22_1 U622 (.X(n196), 
	.B2(n85), 
	.B1(n242), 
	.A2(n130), 
	.A1(n41));
   SEN_AOI221_1 U623 (.X(n242), 
	.C(n245), 
	.B2(X[17]), 
	.B1(n244), 
	.A2(X[1]), 
	.A1(n243));
   SEN_INV_S_1 U624 (.X(n48), 
	.A(X[25]));
   SEN_OAI221_1 U625 (.X(Z[19]), 
	.C(n202), 
	.B2(n352), 
	.B1(n55), 
	.A2(n353), 
	.A1(n201));
   SEN_INV_S_1 U626 (.X(n55), 
	.A(X[19]));
   SEN_AOI222_1 U627 (.X(n202), 
	.C2(n186), 
	.C1(n347), 
	.B2(n195), 
	.B1(n350), 
	.A2(n191), 
	.A1(n355));
   SEN_OAI221_1 U628 (.X(Z[27]), 
	.C(n157), 
	.B2(n351), 
	.B1(n46), 
	.A2(n354), 
	.A1(n29));
   SEN_INV_S_1 U629 (.X(n46), 
	.A(X[27]));
   SEN_INV_S_1 U630 (.X(n71), 
	.A(X[3]));
   SEN_OAI221_1 U631 (.X(Z[18]), 
	.C(n205), 
	.B2(n352), 
	.B1(n56), 
	.A2(n353), 
	.A1(n4));
   SEN_INV_S_1 U632 (.X(n56), 
	.A(X[18]));
   SEN_AOI222_1 U633 (.X(n205), 
	.C2(n191), 
	.C1(n347), 
	.B2(n15), 
	.B1(n350), 
	.A2(n195), 
	.A1(n355));
   SEN_OAI221_1 U634 (.X(Z[11]), 
	.C(n231), 
	.B2(n352), 
	.B1(n63), 
	.A2(n353), 
	.A1(n13));
   SEN_INV_S_1 U635 (.X(n63), 
	.A(X[11]));
   SEN_INV_S_1 U636 (.X(n13), 
	.A(n90));
   SEN_AOI222_1 U637 (.X(n231), 
	.C2(n224), 
	.C1(n348), 
	.B2(n94), 
	.B1(n349), 
	.A2(n227), 
	.A1(n316));
   SEN_OAI221_1 U638 (.X(Z[26]), 
	.C(n163), 
	.B2(n351), 
	.B1(n47), 
	.A2(n354), 
	.A1(n27));
   SEN_INV_S_1 U639 (.X(n47), 
	.A(X[26]));
   SEN_AOI222_1 U640 (.X(n163), 
	.C2(n34), 
	.C1(n348), 
	.B2(n162), 
	.B1(n349), 
	.A2(n33), 
	.A1(n316));
   SEN_OAI221_1 U641 (.X(Z[2]), 
	.C(n145), 
	.B2(n351), 
	.B1(n72), 
	.A2(n354), 
	.A1(n43));
   SEN_INV_S_1 U642 (.X(n72), 
	.A(X[2]));
   SEN_AOI222_1 U643 (.X(n145), 
	.C2(n117), 
	.C1(n348), 
	.B2(n146), 
	.B1(n349), 
	.A2(n321), 
	.A1(n316));
   SEN_INV_S_1 U644 (.X(n45), 
	.A(X[28]));
   SEN_INV_S_1 U645 (.X(n42), 
	.A(X[30]));
   SEN_INV_S_1 U646 (.X(n44), 
	.A(X[29]));
   SEN_INV_S_1 U647 (.X(n62), 
	.A(X[12]));
   SEN_INV_S_1 U648 (.X(n60), 
	.A(X[14]));
   SEN_INV_S_1 U649 (.X(n65), 
	.A(X[9]));
   SEN_INV_S_1 U650 (.X(n66), 
	.A(X[8]));
   SEN_INV_S_1 U651 (.X(n64), 
	.A(X[10]));
   SEN_INV_S_1 U652 (.X(n61), 
	.A(X[13]));
   SEN_INV_S_1 U653 (.X(n51), 
	.A(X[23]));
   SEN_INV_S_1 U654 (.X(n54), 
	.A(X[20]));
   SEN_INV_S_1 U655 (.X(n70), 
	.A(X[4]));
   SEN_INV_S_1 U656 (.X(n53), 
	.A(X[21]));
   SEN_INV_S_1 U657 (.X(n52), 
	.A(X[22]));
   SEN_INV_S_1 U658 (.X(n59), 
	.A(X[15]));
   SEN_INV_S_1 U659 (.X(n67), 
	.A(X[7]));
   SEN_INV_S_1 U660 (.X(n69), 
	.A(X[5]));
   SEN_INV_S_1 U661 (.X(n68), 
	.A(X[6]));
   SEN_OAI211_1 U662 (.X(n176), 
	.B2(n177), 
	.B1(n39), 
	.A2(n158), 
	.A1(n67));
   SEN_BUF_S_1 U663 (.X(n344), 
	.A(X[24]));
endmodule

