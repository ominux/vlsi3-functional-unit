
module Alu ( Z, A, B, INST, SEL );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  input SEL;
  wire   n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926;

  SEN_NR2_1 U345 ( .A1(n818), .A2(n817), .X(n576) );
  SEN_ND2_G_1 U346 ( .A1(n777), .A2(n776), .X(n502) );
  SEN_ND2_G_1 U347 ( .A1(n841), .A2(n840), .X(n556) );
  SEN_NR2_S_5 U348 ( .A1(n893), .A2(n754), .X(n653) );
  SEN_NR2_T_1 U349 ( .A1(n717), .A2(n716), .X(n508) );
  SEN_AOI21_T_1 U350 ( .A1(n585), .A2(n584), .B(n583), .X(n586) );
  SEN_INV_S_1 U351 ( .A(n579), .X(n584) );
  SEN_NR2_S_5 U352 ( .A1(n577), .A2(n327), .X(n666) );
  SEN_INV_S_1 U353 ( .A(n342), .X(n456) );
  SEN_ND2_G_1 U354 ( .A1(n717), .A2(n716), .X(n526) );
  SEN_INV_S_1 U355 ( .A(n501), .X(n340) );
  SEN_NR2_1 U356 ( .A1(n559), .A2(n558), .X(n580) );
  SEN_NR2_2 U357 ( .A1(n426), .A2(n872), .X(n623) );
  SEN_INV_S_1 U358 ( .A(n666), .X(n668) );
  SEN_NR2_1 U359 ( .A1(n701), .A2(n336), .X(n382) );
  SEN_INV_2 U360 ( .A(n708), .X(n522) );
  SEN_NR2_T_1 U361 ( .A1(n732), .A2(n731), .X(n536) );
  SEN_ND3_1 U362 ( .A1(n562), .A2(n545), .A3(n544), .X(n547) );
  SEN_OAI21_G_1 U363 ( .A1(n419), .A2(n557), .B(n579), .X(n614) );
  SEN_INV_S_1 U364 ( .A(n432), .X(n615) );
  SEN_AOI21B_2 U365 ( .A1(n350), .A2(n854), .B(n326), .X(n351) );
  SEN_AN2_DG_4 U366 ( .A1(n674), .A2(n593), .X(n630) );
  SEN_INV_S_1 U367 ( .A(n459), .X(n686) );
  SEN_EO2_S_0P5 U368 ( .A1(n725), .A2(n726), .X(n723) );
  SEN_BUF_S_1 U369 ( .A(n726), .X(n335) );
  SEN_EO2_S_0P5 U370 ( .A1(n731), .A2(n732), .X(n734) );
  SEN_MUXI2_S_2 U371 ( .D0(n438), .D1(n435), .S(A[5]), .X(n740) );
  SEN_EN2_0P5 U372 ( .A1(n747), .A2(n420), .X(n752) );
  SEN_BUF_S_1 U373 ( .A(n748), .X(n420) );
  SEN_EO2_S_0P5 U374 ( .A1(n763), .A2(n764), .X(n761) );
  SEN_MUXI2_DG_5 U375 ( .D0(n441), .D1(n442), .S(n339), .X(n771) );
  SEN_INV_S_1 U376 ( .A(B[9]), .X(n339) );
  SEN_EO2_S_0P5 U377 ( .A1(n776), .A2(n777), .X(n779) );
  SEN_EO2_S_0P5 U378 ( .A1(n783), .A2(n784), .X(n786) );
  SEN_EO2_S_0P5 U379 ( .A1(n790), .A2(n346), .X(n792) );
  SEN_EO2_S_0P5 U380 ( .A1(n796), .A2(n797), .X(n799) );
  SEN_INV_S_1 U381 ( .A(n544), .X(n806) );
  SEN_INV_S_1 U382 ( .A(n533), .X(n811) );
  SEN_EO2_S_0P5 U383 ( .A1(n810), .A2(n811), .X(n813) );
  SEN_MUXI2_S_2 U384 ( .D0(n439), .D1(n436), .S(A[17]), .X(n825) );
  SEN_MUXI2_S_2 U385 ( .D0(n443), .D1(n344), .S(B[17]), .X(n826) );
  SEN_EO2_S_0P5 U386 ( .A1(n825), .A2(n826), .X(n828) );
  SEN_MUXI2_S_2 U387 ( .D0(n439), .D1(n436), .S(A[19]), .X(n840) );
  SEN_MUXI2_S_2 U388 ( .D0(n439), .D1(n436), .S(A[20]), .X(n847) );
  SEN_EO2_S_0P5 U389 ( .A1(n847), .A2(n848), .X(n850) );
  SEN_EO2_S_0P5 U390 ( .A1(n854), .A2(n855), .X(n857) );
  SEN_MUXI2_S_2 U391 ( .D0(n439), .D1(n436), .S(A[21]), .X(n854) );
  SEN_EO2_1 U392 ( .A1(n857), .A2(n350), .X(n860) );
  SEN_INV_S_1 U393 ( .A(n900), .X(n445) );
  SEN_ND2_G_1 U394 ( .A1(n414), .A2(n416), .X(n862) );
  SEN_ND2_G_1 U395 ( .A1(n439), .A2(n415), .X(n416) );
  SEN_ND2_G_1 U396 ( .A1(n436), .A2(A[22]), .X(n414) );
  SEN_EO2_S_0P5 U397 ( .A1(n660), .A2(n659), .X(n861) );
  SEN_EO2_S_0P5 U398 ( .A1(n872), .A2(n426), .X(n874) );
  SEN_MUXI2_S_1 U399 ( .D0(n345), .D1(n444), .S(n879), .X(n877) );
  SEN_MUXI2_S_1 U400 ( .D0(n345), .D1(n444), .S(n889), .X(n886) );
  SEN_EO2_S_0P5 U401 ( .A1(n640), .A2(n639), .X(n891) );
  SEN_EO2_S_0P5 U402 ( .A1(n894), .A2(n895), .X(n896) );
  SEN_INV_S_1 U403 ( .A(n926), .X(n333) );
  SEN_INV_S_1 U404 ( .A(n917), .X(n897) );
  SEN_NR2_1 U405 ( .A1(n418), .A2(n693), .X(n900) );
  SEN_INV_S_1 U406 ( .A(n926), .X(n906) );
  SEN_INV_S_1 U407 ( .A(n704), .X(n910) );
  SEN_EN2_0P5 U408 ( .A1(n920), .A2(n921), .X(n925) );
  SEN_INV_S_1 U409 ( .A(n900), .X(n919) );
  SEN_INV_S_1 U410 ( .A(n428), .X(n447) );
  SEN_NR2_1 U411 ( .A1(n865), .A2(n866), .X(n329) );
  SEN_AOI22_0P5 U412 ( .A1(n353), .A2(n917), .B1(n906), .B2(n861), .X(n312) );
  SEN_OAI21_0P5 U413 ( .A1(A[22]), .A2(B[22]), .B(n447), .X(n313) );
  SEN_ND3_S_0P5 U414 ( .A1(n863), .A2(n862), .A3(n900), .X(n314) );
  SEN_ND3_S_0P5 U415 ( .A1(n312), .A2(n313), .A3(n314), .X(Z[22]) );
  SEN_NR3_0P5 U416 ( .A1(n865), .A2(n866), .A3(n919), .X(n315) );
  SEN_OAOI211_0P5 U417 ( .A1(B[23]), .A2(A[23]), .B(n447), .C(n315), .X(n316)
         );
  SEN_ND2_0P5 U418 ( .A1(n864), .A2(n917), .X(n317) );
  SEN_OAI211_0P5 U419 ( .A1(n867), .A2(n926), .B1(n316), .B2(n317), .X(Z[23])
         );
  SEN_OR2_1 U420 ( .A1(n741), .A2(n740), .X(n514) );
  SEN_INV_0P5 U421 ( .A(n906), .X(n318) );
  SEN_OAI22_0P5 U422 ( .A1(n871), .A2(n897), .B1(n870), .B2(n318), .X(n319) );
  SEN_OAOI211_0P5 U423 ( .A1(A[24]), .A2(B[24]), .B(n447), .C(n319), .X(n320)
         );
  SEN_OAI31_0P5 U424 ( .A1(n868), .A2(n869), .A3(n919), .B(n320), .X(Z[24]) );
  SEN_AN2_1 U425 ( .A1(n346), .A2(n790), .X(n363) );
  SEN_AO2BB2_0P5 U426 ( .A1(n875), .A2(n897), .B1(n874), .B2(n906), .X(n321)
         );
  SEN_OAOI211_0P5 U427 ( .A1(B[25]), .A2(A[25]), .B(n446), .C(n321), .X(n322)
         );
  SEN_OAI31_0P5 U428 ( .A1(n872), .A2(n426), .A3(n919), .B(n322), .X(Z[25]) );
  SEN_AN2_1 U429 ( .A1(n509), .A2(n514), .X(n510) );
  SEN_MUX2_DG_1 U430 ( .D0(n601), .D1(n602), .S(n603), .X(n604) );
  SEN_OA2BB2_0P5 U431 ( .A1(n806), .A2(n549), .B1(n548), .B2(n806), .X(n550)
         );
  SEN_OA2BB2_0P5 U432 ( .A1(n675), .A2(n676), .B1(n674), .B2(n675), .X(n677)
         );
  SEN_AOI21_0P5 U433 ( .A1(n329), .A2(n337), .B(n648), .X(n323) );
  SEN_ND2_0P5 U434 ( .A1(n874), .A2(n323), .X(n649) );
  SEN_EN2_0P5 U435 ( .A1(n599), .A2(n756), .X(n753) );
  SEN_EO2_S_0P5 U436 ( .A1(n901), .A2(n899), .X(n907) );
  SEN_AO2BB2_0P5 U437 ( .A1(n898), .A2(n897), .B1(n896), .B2(n333), .X(n324)
         );
  SEN_OAOI211_0P5 U438 ( .A1(A[28]), .A2(B[28]), .B(n447), .C(n324), .X(n325)
         );
  SEN_OAI31_0P5 U439 ( .A1(n894), .A2(n895), .A3(n919), .B(n325), .X(Z[28]) );
  SEN_INV_S_1 U440 ( .A(n855), .X(n326) );
  SEN_OAI21_3 U441 ( .A1(n661), .A2(n641), .B(n663), .X(n635) );
  SEN_AN2_S_1 U442 ( .A1(n533), .A2(n498), .X(n327) );
  SEN_INV_S_1 U443 ( .A(n428), .X(n446) );
  SEN_OR2_1 U444 ( .A1(n693), .A2(n696), .X(n428) );
  SEN_OR4_1 U445 ( .A1(n646), .A2(n874), .A3(n329), .A4(n648), .X(n328) );
  SEN_MUXI2_S_2 U446 ( .D0(n442), .D1(n344), .S(B[16]), .X(n818) );
  SEN_EN2_S_2 U447 ( .A1(n400), .A2(n401), .X(n909) );
  SEN_ND2_G_4 U448 ( .A1(n697), .A2(n921), .X(n701) );
  SEN_NR2_T_3 U449 ( .A1(n697), .A2(n921), .X(n699) );
  SEN_ND2_T_1 U450 ( .A1(n563), .A2(n562), .X(n564) );
  SEN_ND2_S_2 U451 ( .A1(n824), .A2(n795), .X(n540) );
  SEN_ND4_S_3 U452 ( .A1(n534), .A2(n737), .A3(n789), .A4(n816), .X(n539) );
  SEN_ND2_S_2 U453 ( .A1(n609), .A2(n608), .X(n610) );
  SEN_EN2_1 U454 ( .A1(n738), .A2(n538), .X(n739) );
  SEN_ND2_T_4 U455 ( .A1(n394), .A2(n330), .X(n631) );
  SEN_OAI21_G_1 U456 ( .A1(n715), .A2(n332), .B(n714), .X(Z[1]) );
  SEN_AOI21_G_1 U457 ( .A1(n891), .A2(n906), .B(n890), .X(n892) );
  SEN_ND2_S_1 U458 ( .A1(n792), .A2(n906), .X(n793) );
  SEN_ND2_4 U459 ( .A1(n575), .A2(n585), .X(n588) );
  SEN_INV_1 U460 ( .A(n576), .X(n431) );
  SEN_INV_0P8 U461 ( .A(n738), .X(n745) );
  SEN_INV_2 U462 ( .A(n863), .X(n659) );
  SEN_INV_0P8 U463 ( .A(n723), .X(n730) );
  SEN_NR3_1 U464 ( .A1(n818), .A2(n817), .A3(n919), .X(n819) );
  SEN_INV_2 U465 ( .A(n498), .X(n810) );
  SEN_INV_2 U466 ( .A(n862), .X(n660) );
  SEN_EN2_1 U467 ( .A1(n865), .A2(n866), .X(n867) );
  SEN_NR2_T_2 U468 ( .A1(n833), .A2(n832), .X(n555) );
  SEN_INV_1P25 U469 ( .A(n854), .X(n590) );
  SEN_INV_0P5 U470 ( .A(n920), .X(n385) );
  SEN_ND2_2 U471 ( .A1(n443), .A2(n412), .X(n413) );
  SEN_ND2_G_1 U472 ( .A1(SEL), .A2(n686), .X(n457) );
  SEN_INV_6 U473 ( .A(n682), .X(n437) );
  SEN_AOI21_G_1 U474 ( .A1(n688), .A2(n687), .B(n686), .X(n926) );
  SEN_ND3_T_3 U475 ( .A1(n455), .A2(n454), .A3(n453), .X(n682) );
  SEN_NR2_G_1 U476 ( .A1(n331), .A2(n422), .X(n687) );
  SEN_ND2_T_0P5 U477 ( .A1(n331), .A2(n422), .X(n700) );
  SEN_AOI211_G_2 U478 ( .A1(n386), .A2(n917), .B1(n387), .B2(n388), .X(n374)
         );
  SEN_AOI211_G_2 U479 ( .A1(n699), .A2(n698), .B1(n383), .B2(n382), .X(n381)
         );
  SEN_OAI211_0P5 U480 ( .A1(n926), .A2(n925), .B1(n924), .B2(n923), .X(Z[31])
         );
  SEN_OAI211_0P5 U481 ( .A1(n926), .A2(n916), .B1(n915), .B2(n914), .X(Z[30])
         );
  SEN_EO2_3 U482 ( .A1(n843), .A2(n570), .X(n846) );
  SEN_ND3_T_2 U483 ( .A1(n679), .A2(n867), .A3(n417), .X(n673) );
  SEN_ND2_0P65 U484 ( .A1(n910), .A2(n917), .X(n915) );
  SEN_ND2_S_1 U485 ( .A1(n918), .A2(n917), .X(n924) );
  SEN_OAI211_0P5 U486 ( .A1(n926), .A2(n775), .B1(n774), .B2(n773), .X(Z[9])
         );
  SEN_NR3_T_2 U487 ( .A1(n739), .A2(n540), .A3(n539), .X(n565) );
  SEN_EN2_S_3 U488 ( .A1(n430), .A2(n644), .X(n893) );
  SEN_OAI211_0P5 U489 ( .A1(n926), .A2(n768), .B1(n767), .B2(n766), .X(Z[8])
         );
  SEN_NR2_G_2 U490 ( .A1(n607), .A2(n606), .X(n769) );
  SEN_OAI211_0P5 U491 ( .A1(n926), .A2(n745), .B1(n744), .B2(n743), .X(Z[5])
         );
  SEN_NR2_S_4 U492 ( .A1(n631), .A2(n665), .X(n641) );
  SEN_ND2_3 U493 ( .A1(n349), .A2(n372), .X(n370) );
  SEN_OAI211_0P5 U494 ( .A1(n926), .A2(n760), .B1(n759), .B2(n758), .X(Z[7])
         );
  SEN_ND2_4 U495 ( .A1(n497), .A2(n533), .X(n566) );
  SEN_ND4_S_3 U496 ( .A1(n782), .A2(n722), .A3(n715), .A4(n525), .X(n529) );
  SEN_OAI211_0P5 U497 ( .A1(n926), .A2(n752), .B1(n751), .B2(n750), .X(Z[6])
         );
  SEN_OAI211_0P5 U498 ( .A1(n926), .A2(n730), .B1(n729), .B2(n728), .X(Z[3])
         );
  SEN_ND2_0P65 U499 ( .A1(n724), .A2(n917), .X(n729) );
  SEN_ND2_T_2 U500 ( .A1(n366), .A2(n367), .X(n361) );
  SEN_INV_4 U501 ( .A(n664), .X(n330) );
  SEN_ND2_4 U502 ( .A1(n499), .A2(n429), .X(n334) );
  SEN_INV_2 U503 ( .A(n481), .X(n369) );
  SEN_NR2_G_1 U504 ( .A1(n521), .A2(n508), .X(n528) );
  SEN_AOI211_3 U505 ( .A1(n504), .A2(n494), .B1(n495), .B2(n368), .X(n367) );
  SEN_INV_1 U506 ( .A(n891), .X(n430) );
  SEN_AOI21_G_1 U507 ( .A1(n882), .A2(n906), .B(n881), .X(n883) );
  SEN_OAOI211_1 U508 ( .A1(B[15]), .A2(A[15]), .B(n446), .C(n812), .X(n815) );
  SEN_NR2_G_3 U509 ( .A1(n588), .A2(n576), .X(n578) );
  SEN_OAOI211_1 U510 ( .A1(B[14]), .A2(A[14]), .B(n447), .C(n805), .X(n808) );
  SEN_NR2_G_3 U511 ( .A1(n486), .A2(n485), .X(n487) );
  SEN_AOI21_G_0P75 U512 ( .A1(n907), .A2(n906), .B(n905), .X(n908) );
  SEN_NR2_T_2 U513 ( .A1(n478), .A2(n483), .X(n482) );
  SEN_OAOI211_1 U514 ( .A1(B[13]), .A2(A[13]), .B(n446), .C(n798), .X(n801) );
  SEN_ND2_0P8 U515 ( .A1(n821), .A2(n906), .X(n822) );
  SEN_AOAI211_1 U516 ( .A1(n904), .A2(n903), .B(n428), .C(n902), .X(n905) );
  SEN_AOAI211_1 U517 ( .A1(n880), .A2(n879), .B(n428), .C(n878), .X(n881) );
  SEN_AOAI211_1 U518 ( .A1(n889), .A2(n888), .B(n428), .C(n887), .X(n890) );
  SEN_INV_1 U519 ( .A(n650), .X(n337) );
  SEN_EO2_1 U520 ( .A1(n619), .A2(n618), .X(n882) );
  SEN_NR3_1 U521 ( .A1(n797), .A2(n796), .A3(n445), .X(n798) );
  SEN_OAOI211_1 U522 ( .A1(B[6]), .A2(A[6]), .B(n447), .C(n749), .X(n750) );
  SEN_ND2_T_4 U523 ( .A1(n602), .A2(n477), .X(n483) );
  SEN_OAOI211_1 U524 ( .A1(B[3]), .A2(A[3]), .B(n446), .C(n727), .X(n728) );
  SEN_NR3_1 U525 ( .A1(n811), .A2(n810), .A3(n445), .X(n812) );
  SEN_INV_0P8 U526 ( .A(n753), .X(n760) );
  SEN_INV_1 U527 ( .A(n580), .X(n582) );
  SEN_OAOI211_1 U528 ( .A1(A[12]), .A2(B[12]), .B(n446), .C(n791), .X(n794) );
  SEN_INV_1 U529 ( .A(n820), .X(n821) );
  SEN_OAOI211_1 U530 ( .A1(B[16]), .A2(A[16]), .B(n447), .C(n819), .X(n823) );
  SEN_ND2_3 U531 ( .A1(n548), .A2(n493), .X(n495) );
  SEN_EN2_1 U532 ( .A1(n803), .A2(n804), .X(n544) );
  SEN_NR3_1 U533 ( .A1(n804), .A2(n803), .A3(n445), .X(n805) );
  SEN_INV_0P8 U534 ( .A(n761), .X(n768) );
  SEN_OAI22_T_2 U535 ( .A1(n784), .A2(n783), .B1(n346), .B2(n790), .X(n368) );
  SEN_OAOI211_1 U536 ( .A1(B[4]), .A2(A[4]), .B(n446), .C(n733), .X(n736) );
  SEN_OAOI211_1 U537 ( .A1(A[8]), .A2(B[8]), .B(n446), .C(n765), .X(n766) );
  SEN_AN2_1 U538 ( .A1(n901), .A2(n899), .X(n402) );
  SEN_INV_1 U539 ( .A(n506), .X(n507) );
  SEN_ND2_3 U540 ( .A1(n473), .A2(n472), .X(n484) );
  SEN_INV_1 U541 ( .A(n867), .X(n675) );
  SEN_OAOI211_1 U542 ( .A1(B[31]), .A2(A[31]), .B(n447), .C(n922), .X(n923) );
  SEN_AN2_1 U543 ( .A1(n568), .A2(n556), .X(n579) );
  SEN_INV_1 U544 ( .A(n886), .X(n639) );
  SEN_OAOI211_1 U545 ( .A1(A[7]), .A2(B[7]), .B(n447), .C(n757), .X(n758) );
  SEN_OAOI211_1 U546 ( .A1(A[5]), .A2(B[5]), .B(n446), .C(n742), .X(n743) );
  SEN_INV_3 U547 ( .A(n425), .X(n426) );
  SEN_INV_1 U548 ( .A(n512), .X(n513) );
  SEN_OAOI211_1 U549 ( .A1(A[2]), .A2(B[2]), .B(n446), .C(n718), .X(n721) );
  SEN_OAOI211_1 U550 ( .A1(A[17]), .A2(B[17]), .B(n447), .C(n827), .X(n830) );
  SEN_INV_1 U551 ( .A(n775), .X(n603) );
  SEN_INV_1 U552 ( .A(n877), .X(n618) );
  SEN_OAOI211_1 U553 ( .A1(A[30]), .A2(B[30]), .B(n447), .C(n913), .X(n914) );
  SEN_AN2_1 U554 ( .A1(n863), .A2(n862), .X(n676) );
  SEN_OAOI211_1 U555 ( .A1(A[9]), .A2(B[9]), .B(n446), .C(n772), .X(n773) );
  SEN_OAOI211_1 U556 ( .A1(A[10]), .A2(B[10]), .B(n446), .C(n778), .X(n781) );
  SEN_INV_1 U557 ( .A(n612), .X(n613) );
  SEN_OAOI211_1 U558 ( .A1(B[18]), .A2(A[18]), .B(n447), .C(n834), .X(n838) );
  SEN_NR3_1 U559 ( .A1(n335), .A2(n725), .A3(n445), .X(n727) );
  SEN_OAOI211_1 U560 ( .A1(B[11]), .A2(A[11]), .B(n446), .C(n785), .X(n788) );
  SEN_AOI21_G_1 U561 ( .A1(n713), .A2(n906), .B(n712), .X(n714) );
  SEN_NR2_T_3 U562 ( .A1(n536), .A2(n463), .X(n509) );
  SEN_OAOI211_1 U563 ( .A1(A[21]), .A2(B[21]), .B(n446), .C(n856), .X(n859) );
  SEN_OAOI211_1 U564 ( .A1(A[19]), .A2(B[19]), .B(n447), .C(n842), .X(n845) );
  SEN_OAOI211_1 U565 ( .A1(B[20]), .A2(A[20]), .B(n447), .C(n849), .X(n852) );
  SEN_INV_1 U566 ( .A(n835), .X(n836) );
  SEN_NR3_1 U567 ( .A1(n912), .A2(n911), .A3(n919), .X(n913) );
  SEN_EN2_DG_2 U568 ( .A1(n911), .A2(n912), .X(n916) );
  SEN_NR3_1 U569 ( .A1(n921), .A2(n920), .A3(n919), .X(n922) );
  SEN_NR2_G_2 U570 ( .A1(n841), .A2(n840), .X(n612) );
  SEN_INV_1 U571 ( .A(n885), .X(n640) );
  SEN_ND2_T_2 U572 ( .A1(n411), .A2(n413), .X(n863) );
  SEN_ND2_2 U573 ( .A1(n726), .A2(n725), .X(n468) );
  SEN_AOAI211_1 U574 ( .A1(n711), .A2(n710), .B(n428), .C(n709), .X(n712) );
  SEN_NR2_G_3 U575 ( .A1(n826), .A2(n825), .X(n571) );
  SEN_EO2_1 U576 ( .A1(n523), .A2(n522), .X(n713) );
  SEN_INV_1 U577 ( .A(n817), .X(n638) );
  SEN_ND2_2 U578 ( .A1(n404), .A2(n406), .X(n498) );
  SEN_ND2_3 U579 ( .A1(n458), .A2(n457), .X(n692) );
  SEN_INV_S_2 U580 ( .A(n707), .X(n523) );
  SEN_INV_S_2 U581 ( .A(n763), .X(n475) );
  SEN_INV_12 U582 ( .A(n437), .X(n435) );
  SEN_OAI21_T_0P5 U583 ( .A1(A[0]), .A2(B[0]), .B(n447), .X(n390) );
  SEN_INV_4 U584 ( .A(n683), .X(n440) );
  SEN_MUXI2_D_1 U585 ( .D0(n688), .D1(n461), .S(n424), .X(n462) );
  SEN_INV_S_0P5 U586 ( .A(n456), .X(n336) );
  SEN_ND2_2 U587 ( .A1(n451), .A2(n671), .X(n454) );
  SEN_ND2_3 U588 ( .A1(n696), .A2(n671), .X(n460) );
  SEN_INV_10 U589 ( .A(n434), .X(n705) );
  SEN_INV_1 U590 ( .A(B[15]), .X(n496) );
  SEN_INV_1 U591 ( .A(B[26]), .X(n879) );
  SEN_INV_1 U592 ( .A(A[29]), .X(n904) );
  SEN_INV_1 U593 ( .A(A[1]), .X(n710) );
  SEN_INV_1 U594 ( .A(A[14]), .X(n492) );
  SEN_INV_1 U595 ( .A(B[27]), .X(n889) );
  SEN_INV_1 U596 ( .A(B[1]), .X(n711) );
  SEN_INV_1 U597 ( .A(B[14]), .X(n491) );
  SEN_INV_1 U598 ( .A(B[29]), .X(n903) );
  SEN_INV_1 U599 ( .A(B[13]), .X(n489) );
  SEN_INV_1 U600 ( .A(A[27]), .X(n888) );
  SEN_INV_1 U601 ( .A(A[13]), .X(n490) );
  SEN_INV_1 U602 ( .A(A[26]), .X(n880) );
  SEN_INV_4 U603 ( .A(INST[2]), .X(n331) );
  SEN_INV_1 U604 ( .A(n917), .X(n332) );
  SEN_MUXI2_DG_2 U605 ( .D0(n345), .D1(n444), .S(n491), .X(n542) );
  SEN_MUXI2_DG_2 U606 ( .D0(n345), .D1(n444), .S(n489), .X(n561) );
  SEN_ND2_T_4 U607 ( .A1(n349), .A2(n431), .X(n432) );
  SEN_ND2_T_5 U608 ( .A1(n348), .A2(n498), .X(n349) );
  SEN_AOI211_2 U609 ( .A1(n706), .A2(n331), .B1(n418), .B2(n705), .X(n378) );
  SEN_ND2_G_3 U610 ( .A1(n702), .A2(n701), .X(n706) );
  SEN_MUXI2_D_1 U611 ( .D0(n443), .D1(n441), .S(B[24]), .X(n869) );
  SEN_ND2_T_1 U612 ( .A1(n441), .A2(B[22]), .X(n411) );
  SEN_INV_4 U613 ( .A(n755), .X(n599) );
  SEN_MUXI2_DG_2 U614 ( .D0(n442), .D1(n344), .S(B[2]), .X(n717) );
  SEN_MUXI2_DG_2 U615 ( .D0(n442), .D1(n344), .S(B[3]), .X(n726) );
  SEN_MUXI2_DG_2 U616 ( .D0(n442), .D1(n344), .S(B[4]), .X(n732) );
  SEN_MUXI2_DG_2 U617 ( .D0(n442), .D1(n344), .S(B[5]), .X(n741) );
  SEN_MUXI2_DG_3 U618 ( .D0(n442), .D1(n344), .S(B[6]), .X(n748) );
  SEN_MUXI2_DG_3 U619 ( .D0(n442), .D1(n344), .S(B[8]), .X(n764) );
  SEN_MUXI2_DG_2 U620 ( .D0(n442), .D1(n344), .S(B[10]), .X(n777) );
  SEN_MUXI2_DG_3 U621 ( .D0(n442), .D1(n344), .S(B[7]), .X(n756) );
  SEN_MAJI3_2 U622 ( .A1(n725), .A2(n335), .A3(n531), .X(n537) );
  SEN_INV_2 U623 ( .A(n631), .X(n627) );
  SEN_AN3_S_2 U624 ( .A1(n488), .A2(n487), .A3(n514), .X(n429) );
  SEN_ND3_T_2 U625 ( .A1(n348), .A2(n330), .A3(n669), .X(n396) );
  SEN_ND2_T_4 U626 ( .A1(n566), .A2(n575), .X(n611) );
  SEN_ND2_T_4 U627 ( .A1(n642), .A2(n634), .X(n661) );
  SEN_AO2BB2_4 U628 ( .A1(n598), .A2(n599), .B1(n748), .B2(n747), .X(n474) );
  SEN_INV_3 U629 ( .A(n756), .X(n598) );
  SEN_MUXI2_S_4 U630 ( .D0(n438), .D1(n435), .S(A[7]), .X(n755) );
  SEN_NR3_T_3 U631 ( .A1(n499), .A2(n340), .A3(n481), .X(n360) );
  SEN_BUF_6 U632 ( .A(INST[3]), .X(n434) );
  SEN_MUX2_G_4 U633 ( .D0(n440), .D1(n437), .S(A[8]), .X(n763) );
  SEN_INV_3 U634 ( .A(n341), .X(n671) );
  SEN_ND3_T_2 U635 ( .A1(n500), .A2(n494), .A3(n502), .X(n481) );
  SEN_MUXI2_DG_4 U636 ( .D0(n439), .D1(n436), .S(A[18]), .X(n832) );
  SEN_MUXI2_DG_3 U637 ( .D0(n439), .D1(n436), .S(A[23]), .X(n865) );
  SEN_NR3_0P5 U638 ( .A1(n764), .A2(n763), .A3(n445), .X(n765) );
  SEN_MUXI2_DG_2 U639 ( .D0(n438), .D1(n435), .S(A[4]), .X(n731) );
  SEN_INV_2P5 U640 ( .A(n435), .X(n338) );
  SEN_MUXI2_DG_5 U641 ( .D0(n438), .D1(n435), .S(A[0]), .X(n458) );
  SEN_OAOI211_3 U642 ( .A1(n549), .A2(n363), .B(n364), .C(n365), .X(n362) );
  SEN_NR3_0P5 U643 ( .A1(n833), .A2(n832), .A3(n919), .X(n834) );
  SEN_NR3_0P5 U644 ( .A1(n848), .A2(n847), .A3(n919), .X(n849) );
  SEN_EO2_DG_1 U645 ( .A1(n840), .A2(n841), .X(n843) );
  SEN_NR3_0P5 U646 ( .A1(n826), .A2(n825), .A3(n919), .X(n827) );
  SEN_NR3_0P5 U647 ( .A1(n717), .A2(n716), .A3(n445), .X(n718) );
  SEN_ND2_T_1 U648 ( .A1(n784), .A2(n783), .X(n494) );
  SEN_NR3_0P5 U649 ( .A1(n777), .A2(n776), .A3(n445), .X(n778) );
  SEN_NR3_0P5 U650 ( .A1(n346), .A2(n790), .A3(n445), .X(n791) );
  SEN_NR3_0P5 U651 ( .A1(n756), .A2(n755), .A3(n445), .X(n757) );
  SEN_EO2_0P5 U652 ( .A1(n740), .A2(n741), .X(n738) );
  SEN_ND3_S_4 U653 ( .A1(n578), .A2(n811), .A3(n810), .X(n587) );
  SEN_ND2_S_1P5 U654 ( .A1(n869), .A2(n868), .X(n647) );
  SEN_BUF_6 U655 ( .A(INST[1]), .X(n341) );
  SEN_NR2_T_3 U656 ( .A1(n726), .A2(n725), .X(n463) );
  SEN_ND2_2 U657 ( .A1(n474), .A2(n484), .X(n478) );
  SEN_ND2_T_4 U658 ( .A1(n598), .A2(n599), .X(n477) );
  SEN_ND2_2 U659 ( .A1(n561), .A2(n560), .X(n548) );
  SEN_MUXI2_S_6 U660 ( .D0(n438), .D1(n435), .S(A[9]), .X(n770) );
  SEN_INV_12 U661 ( .A(n343), .X(n344) );
  SEN_INV_10 U662 ( .A(n355), .X(n343) );
  SEN_INV_10 U663 ( .A(n440), .X(n438) );
  SEN_OAI21_8 U664 ( .A1(n356), .A2(n422), .B(n459), .X(n355) );
  SEN_NR2_T_4 U665 ( .A1(n357), .A2(n358), .X(n356) );
  SEN_MUXI2_S_4 U666 ( .D0(n433), .D1(n342), .S(n452), .X(n358) );
  SEN_ND2_2 U667 ( .A1(n408), .A2(n689), .X(n410) );
  SEN_INV_3 U668 ( .A(n482), .X(n501) );
  SEN_ND2_T_2 U669 ( .A1(n347), .A2(n666), .X(n394) );
  SEN_ND3_T_1 U670 ( .A1(n376), .A2(n375), .A3(n374), .X(Z[0]) );
  SEN_ND2_G_4 U671 ( .A1(n433), .A2(n341), .X(n342) );
  SEN_NR4_1 U672 ( .A1(n910), .A2(n341), .A3(n331), .A4(n705), .X(n379) );
  SEN_OAI211_1 U673 ( .A1(n341), .A2(n706), .B1(n377), .B2(n378), .X(n376) );
  SEN_NR2_2 U674 ( .A1(n451), .A2(n341), .X(n683) );
  SEN_ND2_S_1P5 U675 ( .A1(n450), .A2(n341), .X(n455) );
  SEN_NR2_1 U676 ( .A1(n696), .A2(n341), .X(n698) );
  SEN_ND2_G_1 U677 ( .A1(n331), .A2(n341), .X(n690) );
  SEN_OAOI211_G_1 U678 ( .A1(n702), .A2(n336), .B(n381), .C(n700), .X(n380) );
  SEN_NR2_S_2 U679 ( .A1(n342), .A2(n331), .X(n448) );
  SEN_MUXI2_S_2 U680 ( .D0(n343), .D1(n444), .S(n711), .X(n708) );
  SEN_INV_5 U681 ( .A(n343), .X(n441) );
  SEN_INV_4 U682 ( .A(n344), .X(n345) );
  SEN_MUXI2_DG_2 U683 ( .D0(n344), .D1(n442), .S(n409), .X(n689) );
  SEN_MUXI2_S_1 U684 ( .D0(n442), .D1(n344), .S(B[21]), .X(n855) );
  SEN_MUXI2_S_4 U685 ( .D0(n442), .D1(n344), .S(B[11]), .X(n784) );
  SEN_MUX2_S_2 U686 ( .D0(n444), .D1(n345), .S(B[12]), .X(n346) );
  SEN_AOI21B_2 U687 ( .A1(n345), .A2(B[15]), .B(n403), .X(n533) );
  SEN_MUXI2_S_1 U688 ( .D0(n345), .D1(n444), .S(n903), .X(n901) );
  SEN_OAI21_S_2 U689 ( .A1(n546), .A2(n790), .B(n346), .X(n563) );
  SEN_OAI21_5 U690 ( .A1(n360), .A2(n361), .B(n362), .X(n347) );
  SEN_INV_3 U691 ( .A(n347), .X(n348) );
  SEN_EO2_1 U692 ( .A1(n813), .A2(n347), .X(n816) );
  SEN_ND2_2 U693 ( .A1(n347), .A2(n810), .X(n497) );
  SEN_ND2_2 U694 ( .A1(n349), .A2(n566), .X(n636) );
  SEN_OAI21_5 U695 ( .A1(n611), .A2(n370), .B(n371), .X(n350) );
  SEN_NR2_T_3 U696 ( .A1(n350), .A2(n854), .X(n672) );
  SEN_NR2_T_1P5 U697 ( .A1(n351), .A2(n672), .X(n373) );
  SEN_MUXI2_S_1 U698 ( .D0(n673), .D1(n678), .S(n351), .X(n681) );
  SEN_EO2_2 U699 ( .A1(n861), .A2(n373), .X(n352) );
  SEN_INV_3 U700 ( .A(n352), .X(n353) );
  SEN_ND3_T_1 U701 ( .A1(n352), .A2(n704), .A3(n393), .X(n392) );
  SEN_NR4_6 U702 ( .A1(n695), .A2(n864), .A3(n353), .A4(n909), .X(n354) );
  SEN_AOI31_1 U703 ( .A1(n354), .A2(n379), .A3(n703), .B(n380), .X(n375) );
  SEN_ND3_T_2 U704 ( .A1(n354), .A2(n704), .A3(n703), .X(n377) );
  SEN_ND2_S_2 U705 ( .A1(n460), .A2(n690), .X(n357) );
  SEN_ND3_2 U706 ( .A1(n488), .A2(n487), .A3(n514), .X(n359) );
  SEN_NR2_1 U707 ( .A1(n542), .A2(n541), .X(n365) );
  SEN_INV_3 U708 ( .A(n495), .X(n364) );
  SEN_ND3_2 U709 ( .A1(n369), .A2(n501), .A3(n359), .X(n366) );
  SEN_AN2_S_1 U710 ( .A1(n585), .A2(n431), .X(n372) );
  SEN_AOI21_S_1 U711 ( .A1(n614), .A2(n585), .B(n580), .X(n371) );
  SEN_ND2_G_1 U712 ( .A1(n385), .A2(n698), .X(n384) );
  SEN_INV_1 U713 ( .A(n689), .X(n391) );
  SEN_NR4_1 U714 ( .A1(n909), .A2(n418), .A3(n671), .A4(n700), .X(n393) );
  SEN_AOI21_2 U715 ( .A1(n697), .A2(n921), .B(n384), .X(n383) );
  SEN_ND3_S_0P5 U716 ( .A1(n391), .A2(n900), .A3(n692), .X(n389) );
  SEN_OAI211_1 U717 ( .A1(n694), .A2(n926), .B1(n389), .B2(n390), .X(n388) );
  SEN_NR4_3 U718 ( .A1(n695), .A2(n392), .A3(n864), .A4(n918), .X(n387) );
  SEN_INV_S_1 U719 ( .A(n525), .X(n386) );
  SEN_ND2B_4 U720 ( .A(n699), .B(n920), .X(n702) );
  SEN_AN2_6 U721 ( .A1(n417), .A2(n592), .X(n622) );
  SEN_AOI21B_3 U722 ( .A1(n631), .A2(n622), .B(n630), .X(n646) );
  SEN_NR2_2 U723 ( .A1(n646), .A2(n329), .X(n395) );
  SEN_INV_AS_2 U724 ( .A(n395), .X(n594) );
  SEN_INV_2 U725 ( .A(n630), .X(n621) );
  SEN_AOI31_3 U726 ( .A1(n330), .A2(n668), .A3(n669), .B(n667), .X(n397) );
  SEN_ND2_G_1 U727 ( .A1(n662), .A2(n663), .X(n670) );
  SEN_INV_1 U728 ( .A(n670), .X(n398) );
  SEN_ND2_T_4 U729 ( .A1(n661), .A2(n398), .X(n399) );
  SEN_ND3_T_4 U730 ( .A1(n396), .A2(n397), .A3(n399), .X(n400) );
  SEN_INV_1 U731 ( .A(n907), .X(n401) );
  SEN_OAI22_T_4 U732 ( .A1(n400), .A2(n402), .B1(n901), .B2(n899), .X(n685) );
  SEN_ND2_T_1 U733 ( .A1(n444), .A2(n496), .X(n403) );
  SEN_ND2_T_1 U734 ( .A1(n436), .A2(A[15]), .X(n404) );
  SEN_INV_1 U735 ( .A(A[15]), .X(n405) );
  SEN_ND2_T_1 U736 ( .A1(n438), .A2(n405), .X(n406) );
  SEN_ND2_T_1 U737 ( .A1(n438), .A2(n331), .X(n407) );
  SEN_ND2B_V1_3 U738 ( .A(n442), .B(n407), .X(n464) );
  SEN_ND2_G_1 U739 ( .A1(n692), .A2(n464), .X(n408) );
  SEN_INV_1 U740 ( .A(B[0]), .X(n409) );
  SEN_ND2_S_1P5 U741 ( .A1(n465), .A2(n410), .X(n467) );
  SEN_ND2_T_1P5 U742 ( .A1(n507), .A2(n410), .X(n524) );
  SEN_INV_1 U743 ( .A(B[22]), .X(n412) );
  SEN_INV_1 U744 ( .A(A[22]), .X(n415) );
  SEN_INV_2 U745 ( .A(n676), .X(n417) );
  SEN_INV_2 U746 ( .A(SEL), .X(n452) );
  SEN_ND2_T_1 U747 ( .A1(n501), .A2(n500), .X(n518) );
  SEN_INV_S_1 U748 ( .A(n696), .X(n418) );
  SEN_BUF_S_6 U749 ( .A(INST[0]), .X(n433) );
  SEN_ND2_S_2 U750 ( .A1(n705), .A2(n433), .X(n451) );
  SEN_ND3_S_4 U751 ( .A1(n853), .A2(n884), .A3(n898), .X(n655) );
  SEN_OAI21_3 U752 ( .A1(n567), .A2(n432), .B(n419), .X(n573) );
  SEN_MAJ3_2 U753 ( .A1(n638), .A2(n637), .A3(n636), .X(n427) );
  SEN_EO2_2 U754 ( .A1(n820), .A2(n636), .X(n824) );
  SEN_NR3_0P5 U755 ( .A1(n732), .A2(n731), .A3(n445), .X(n733) );
  SEN_NR2_T_4 U756 ( .A1(n655), .A2(n654), .X(n656) );
  SEN_ND4_S_4 U757 ( .A1(n565), .A2(n809), .A3(n860), .A4(n802), .X(n596) );
  SEN_MUXI2_DG_3 U758 ( .D0(n438), .D1(n435), .S(A[12]), .X(n790) );
  SEN_MUXI2_S_2 U759 ( .D0(n438), .D1(n435), .S(A[16]), .X(n817) );
  SEN_MUXI2_S_2 U760 ( .D0(n438), .D1(n435), .S(A[10]), .X(n776) );
  SEN_ND3_T_4 U761 ( .A1(n831), .A2(n653), .A3(n875), .X(n654) );
  SEN_ND2_S_0P5 U762 ( .A1(n739), .A2(n917), .X(n744) );
  SEN_ND3_4 U763 ( .A1(n471), .A2(n470), .A3(n469), .X(n499) );
  SEN_ND2_2 U764 ( .A1(n509), .A2(n511), .X(n469) );
  SEN_AOI22_1 U765 ( .A1(n825), .A2(n826), .B1(n818), .B2(n817), .X(n419) );
  SEN_NR3_0P5 U766 ( .A1(n420), .A2(n747), .A3(n445), .X(n749) );
  SEN_EO2_2 U767 ( .A1(n896), .A2(n635), .X(n898) );
  SEN_INV_2 U768 ( .A(n764), .X(n476) );
  SEN_OAI21_S_3 U769 ( .A1(n452), .A2(n434), .B(n696), .X(n453) );
  SEN_MUXI2_DG_4 U770 ( .D0(n438), .D1(n435), .S(A[11]), .X(n783) );
  SEN_OAI21_G_2 U771 ( .A1(n449), .A2(n434), .B(n424), .X(n450) );
  SEN_INV_AS_2 U772 ( .A(n611), .X(n616) );
  SEN_NR3_T_2 U773 ( .A1(n746), .A2(n529), .A3(n724), .X(n534) );
  SEN_MUXI2_S_2 U774 ( .D0(n438), .D1(n435), .S(A[2]), .X(n716) );
  SEN_MUXI2_S_4 U775 ( .D0(n438), .D1(n435), .S(A[6]), .X(n747) );
  SEN_INV_S_1 U776 ( .A(n436), .X(n421) );
  SEN_ND3_T_4 U777 ( .A1(n456), .A2(n424), .A3(n422), .X(n459) );
  SEN_NR2_3 U778 ( .A1(n877), .A2(n876), .X(n628) );
  SEN_AOI22_T_3 U779 ( .A1(n633), .A2(n632), .B1(n877), .B2(n876), .X(n642) );
  SEN_INV_10 U780 ( .A(n705), .X(n422) );
  SEN_MUXI2_S_2 U781 ( .D0(n437), .D1(n440), .S(n710), .X(n707) );
  SEN_NR2_T_3 U782 ( .A1(n692), .A2(n464), .X(n506) );
  SEN_MAJI3_2 U783 ( .A1(n784), .A2(n783), .A3(n532), .X(n543) );
  SEN_EN2_DG_1 U784 ( .A1(n792), .A2(n543), .X(n795) );
  SEN_ND3_2 U785 ( .A1(n652), .A2(n328), .A3(n651), .X(n875) );
  SEN_EO2_2 U786 ( .A1(n753), .A2(n645), .X(n754) );
  SEN_ND2_G_4 U787 ( .A1(n645), .A2(n599), .X(n608) );
  SEN_MAJI3_3 U788 ( .A1(n420), .A2(n747), .A3(n597), .X(n645) );
  SEN_EN2_3 U789 ( .A1(n828), .A2(n427), .X(n831) );
  SEN_EN2_S_2 U790 ( .A1(n734), .A2(n537), .X(n737) );
  SEN_EN2_S_2 U791 ( .A1(n925), .A2(n697), .X(n918) );
  SEN_INV_2 U792 ( .A(n918), .X(n703) );
  SEN_ND3_T_4 U793 ( .A1(n658), .A2(n657), .A3(n656), .X(n695) );
  SEN_OAI211_0P5 U794 ( .A1(n795), .A2(n897), .B1(n794), .B2(n793), .X(Z[12])
         );
  SEN_INV_4 U795 ( .A(n331), .X(n424) );
  SEN_ND3_S_8 U796 ( .A1(n846), .A2(n839), .A3(n871), .X(n595) );
  SEN_OAI211_3 U797 ( .A1(n589), .A2(n588), .B1(n587), .B2(n586), .X(n664) );
  SEN_INV_AS_2 U798 ( .A(n873), .X(n425) );
  SEN_ND2_T_1P5 U799 ( .A1(n433), .A2(SEL), .X(n449) );
  SEN_ND2_T_4 U800 ( .A1(n632), .A2(n630), .X(n665) );
  SEN_NR2_T_4 U801 ( .A1(n629), .A2(n628), .X(n632) );
  SEN_NR3_T_2 U802 ( .A1(n329), .A2(n648), .A3(n623), .X(n620) );
  SEN_EN2_3 U803 ( .A1(n850), .A2(n617), .X(n853) );
  SEN_EO2_1 U804 ( .A1(n882), .A2(n626), .X(n884) );
  SEN_OAI21_T_3 U805 ( .A1(n622), .A2(n621), .B(n620), .X(n633) );
  SEN_ND3_T_2 U806 ( .A1(n467), .A2(n509), .A3(n466), .X(n471) );
  SEN_AOI21_2 U807 ( .A1(n708), .A2(n707), .B(n508), .X(n466) );
  SEN_NR3_0P5 U808 ( .A1(n841), .A2(n840), .A3(n919), .X(n842) );
  SEN_NR2_T_1 U809 ( .A1(n777), .A2(n776), .X(n504) );
  SEN_INV_2 U810 ( .A(n484), .X(n486) );
  SEN_INV_2 U811 ( .A(n672), .X(n679) );
  SEN_NR2_2 U812 ( .A1(n448), .A2(n705), .X(n684) );
  SEN_INV_5 U813 ( .A(n684), .X(n444) );
  SEN_INV_4 U814 ( .A(n771), .X(n473) );
  SEN_EO2_1 U815 ( .A1(n752), .A2(n597), .X(n746) );
  SEN_EO2_S_0P5 U816 ( .A1(n716), .A2(n717), .X(n719) );
  SEN_NR2_S_5 U817 ( .A1(n571), .A2(n555), .X(n575) );
  SEN_AN2_2 U818 ( .A1(n535), .A2(n512), .X(n470) );
  SEN_ND2_2 U819 ( .A1(n771), .A2(n770), .X(n479) );
  SEN_AOI21_3 U820 ( .A1(n647), .A2(n624), .B(n623), .X(n629) );
  SEN_ND2_T_1P5 U821 ( .A1(n426), .A2(n872), .X(n624) );
  SEN_ND2_2 U822 ( .A1(n764), .A2(n763), .X(n601) );
  SEN_ND2_G_3 U823 ( .A1(n476), .A2(n475), .X(n602) );
  SEN_EO2_2 U824 ( .A1(n799), .A2(n564), .X(n802) );
  SEN_NR2_T_3 U825 ( .A1(n612), .A2(n554), .X(n585) );
  SEN_NR2_2 U826 ( .A1(n553), .A2(n552), .X(n809) );
  SEN_NR2_T_3 U827 ( .A1(n596), .A2(n595), .X(n658) );
  SEN_ND2_2 U828 ( .A1(n526), .A2(n468), .X(n511) );
  SEN_INV_6 U829 ( .A(n437), .X(n436) );
  SEN_ND2_G_3 U830 ( .A1(n833), .A2(n832), .X(n568) );
  SEN_INV_AS_2 U831 ( .A(n566), .X(n567) );
  SEN_NR3_0P5 U832 ( .A1(n784), .A2(n783), .A3(n445), .X(n785) );
  SEN_MUXI2_S_3 U833 ( .D0(n438), .D1(n435), .S(A[3]), .X(n725) );
  SEN_ND2_2 U834 ( .A1(n591), .A2(n590), .X(n592) );
  SEN_INV_6 U835 ( .A(n444), .X(n442) );
  SEN_OAI21_S_3 U836 ( .A1(n645), .A2(n599), .B(n598), .X(n609) );
  SEN_EO2_2 U837 ( .A1(n761), .A2(n610), .X(n762) );
  SEN_EO2_2 U838 ( .A1(n835), .A2(n574), .X(n839) );
  SEN_AOI21_3 U839 ( .A1(n334), .A2(n505), .B(n504), .X(n532) );
  SEN_NR2_T_1P5 U840 ( .A1(n528), .A2(n527), .X(n530) );
  SEN_EO2_2 U841 ( .A1(n723), .A2(n530), .X(n724) );
  SEN_MUXI2_DG_3 U842 ( .D0(n443), .D1(n441), .S(B[23]), .X(n866) );
  SEN_MUXI2_DG_3 U843 ( .D0(n443), .D1(n441), .S(B[19]), .X(n841) );
  SEN_NR2_2 U844 ( .A1(n665), .A2(n670), .X(n669) );
  SEN_NR2_2 U845 ( .A1(n848), .A2(n847), .X(n554) );
  SEN_ND3_T_2 U846 ( .A1(n608), .A2(n602), .A3(n775), .X(n600) );
  SEN_INV_6 U847 ( .A(n440), .X(n439) );
  SEN_ND2_2 U848 ( .A1(n601), .A2(n479), .X(n480) );
  SEN_ND3_1 U849 ( .A1(n646), .A2(n874), .A3(n337), .X(n652) );
  SEN_MUXI2_S_3 U850 ( .D0(n443), .D1(n441), .S(B[18]), .X(n833) );
  SEN_OAI21_S_3 U851 ( .A1(n679), .A2(n678), .B(n677), .X(n680) );
  SEN_MUXI2_S_3 U852 ( .D0(n443), .D1(n441), .S(B[20]), .X(n848) );
  SEN_INV_2 U853 ( .A(n578), .X(n577) );
  SEN_NR2_2 U854 ( .A1(n769), .A2(n762), .X(n657) );
  SEN_ND2_T_1P5 U855 ( .A1(n517), .A2(n516), .X(n597) );
  SEN_AOI21_T_1 U856 ( .A1(n522), .A2(n523), .B(n506), .X(n465) );
  SEN_ND2_2 U857 ( .A1(n659), .A2(n660), .X(n674) );
  SEN_EN2_4 U858 ( .A1(n916), .A2(n685), .X(n704) );
  SEN_MUXI2_S_2 U859 ( .D0(n551), .D1(n547), .S(n563), .X(n553) );
  SEN_INV_4 U860 ( .A(n444), .X(n443) );
  SEN_OAI211_0P5 U861 ( .A1(n802), .A2(n897), .B1(n801), .B2(n800), .X(Z[13])
         );
  SEN_INV_2 U862 ( .A(n543), .X(n546) );
  SEN_INV_2 U863 ( .A(n770), .X(n472) );
  SEN_NR2_T_3 U864 ( .A1(n681), .A2(n680), .X(n864) );
  SEN_MAJI3_T_1 U865 ( .A1(n523), .A2(n522), .A3(n524), .X(n521) );
  SEN_INV_2 U866 ( .A(n530), .X(n531) );
  SEN_MAJI3_T_4 U867 ( .A1(n911), .A2(n912), .A3(n685), .X(n697) );
  SEN_OAI211_0P5 U868 ( .A1(n824), .A2(n897), .B1(n823), .B2(n822), .X(Z[16])
         );
  SEN_NR2_T_1P5 U869 ( .A1(n518), .A2(n503), .X(n505) );
  SEN_ND2_2 U870 ( .A1(n546), .A2(n790), .X(n562) );
  SEN_ND2_2 U871 ( .A1(n480), .A2(n484), .X(n500) );
  SEN_INV_2 U872 ( .A(n483), .X(n488) );
  SEN_EO2_2 U873 ( .A1(n870), .A2(n594), .X(n871) );
  SEN_ND2_2 U874 ( .A1(n569), .A2(n568), .X(n570) );
  SEN_AOAI211_3 U875 ( .A1(n616), .A2(n615), .B(n614), .C(n613), .X(n617) );
  SEN_EO2_2 U876 ( .A1(n779), .A2(n520), .X(n782) );
  SEN_ND2_T_1 U877 ( .A1(n334), .A2(n519), .X(n520) );
  SEN_ND2_2 U878 ( .A1(n643), .A2(n642), .X(n644) );
  SEN_NR3_G_1 U879 ( .A1(n771), .A2(n770), .A3(n445), .X(n772) );
  SEN_NR2_1 U880 ( .A1(n671), .A2(n422), .X(n461) );
  SEN_ND2_G_1 U881 ( .A1(n806), .A2(n548), .X(n551) );
  SEN_ND2_G_1 U882 ( .A1(n462), .A2(n440), .X(n917) );
  SEN_INV_2 U883 ( .A(n433), .X(n696) );
  SEN_OAI21_G_1 U884 ( .A1(n884), .A2(n332), .B(n883), .X(Z[26]) );
  SEN_OAI211_1 U885 ( .A1(n839), .A2(n897), .B1(n838), .B2(n837), .X(Z[18]) );
  SEN_ND2_G_1 U886 ( .A1(n836), .A2(n906), .X(n837) );
  SEN_OAI211_1 U887 ( .A1(n846), .A2(n897), .B1(n845), .B2(n844), .X(Z[19]) );
  SEN_ND2_G_1 U888 ( .A1(n843), .A2(n906), .X(n844) );
  SEN_OAI211_1 U889 ( .A1(n332), .A2(n853), .B1(n852), .B2(n851), .X(Z[20]) );
  SEN_ND2_G_1 U890 ( .A1(n850), .A2(n906), .X(n851) );
  SEN_OAI211_1 U891 ( .A1(n332), .A2(n831), .B1(n830), .B2(n829), .X(Z[17]) );
  SEN_ND2_G_1 U892 ( .A1(n828), .A2(n333), .X(n829) );
  SEN_OAI211_1 U893 ( .A1(n782), .A2(n897), .B1(n781), .B2(n780), .X(Z[10]) );
  SEN_ND2_G_1 U894 ( .A1(n779), .A2(n333), .X(n780) );
  SEN_OAI211_1 U895 ( .A1(n809), .A2(n897), .B1(n808), .B2(n807), .X(Z[14]) );
  SEN_ND2_G_1 U896 ( .A1(n806), .A2(n906), .X(n807) );
  SEN_OAI211_1 U897 ( .A1(n737), .A2(n897), .B1(n736), .B2(n735), .X(Z[4]) );
  SEN_ND2_G_1 U898 ( .A1(n734), .A2(n333), .X(n735) );
  SEN_ND2_G_1 U899 ( .A1(n799), .A2(n906), .X(n800) );
  SEN_ND2_G_1 U900 ( .A1(n762), .A2(n917), .X(n767) );
  SEN_OAI211_1 U901 ( .A1(n722), .A2(n897), .B1(n721), .B2(n720), .X(Z[2]) );
  SEN_ND2_G_1 U902 ( .A1(n719), .A2(n333), .X(n720) );
  SEN_OAI211_1 U903 ( .A1(n789), .A2(n897), .B1(n788), .B2(n787), .X(Z[11]) );
  SEN_ND2_G_1 U904 ( .A1(n786), .A2(n906), .X(n787) );
  SEN_OAI211_1 U905 ( .A1(n860), .A2(n897), .B1(n859), .B2(n858), .X(Z[21]) );
  SEN_ND2_G_1 U906 ( .A1(n857), .A2(n333), .X(n858) );
  SEN_NR3_G_1 U907 ( .A1(n855), .A2(n854), .A3(n445), .X(n856) );
  SEN_OAI211_1 U908 ( .A1(n816), .A2(n897), .B1(n815), .B2(n814), .X(Z[15]) );
  SEN_ND2_G_1 U909 ( .A1(n813), .A2(n333), .X(n814) );
  SEN_NR3_G_1 U910 ( .A1(n741), .A2(n740), .A3(n445), .X(n742) );
  SEN_ND2_G_1 U911 ( .A1(n746), .A2(n917), .X(n751) );
  SEN_ND2_G_1 U912 ( .A1(n754), .A2(n917), .X(n759) );
  SEN_ND2_G_1 U913 ( .A1(n769), .A2(n917), .X(n774) );
  SEN_ND2_G_1 U914 ( .A1(n691), .A2(n705), .X(n693) );
  SEN_INV_S_1 U915 ( .A(n460), .X(n688) );
  SEN_ND2_G_1 U916 ( .A1(n675), .A2(n674), .X(n678) );
  SEN_OAI21_G_1 U917 ( .A1(n650), .A2(n874), .B(n649), .X(n651) );
  SEN_AOAI211_G_1 U918 ( .A1(n627), .A2(n630), .B(n633), .C(n625), .X(n626) );
  SEN_OAI21_G_1 U919 ( .A1(n608), .A2(n605), .B(n604), .X(n606) );
  SEN_ND2_G_1 U920 ( .A1(n603), .A2(n601), .X(n605) );
  SEN_ND2_G_1 U921 ( .A1(n573), .A2(n572), .X(n574) );
  SEN_ND2_G_1 U922 ( .A1(n573), .A2(n575), .X(n569) );
  SEN_OAI21_G_1 U923 ( .A1(n562), .A2(n551), .B(n550), .X(n552) );
  SEN_OAI21_G_1 U924 ( .A1(n537), .A2(n536), .B(n535), .X(n538) );
  SEN_OAI21_G_1 U925 ( .A1(n528), .A2(n511), .B(n510), .X(n517) );
  SEN_NR2_1 U926 ( .A1(n895), .A2(n894), .X(n667) );
  SEN_ND2_G_1 U927 ( .A1(n582), .A2(n581), .X(n583) );
  SEN_ND2_G_1 U928 ( .A1(n855), .A2(n854), .X(n581) );
  SEN_NR2_1 U929 ( .A1(n561), .A2(n560), .X(n549) );
  SEN_ND2_G_1 U930 ( .A1(n542), .A2(n541), .X(n493) );
  SEN_NR2_1 U931 ( .A1(n748), .A2(n747), .X(n485) );
  SEN_ND2_G_1 U932 ( .A1(n741), .A2(n740), .X(n512) );
  SEN_ND2_G_1 U933 ( .A1(n732), .A2(n731), .X(n535) );
  SEN_ND2_G_1 U934 ( .A1(n895), .A2(n894), .X(n662) );
  SEN_ND2_G_1 U935 ( .A1(n639), .A2(n640), .X(n663) );
  SEN_ND2_G_1 U936 ( .A1(n886), .A2(n885), .X(n634) );
  SEN_NR2_1 U937 ( .A1(n869), .A2(n868), .X(n648) );
  SEN_ND2_G_1 U938 ( .A1(n866), .A2(n865), .X(n593) );
  SEN_ND3_S_0P5 U939 ( .A1(n901), .A2(n900), .A3(n899), .X(n902) );
  SEN_ND3_S_0P5 U940 ( .A1(n886), .A2(n900), .A3(n885), .X(n887) );
  SEN_ND3_S_0P5 U941 ( .A1(n877), .A2(n876), .A3(n900), .X(n878) );
  SEN_ND3_S_0P5 U942 ( .A1(n708), .A2(n900), .A3(n707), .X(n709) );
  SEN_INV_S_1 U943 ( .A(n690), .X(n691) );
  SEN_INV_S_1 U944 ( .A(n647), .X(n650) );
  SEN_INV_S_1 U945 ( .A(n641), .X(n643) );
  SEN_INV_S_1 U946 ( .A(n818), .X(n637) );
  SEN_INV_S_1 U947 ( .A(n629), .X(n625) );
  SEN_INV_S_1 U948 ( .A(n876), .X(n619) );
  SEN_MUXI2_S_1 U949 ( .D0(n605), .D1(n600), .S(n609), .X(n607) );
  SEN_EN2_0P5 U950 ( .A1(n770), .A2(n771), .X(n775) );
  SEN_EN2_0P5 U951 ( .A1(n868), .A2(n869), .X(n870) );
  SEN_INV_S_1 U952 ( .A(n571), .X(n572) );
  SEN_EN2_0P5 U953 ( .A1(n832), .A2(n833), .X(n835) );
  SEN_INV_S_1 U954 ( .A(n561), .X(n797) );
  SEN_INV_S_1 U955 ( .A(n560), .X(n796) );
  SEN_INV_S_1 U956 ( .A(n575), .X(n557) );
  SEN_INV_S_1 U957 ( .A(n549), .X(n545) );
  SEN_INV_S_1 U958 ( .A(n542), .X(n804) );
  SEN_INV_S_1 U959 ( .A(n541), .X(n803) );
  SEN_EO2_S_0P5 U960 ( .A1(n786), .A2(n532), .X(n789) );
  SEN_INV_S_1 U961 ( .A(n526), .X(n527) );
  SEN_EO2_S_0P5 U962 ( .A1(n464), .A2(n694), .X(n525) );
  SEN_EO2_S_0P5 U963 ( .A1(n692), .A2(n689), .X(n694) );
  SEN_EO2_S_0P5 U964 ( .A1(n713), .A2(n524), .X(n715) );
  SEN_EN2_0P5 U965 ( .A1(n719), .A2(n521), .X(n722) );
  SEN_INV_S_1 U966 ( .A(n518), .X(n519) );
  SEN_AOI21_S_1 U967 ( .A1(n515), .A2(n514), .B(n513), .X(n516) );
  SEN_INV_S_1 U968 ( .A(n535), .X(n515) );
  SEN_INV_S_1 U969 ( .A(n502), .X(n503) );
  SEN_EN2_0P5 U970 ( .A1(n817), .A2(n818), .X(n820) );
  SEN_MUXI2_S_1 U971 ( .D0(n439), .D1(n436), .S(A[31]), .X(n920) );
  SEN_MUXI2_S_1 U972 ( .D0(n443), .D1(n441), .S(B[31]), .X(n921) );
  SEN_INV_S_1 U973 ( .A(n847), .X(n558) );
  SEN_INV_S_1 U974 ( .A(n848), .X(n559) );
  SEN_AOI22_1 U975 ( .A1(n825), .A2(n826), .B1(n818), .B2(n817), .X(n589) );
  SEN_MUXI2_S_1 U976 ( .D0(n437), .D1(n440), .S(n492), .X(n541) );
  SEN_MUXI2_S_1 U977 ( .D0(n437), .D1(n440), .S(n490), .X(n560) );
  SEN_MUXI2_S_1 U978 ( .D0(n439), .D1(n436), .S(A[28]), .X(n894) );
  SEN_MUXI2_S_1 U979 ( .D0(n443), .D1(n441), .S(B[28]), .X(n895) );
  SEN_MUXI2_S_1 U980 ( .D0(n338), .D1(n440), .S(n888), .X(n885) );
  SEN_MUXI2_S_1 U981 ( .D0(n338), .D1(n440), .S(n880), .X(n876) );
  SEN_MUXI2_S_1 U982 ( .D0(n439), .D1(n436), .S(A[25]), .X(n872) );
  SEN_MUXI2_S_1 U983 ( .D0(n443), .D1(n441), .S(B[25]), .X(n873) );
  SEN_MUXI2_S_1 U984 ( .D0(n439), .D1(n436), .S(A[24]), .X(n868) );
  SEN_INV_S_1 U985 ( .A(n855), .X(n591) );
  SEN_MUXI2_S_1 U986 ( .D0(n421), .D1(n440), .S(n904), .X(n899) );
  SEN_MUXI2_S_1 U987 ( .D0(n443), .D1(n441), .S(B[30]), .X(n912) );
  SEN_MUXI2_S_1 U988 ( .D0(n439), .D1(n436), .S(A[30]), .X(n911) );
  SEN_AO21B_1 U989 ( .A1(n909), .A2(n917), .B(n908), .X(Z[29]) );
  SEN_AO21B_1 U990 ( .A1(n893), .A2(n917), .B(n892), .X(Z[27]) );
endmodule

