
module Alu ( Z, A, B, INST, FLAGS );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  output [3:0] FLAGS;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062;

  SEN_INV_2 U416 ( .A(n362), .X(n364) );
  SEN_INV_2 U417 ( .A(n362), .X(n363) );
  SEN_ND2_G_1 U418 ( .A1(n540), .A2(A[8]), .X(n592) );
  SEN_ND2_G_1 U419 ( .A1(n701), .A2(n700), .X(n907) );
  SEN_ND2_G_1 U420 ( .A1(n623), .A2(n622), .X(n939) );
  SEN_ND2_G_1 U421 ( .A1(n536), .A2(n609), .X(n610) );
  SEN_INV_S_1 U422 ( .A(n985), .X(n978) );
  SEN_ND3_S_0P5 U423 ( .A1(n736), .A2(n779), .A3(n735), .X(n737) );
  SEN_ND2_G_1 U424 ( .A1(n533), .A2(n734), .X(n735) );
  SEN_NR2_1 U425 ( .A1(n738), .A2(n546), .X(n825) );
  SEN_ND3_S_0P5 U426 ( .A1(n755), .A2(n779), .A3(n754), .X(n756) );
  SEN_ND2_G_1 U427 ( .A1(n533), .A2(n753), .X(n754) );
  SEN_NR2_1 U428 ( .A1(n751), .A2(n546), .X(n861) );
  SEN_NR2_1 U429 ( .A1(n862), .A2(n861), .X(n820) );
  SEN_ND3_S_0P5 U430 ( .A1(n760), .A2(n779), .A3(n759), .X(n761) );
  SEN_ND2_G_1 U431 ( .A1(n533), .A2(n758), .X(n759) );
  SEN_INV_S_1 U432 ( .A(n793), .X(n782) );
  SEN_INV_S_1 U433 ( .A(n1057), .X(n552) );
  SEN_INV_S_1 U434 ( .A(n1010), .X(n1053) );
  SEN_EO2_G_2 U435 ( .A1(n917), .A2(n918), .X(n919) );
  SEN_NR2_1 U436 ( .A1(n851), .A2(n858), .X(n850) );
  SEN_EO2_2 U437 ( .A1(n916), .A2(n915), .X(n914) );
  SEN_INV_S_1 U438 ( .A(n914), .X(n496) );
  SEN_INV_2 U439 ( .A(n1036), .X(n548) );
  SEN_INV_S_1 U440 ( .A(n778), .X(n806) );
  SEN_INV_S_1 U441 ( .A(n1010), .X(n366) );
  SEN_EO2_S_0P5 U442 ( .A1(n805), .A2(n778), .X(n810) );
  SEN_INV_S_1 U443 ( .A(n552), .X(n551) );
  SEN_INV_2 U444 ( .A(n556), .X(n553) );
  SEN_EO2_S_0P5 U445 ( .A1(n792), .A2(n782), .X(n796) );
  SEN_NR2_1 U446 ( .A1(n806), .A2(n805), .X(n799) );
  SEN_INV_S_1 U447 ( .A(n796), .X(n788) );
  SEN_INV_S_1 U448 ( .A(n799), .X(n787) );
  SEN_INV_S_1 U449 ( .A(n552), .X(n550) );
  SEN_NR2_2 U450 ( .A1(n786), .A2(n790), .X(n1044) );
  SEN_INV_S_1 U451 ( .A(n548), .X(n549) );
  SEN_NR2_1 U452 ( .A1(n955), .A2(n954), .X(n676) );
  SEN_ND2_2 U453 ( .A1(n656), .A2(n840), .X(n661) );
  SEN_EO2_S_0P5 U454 ( .A1(n554), .A2(A[3]), .X(n616) );
  SEN_NR2_2 U455 ( .A1(n1031), .A2(n388), .X(n389) );
  SEN_EO2_S_0P5 U456 ( .A1(n554), .A2(A[14]), .X(n602) );
  SEN_EO2_S_0P5 U457 ( .A1(n555), .A2(A[15]), .X(n430) );
  SEN_OAI21_G_1 U458 ( .A1(n638), .A2(n553), .B(n789), .X(n1051) );
  SEN_NR2_1 U459 ( .A1(n534), .A2(A[0]), .X(n1047) );
  SEN_INV_S_1 U460 ( .A(n944), .X(n634) );
  SEN_ND3_T_2 U461 ( .A1(n592), .A2(n591), .A3(n590), .X(n999) );
  SEN_AOI21_S_1 U462 ( .A1(n533), .A2(n588), .B(n365), .X(n591) );
  SEN_INV_2 U463 ( .A(n654), .X(n472) );
  SEN_NR2_1 U464 ( .A1(n389), .A2(n935), .X(n469) );
  SEN_EO2_S_0P5 U465 ( .A1(n555), .A2(A[9]), .X(n568) );
  SEN_INV_2 U466 ( .A(n556), .X(n555) );
  SEN_ND2_2 U467 ( .A1(n789), .A2(n1050), .X(n791) );
  SEN_NR2_1 U468 ( .A1(n678), .A2(n546), .X(n986) );
  SEN_ND2_G_1 U469 ( .A1(n914), .A2(n908), .X(n909) );
  SEN_OAI22_1 U470 ( .A1(n905), .A2(n896), .B1(n901), .B2(n900), .X(n885) );
  SEN_NR2_1 U471 ( .A1(n905), .A2(n977), .X(n886) );
  SEN_ND3_S_0P5 U472 ( .A1(n744), .A2(n779), .A3(n743), .X(n745) );
  SEN_NR2_1 U473 ( .A1(n740), .A2(n546), .X(n871) );
  SEN_ND3_S_0P5 U474 ( .A1(n777), .A2(n776), .A3(n775), .X(n778) );
  SEN_EO2_S_0P5 U475 ( .A1(n553), .A2(A[30]), .X(n774) );
  SEN_INV_S_1 U476 ( .A(Z[29]), .X(n502) );
  SEN_EO2_S_0P5 U477 ( .A1(n358), .A2(n1007), .X(n1008) );
  SEN_INV_S_1 U478 ( .A(n998), .X(n997) );
  SEN_EO2_S_0P5 U479 ( .A1(n996), .A2(n989), .X(n990) );
  SEN_OAI21_G_1 U480 ( .A1(n989), .A2(n996), .B(n930), .X(n441) );
  SEN_NR2_1 U481 ( .A1(n933), .A2(n1036), .X(n439) );
  SEN_AN3B_1 U482 ( .B1(n932), .B2(n1010), .A(n931), .X(n440) );
  SEN_NR2_T_1 U483 ( .A1(n584), .A2(n545), .X(n917) );
  SEN_EO2_S_0P5 U484 ( .A1(n919), .A2(n419), .X(n426) );
  SEN_INV_S_1 U485 ( .A(n906), .X(n988) );
  SEN_EO2_S_0P5 U486 ( .A1(n978), .A2(n414), .X(n979) );
  SEN_EO2_1 U487 ( .A1(n980), .A2(n981), .X(n985) );
  SEN_NR2_1 U488 ( .A1(n527), .A2(n549), .X(n446) );
  SEN_EO2_1 U489 ( .A1(n972), .A2(n973), .X(n977) );
  SEN_EO2_1 U490 ( .A1(n889), .A2(n890), .X(n892) );
  SEN_EO2_S_0P5 U491 ( .A1(n871), .A2(n872), .X(n874) );
  SEN_INV_S_1 U492 ( .A(n860), .X(n866) );
  SEN_ND3_S_0P5 U493 ( .A1(n768), .A2(n779), .A3(n767), .X(n769) );
  SEN_EO2_S_0P5 U494 ( .A1(n553), .A2(A[29]), .X(n765) );
  SEN_AO21B_1 U495 ( .A1(n785), .A2(n788), .B(n784), .X(FLAGS[1]) );
  SEN_ND2_G_1 U496 ( .A1(n1041), .A2(n548), .X(n1042) );
  SEN_EO2_S_0P5 U497 ( .A1(n525), .A2(n1029), .X(n1030) );
  SEN_OAI211_1 U498 ( .A1(n1036), .A2(n858), .B1(n857), .B2(n856), .X(Z[14])
         );
  SEN_ND2_G_1 U499 ( .A1(n852), .A2(n367), .X(n857) );
  SEN_OAOI211_G_1 U500 ( .A1(n850), .A2(n847), .B(n846), .C(n845), .X(n848) );
  SEN_OAI21_G_1 U501 ( .A1(n490), .A2(n1044), .B(n491), .X(Z[18]) );
  SEN_EO2_1 U502 ( .A1(n496), .A2(n497), .X(n490) );
  SEN_OAI211_1 U503 ( .A1(n399), .A2(n1044), .B1(n400), .B2(n401), .X(Z[25])
         );
  SEN_ND2_G_1 U504 ( .A1(n868), .A2(n548), .X(n401) );
  SEN_OAI21_G_1 U505 ( .A1(n403), .A2(n1044), .B(n404), .X(Z[28]) );
  SEN_AOI21B_1 U506 ( .A1(n823), .A2(n548), .B(n405), .X(n404) );
  SEN_EO2_S_0P5 U507 ( .A1(n823), .A2(n408), .X(n403) );
  SEN_AOI21B_1 U508 ( .A1(n859), .A2(n860), .B(n409), .X(n408) );
  SEN_ND2_G_1 U509 ( .A1(n800), .A2(n516), .X(Z[31]) );
  SEN_OR2_1 U510 ( .A1(n802), .A2(n801), .X(n516) );
  SEN_OAOI211_G_1 U511 ( .A1(n802), .A2(n799), .B(n798), .C(n797), .X(n800) );
  SEN_ND3_S_0P5 U512 ( .A1(n788), .A2(n1058), .A3(n787), .X(n801) );
  SEN_ND2B_1 U513 ( .A(n972), .B(n973), .X(n896) );
  SEN_INV_0P5 U514 ( .A(n541), .X(n348) );
  SEN_NR2_0P5 U515 ( .A1(n543), .A2(B[31]), .X(n349) );
  SEN_AOI211_0P5 U516 ( .A1(B[31]), .A2(n348), .B1(n547), .B2(n349), .X(n792)
         );
  SEN_NR3B_1 U517 ( .A(n1048), .B1(n364), .B2(n1047), .X(n1055) );
  SEN_ND2B_1 U518 ( .A(n991), .B(n992), .X(n930) );
  SEN_INV_0P5 U519 ( .A(n541), .X(n350) );
  SEN_NR2_0P5 U520 ( .A1(n361), .A2(B[28]), .X(n351) );
  SEN_AOI211_0P5 U521 ( .A1(B[28]), .A2(n350), .B1(n546), .B2(n351), .X(n821)
         );
  SEN_ND2B_1 U522 ( .A(n802), .B(n787), .X(n785) );
  SEN_ND2B_1 U523 ( .A(n792), .B(n782), .X(n784) );
  SEN_OR3_1 U524 ( .A1(n789), .A2(n529), .A3(n790), .X(n1036) );
  SEN_OAI21_0P5 U525 ( .A1(A[19]), .A2(B[19]), .B(n551), .X(n352) );
  SEN_OAI31_0P5 U526 ( .A1(n912), .A2(n911), .A3(n366), .B(n352), .X(n447) );
  SEN_EO2_S_0P5 U527 ( .A1(n1054), .A2(n1055), .X(n1062) );
  SEN_AN3_0P5 U528 ( .A1(n624), .A2(n1011), .A3(n1010), .X(n1012) );
  SEN_EN2_S_2 U529 ( .A1(n955), .A2(n954), .X(n959) );
  SEN_INV_0P5 U530 ( .A(n541), .X(n353) );
  SEN_NR2_0P5 U531 ( .A1(n361), .A2(B[29]), .X(n354) );
  SEN_AOI211_0P5 U532 ( .A1(B[29]), .A2(n353), .B1(n547), .B2(n354), .X(n814)
         );
  SEN_ND2_0P5 U533 ( .A1(n1050), .A2(n1051), .X(n355) );
  SEN_OAI211_0P5 U534 ( .A1(n1050), .A2(n1049), .B1(n355), .B2(n1052), .X(
        n1061) );
  SEN_ND3B_0P5 U535 ( .A(n842), .B1(n373), .B2(n1010), .X(n843) );
  SEN_EO2_S_0P5 U536 ( .A1(n862), .A2(n861), .X(n860) );
  SEN_INV_0P5 U537 ( .A(n541), .X(n356) );
  SEN_NR2_0P5 U538 ( .A1(n543), .A2(B[30]), .X(n357) );
  SEN_AOI211_0P5 U539 ( .A1(B[30]), .A2(n356), .B1(n547), .B2(n357), .X(n805)
         );
  SEN_INV_5 U540 ( .A(n421), .X(n360) );
  SEN_ND2_T_5 U541 ( .A1(n1037), .A2(n1041), .X(n937) );
  SEN_AOI22_2 U542 ( .A1(n642), .A2(n1048), .B1(n1054), .B2(n641), .X(n1037)
         );
  SEN_OAI21_G_2 U543 ( .A1(n1007), .A2(n358), .B(n942), .X(n962) );
  SEN_NR2_2 U544 ( .A1(n643), .A2(n545), .X(n1038) );
  SEN_INV_4 U545 ( .A(n556), .X(n554) );
  SEN_OAI211_2 U546 ( .A1(n1036), .A2(n358), .B1(n1014), .B2(n1013), .X(Z[5])
         );
  SEN_OAI211_2 U547 ( .A1(n1062), .A2(n1061), .B1(n1060), .B2(n1059), .X(Z[0])
         );
  SEN_INV_S_1 U548 ( .A(n1044), .X(n367) );
  SEN_EO2_S_0P5 U549 ( .A1(n1009), .A2(n1011), .X(n358) );
  SEN_INV_2 U550 ( .A(A[31]), .X(n556) );
  SEN_EN2_0P5 U551 ( .A1(n933), .A2(n441), .X(n442) );
  SEN_INV_3 U552 ( .A(n506), .X(n504) );
  SEN_OAI21_G_1 U553 ( .A1(n785), .A2(n784), .B(n783), .X(FLAGS[0]) );
  SEN_NR2_T_1P5 U554 ( .A1(Z[28]), .A2(Z[14]), .X(n507) );
  SEN_OAI31_1 U555 ( .A1(n850), .A2(n374), .A3(n849), .B(n848), .X(Z[15]) );
  SEN_OAI21_T_2 U556 ( .A1(n448), .A2(n444), .B(n449), .X(Z[24]) );
  SEN_ND2_2 U557 ( .A1(n830), .A2(n1058), .X(n835) );
  SEN_AOI21_S_2 U558 ( .A1(n887), .A2(n886), .B(n885), .X(n888) );
  SEN_ND2_3 U559 ( .A1(n411), .A2(n827), .X(n418) );
  SEN_NR2_T_2 U560 ( .A1(n410), .A2(n929), .X(n989) );
  SEN_OAI21_4 U561 ( .A1(n410), .A2(n412), .B(n413), .X(n411) );
  SEN_INV_0P65 U562 ( .A(Z[4]), .X(n499) );
  SEN_AOI21_S_2 U563 ( .A1(n880), .A2(n881), .B(n884), .X(n397) );
  SEN_NR2_0P65 U564 ( .A1(n788), .A2(n1044), .X(n798) );
  SEN_NR2_G_0P8 U565 ( .A1(n841), .A2(n1044), .X(n846) );
  SEN_INV_1 U566 ( .A(n938), .X(n1028) );
  SEN_OAOI211_G_1 U567 ( .A1(B[11]), .A2(A[11]), .B(n550), .C(n923), .X(n926)
         );
  SEN_OAOI211_G_1 U568 ( .A1(A[3]), .A2(B[3]), .B(n550), .C(n458), .X(n457) );
  SEN_OAOI211_G_1 U569 ( .A1(B[20]), .A2(A[20]), .B(n550), .C(n956), .X(n957)
         );
  SEN_ND2_2 U570 ( .A1(n747), .A2(n746), .X(n748) );
  SEN_INV_2 U571 ( .A(n905), .X(n898) );
  SEN_OAOI211_G_1 U572 ( .A1(A[27]), .A2(B[27]), .B(n551), .C(n863), .X(n864)
         );
  SEN_INV_1 U573 ( .A(n625), .X(n526) );
  SEN_OAI21_G_2 U574 ( .A1(n868), .A2(n867), .B(n874), .X(n749) );
  SEN_ND2_3 U575 ( .A1(n918), .A2(n585), .X(n829) );
  SEN_OAOI211_G_1 U576 ( .A1(B[26]), .A2(A[26]), .B(n551), .C(n873), .X(n876)
         );
  SEN_OAOI211_G_1 U577 ( .A1(A[23]), .A2(B[23]), .B(n551), .C(n891), .X(n894)
         );
  SEN_OAOI211_G_1 U578 ( .A1(B[25]), .A2(A[25]), .B(n551), .C(n402), .X(n400)
         );
  SEN_NR2_G_1 U579 ( .A1(n884), .A2(n549), .X(n451) );
  SEN_INV_S_1 U580 ( .A(n828), .X(n460) );
  SEN_NR2_G_1 U581 ( .A1(n914), .A2(n549), .X(n492) );
  SEN_OAOI211_G_1 U582 ( .A1(B[14]), .A2(A[14]), .B(n551), .C(n855), .X(n856)
         );
  SEN_EO2_3 U583 ( .A1(n842), .A2(n373), .X(n374) );
  SEN_NR3_T_0P65 U584 ( .A1(n793), .A2(n792), .A3(n366), .X(n794) );
  SEN_INV_1 U585 ( .A(n821), .X(n762) );
  SEN_INV_1 U586 ( .A(n815), .X(n771) );
  SEN_EO2_4 U587 ( .A1(n1026), .A2(n1027), .X(n938) );
  SEN_INV_1 U588 ( .A(n871), .X(n747) );
  SEN_NR2_1 U589 ( .A1(n821), .A2(n366), .X(n406) );
  SEN_EO2_8 U590 ( .A1(n900), .A2(n718), .X(n905) );
  SEN_NR2_G_2 U591 ( .A1(n883), .A2(n882), .X(n824) );
  SEN_NR2_G_1 U592 ( .A1(n826), .A2(n825), .X(n867) );
  SEN_ND2_S_0P5 U593 ( .A1(n915), .A2(n1010), .X(n494) );
  SEN_NR2_T_2 U594 ( .A1(n600), .A2(n545), .X(n831) );
  SEN_INV_2 U595 ( .A(n622), .X(n1026) );
  SEN_NR2_T_3 U596 ( .A1(n455), .A2(n545), .X(n388) );
  SEN_NR2_S_3 U597 ( .A1(n684), .A2(n546), .X(n980) );
  SEN_NR2_G_2 U598 ( .A1(n727), .A2(n546), .X(n882) );
  SEN_NR2_S_3 U599 ( .A1(n706), .A2(n546), .X(n900) );
  SEN_ND3_T_2 U600 ( .A1(n672), .A2(n779), .A3(n671), .X(n673) );
  SEN_INV_16 U601 ( .A(n360), .X(n545) );
  SEN_ND3_T_2 U602 ( .A1(n583), .A2(n582), .A3(n581), .X(n918) );
  SEN_ND2_2 U603 ( .A1(n372), .A2(A[6]), .X(n612) );
  SEN_INV_8 U604 ( .A(n363), .X(n779) );
  SEN_INV_1 U605 ( .A(n640), .X(n641) );
  SEN_OAI21_G_1 U606 ( .A1(B[6]), .A2(A[6]), .B(n551), .X(n947) );
  SEN_INV_6 U607 ( .A(n1046), .X(n362) );
  SEN_EO2_2 U608 ( .A1(A[5]), .A2(n554), .X(n464) );
  SEN_EO2_S_1 U609 ( .A1(n553), .A2(A[23]), .X(n720) );
  SEN_INV_1 U610 ( .A(A[26]), .X(n742) );
  SEN_INV_1 U611 ( .A(A[20]), .X(n670) );
  SEN_ND4_S_6 U612 ( .A1(n504), .A2(n502), .A3(n501), .A4(n507), .X(n505) );
  SEN_ND2_T_2 U613 ( .A1(n809), .A2(n517), .X(Z[30]) );
  SEN_ND2_2 U614 ( .A1(n804), .A2(n367), .X(n809) );
  SEN_OAI211_2 U615 ( .A1(n819), .A2(n549), .B1(n818), .B2(n817), .X(Z[29]) );
  SEN_NR2_T_4 U616 ( .A1(n803), .A2(n810), .X(n802) );
  SEN_ND2_T_2 U617 ( .A1(n904), .A2(n519), .X(Z[22]) );
  SEN_EO2_2 U618 ( .A1(n892), .A2(n888), .X(n895) );
  SEN_ND2_2 U619 ( .A1(n899), .A2(n367), .X(n904) );
  SEN_ND2_2 U620 ( .A1(n953), .A2(n1058), .X(n958) );
  SEN_AOAI211_G_3 U621 ( .A1(n937), .A2(n469), .B(n470), .C(n471), .X(n468) );
  SEN_AOI22_T_3 U622 ( .A1(n885), .A2(n892), .B1(n726), .B2(n725), .X(n880) );
  SEN_AN2_1 U623 ( .A1(n978), .A2(n909), .X(n415) );
  SEN_ND2_G_0P65 U624 ( .A1(n840), .A2(n367), .X(n849) );
  SEN_INV_1 U625 ( .A(n928), .X(n929) );
  SEN_ND3_T_2 U626 ( .A1(n460), .A2(n827), .A3(n829), .X(n657) );
  SEN_OAOI211_G_1 U627 ( .A1(A[2]), .A2(B[2]), .B(n550), .C(n1032), .X(n1033)
         );
  SEN_OAOI211_1 U628 ( .A1(A[21]), .A2(B[21]), .B(n550), .C(n974), .X(n975) );
  SEN_AOAI211_1 U629 ( .A1(n1058), .A2(n1061), .B(n548), .C(n1062), .X(n1059)
         );
  SEN_OAOI211_G_1 U630 ( .A1(A[1]), .A2(B[1]), .B(n550), .C(n1040), .X(n1043)
         );
  SEN_AOI22_T_1 U631 ( .A1(n823), .A2(n820), .B1(n359), .B2(n762), .X(n763) );
  SEN_OAOI211_1 U632 ( .A1(B[12]), .A2(A[12]), .B(n550), .C(n425), .X(n424) );
  SEN_OAOI211_1 U633 ( .A1(A[9]), .A2(B[9]), .B(n550), .C(n993), .X(n994) );
  SEN_OAOI211_1 U634 ( .A1(A[17]), .A2(B[17]), .B(n550), .C(n982), .X(n983) );
  SEN_OR2_1 U635 ( .A1(n985), .A2(n549), .X(n521) );
  SEN_NR2_G_1 U636 ( .A1(n950), .A2(n676), .X(n698) );
  SEN_AOI22_1 U637 ( .A1(n359), .A2(n406), .B1(n551), .B2(n407), .X(n405) );
  SEN_NR3_1 U638 ( .A1(n1055), .A2(n1054), .A3(n1053), .X(n1056) );
  SEN_INV_1 U639 ( .A(n889), .X(n725) );
  SEN_INV_1 U640 ( .A(n890), .X(n726) );
  SEN_INV_1 U641 ( .A(n980), .X(n696) );
  SEN_INV_2 U642 ( .A(n911), .X(n523) );
  SEN_EO2_G_2 U643 ( .A1(n814), .A2(n815), .X(n812) );
  SEN_INV_2 U644 ( .A(n814), .X(n770) );
  SEN_OAI21_G_1 U645 ( .A1(n494), .A2(n916), .B(n495), .X(n493) );
  SEN_NR3_1 U646 ( .A1(n955), .A2(n954), .A3(n366), .X(n956) );
  SEN_NR3_T_0P65 U647 ( .A1(n862), .A2(n861), .A3(n366), .X(n863) );
  SEN_INV_0P8 U648 ( .A(n872), .X(n746) );
  SEN_NR3_T_0P65 U649 ( .A1(n815), .A2(n814), .A3(n366), .X(n816) );
  SEN_NR2_G_2 U650 ( .A1(n719), .A2(n546), .X(n889) );
  SEN_NR2_T_2 U651 ( .A1(n572), .A2(n545), .X(n991) );
  SEN_NR2_T_2 U652 ( .A1(n594), .A2(n545), .X(n842) );
  SEN_NR2_T_3 U653 ( .A1(n587), .A2(n545), .X(n1001) );
  SEN_NR2_T_2 U654 ( .A1(n668), .A2(n546), .X(n911) );
  SEN_NR2_T_2 U655 ( .A1(n712), .A2(n546), .X(n972) );
  SEN_NR2_S_4 U656 ( .A1(n674), .A2(n546), .X(n954) );
  SEN_ND3_T_2 U657 ( .A1(n711), .A2(n710), .A3(n709), .X(n718) );
  SEN_ND3_T_2 U658 ( .A1(n732), .A2(n731), .A3(n730), .X(n739) );
  SEN_OAI21_G_1 U659 ( .A1(A[8]), .A2(B[8]), .B(n550), .X(n1000) );
  SEN_OAI21_G_1 U660 ( .A1(A[4]), .A2(B[4]), .B(n550), .X(n1018) );
  SEN_OAI21_G_1 U661 ( .A1(B[18]), .A2(A[18]), .B(n551), .X(n495) );
  SEN_INV_1 U662 ( .A(n367), .X(n444) );
  SEN_INV_3 U663 ( .A(n362), .X(n365) );
  SEN_ND2_T_6 U664 ( .A1(n376), .A2(n377), .X(n371) );
  SEN_EO2_1 U665 ( .A1(n555), .A2(A[12]), .X(n580) );
  SEN_NR2_T_2 U666 ( .A1(n1049), .A2(n420), .X(n421) );
  SEN_INV_0P5 U667 ( .A(n1044), .X(n1058) );
  SEN_INV_5 U668 ( .A(n529), .X(n1050) );
  SEN_INV_2 U669 ( .A(n531), .X(n638) );
  SEN_INV_0P8 U670 ( .A(A[17]), .X(n685) );
  SEN_INV_1 U671 ( .A(A[5]), .X(n465) );
  SEN_INV_0P8 U672 ( .A(A[21]), .X(n713) );
  SEN_INV_1 U673 ( .A(A[4]), .X(n384) );
  SEN_INV_0P8 U674 ( .A(A[14]), .X(n601) );
  SEN_INV_0P8 U675 ( .A(A[12]), .X(n579) );
  SEN_NR3_T_2 U676 ( .A1(Z[31]), .A2(n505), .A3(Z[30]), .X(FLAGS[2]) );
  SEN_INV_1 U677 ( .A(Z[15]), .X(n501) );
  SEN_OR4B_2 U678 ( .B1(Z[18]), .B2(Z[10]), .B3(Z[11]), .A(n511), .X(n510) );
  SEN_ND2_2 U679 ( .A1(n813), .A2(n1058), .X(n818) );
  SEN_OAI211_2 U680 ( .A1(n1036), .A2(n836), .B1(n835), .B2(n834), .X(Z[13])
         );
  SEN_INV_S_2 U681 ( .A(n394), .X(n869) );
  SEN_ND2_T_2 U682 ( .A1(n764), .A2(n763), .X(n811) );
  SEN_ND3_T_2 U683 ( .A1(n976), .A2(n975), .A3(n520), .X(Z[21]) );
  SEN_NR2_S_4 U684 ( .A1(n398), .A2(n824), .X(n394) );
  SEN_ND3_T_2 U685 ( .A1(n984), .A2(n983), .A3(n521), .X(Z[17]) );
  SEN_NR2B_V1_2 U686 ( .A(n500), .B(Z[16]), .X(n416) );
  SEN_AOI21_G_2 U687 ( .A1(n839), .A2(n838), .B(n837), .X(n851) );
  SEN_OAI211_2 U688 ( .A1(n927), .A2(n1044), .B1(n926), .B2(n925), .X(Z[11])
         );
  SEN_OAI21_G_2 U689 ( .A1(n970), .A2(n977), .B(n896), .X(n897) );
  SEN_INV_S_2 U690 ( .A(n393), .X(n398) );
  SEN_ND2_4 U691 ( .A1(n467), .A2(n468), .X(n390) );
  SEN_OAI21_0P75 U692 ( .A1(n1024), .A2(n1044), .B(n1023), .X(Z[4]) );
  SEN_NR2_S_4 U693 ( .A1(n472), .A2(n655), .X(n471) );
  SEN_NR2_G_2 U694 ( .A1(n446), .A2(n447), .X(n445) );
  SEN_NR2_G_2 U695 ( .A1(n481), .A2(n661), .X(n479) );
  SEN_OAOI211_1 U696 ( .A1(B[5]), .A2(A[5]), .B(n550), .C(n1012), .X(n1013) );
  SEN_INV_1 U697 ( .A(n829), .X(n607) );
  SEN_OR2_1 U698 ( .A1(n988), .A2(n549), .X(n417) );
  SEN_INV_1 U699 ( .A(n699), .X(n702) );
  SEN_AOI211_G_2 U700 ( .A1(n551), .A2(n450), .B1(n451), .B2(n452), .X(n449)
         );
  SEN_INV_1 U701 ( .A(n913), .X(n498) );
  SEN_ND2_3 U702 ( .A1(n942), .A2(n940), .X(n378) );
  SEN_NR2_G_1 U703 ( .A1(n492), .A2(n493), .X(n491) );
  SEN_AOI211_3 U704 ( .A1(n998), .A2(n928), .B1(n933), .B2(n996), .X(n481) );
  SEN_AOI211_G_2 U705 ( .A1(n550), .A2(n438), .B1(n439), .B2(n440), .X(n437)
         );
  SEN_NR2_G_1 U706 ( .A1(n1004), .A2(n1003), .X(n1005) );
  SEN_ND2_2 U707 ( .A1(n886), .A2(n892), .X(n881) );
  SEN_INV_1 U708 ( .A(n812), .X(n819) );
  SEN_INV_1 U709 ( .A(n660), .X(n487) );
  SEN_OAOI211_1 U710 ( .A1(n553), .A2(B[31]), .B(n550), .C(n794), .X(n795) );
  SEN_INV_1 U711 ( .A(n820), .X(n409) );
  SEN_OAOI211_1 U712 ( .A1(B[30]), .A2(A[30]), .B(n551), .C(n807), .X(n808) );
  SEN_NR2_G_1 U713 ( .A1(n867), .A2(n824), .X(n750) );
  SEN_OR2_1 U714 ( .A1(n977), .A2(n549), .X(n520) );
  SEN_NR2_G_2 U715 ( .A1(n466), .A2(n389), .X(n470) );
  SEN_ND2_2 U716 ( .A1(n874), .A2(n548), .X(n875) );
  SEN_INV_1 U717 ( .A(n676), .X(n677) );
  SEN_OAOI211_1 U718 ( .A1(A[22]), .A2(B[22]), .B(n551), .C(n902), .X(n903) );
  SEN_INV_4 U719 ( .A(n847), .X(n840) );
  SEN_ND2_2 U720 ( .A1(n892), .A2(n548), .X(n893) );
  SEN_OAOI211_1 U721 ( .A1(A[29]), .A2(B[29]), .B(n551), .C(n816), .X(n817) );
  SEN_OAOI211_1 U722 ( .A1(B[13]), .A2(A[13]), .B(n551), .C(n833), .X(n834) );
  SEN_INV_1 U723 ( .A(n838), .X(n836) );
  SEN_OAOI211_1 U724 ( .A1(A[16]), .A2(B[16]), .B(n550), .C(n435), .X(n434) );
  SEN_INV_1 U725 ( .A(n525), .X(n1035) );
  SEN_INV_1 U726 ( .A(n924), .X(n920) );
  SEN_OAOI211_1 U727 ( .A1(A[0]), .A2(B[0]), .B(n551), .C(n1056), .X(n1060) );
  SEN_EO2_4 U728 ( .A1(n1038), .A2(n1039), .X(n1041) );
  SEN_AN2_1 U729 ( .A1(n947), .A2(n946), .X(n522) );
  SEN_NR3_1 U730 ( .A1(n826), .A2(n825), .A3(n366), .X(n402) );
  SEN_EO2_2 U731 ( .A1(n388), .A2(n1031), .X(n466) );
  SEN_EO2_2 U732 ( .A1(n821), .A2(n822), .X(n823) );
  SEN_NR2_T_2 U733 ( .A1(n922), .A2(n921), .X(n828) );
  SEN_INV_1 U734 ( .A(n931), .X(n586) );
  SEN_NR3_1 U735 ( .A1(n883), .A2(n882), .A3(n366), .X(n452) );
  SEN_NR3_1 U736 ( .A1(n806), .A2(n805), .A3(n366), .X(n807) );
  SEN_NR3_1 U737 ( .A1(n832), .A2(n831), .A3(n366), .X(n833) );
  SEN_NR2_G_3 U738 ( .A1(n832), .A2(n831), .X(n837) );
  SEN_INV_1 U739 ( .A(n986), .X(n701) );
  SEN_INV_1 U740 ( .A(n916), .X(n697) );
  SEN_INV_1 U741 ( .A(n987), .X(n700) );
  SEN_EO2_2 U742 ( .A1(n882), .A2(n739), .X(n884) );
  SEN_NR3_1 U743 ( .A1(n890), .A2(n889), .A3(n366), .X(n891) );
  SEN_NR3_1 U744 ( .A1(n922), .A2(n921), .A3(n1053), .X(n923) );
  SEN_EO2_2 U745 ( .A1(n825), .A2(n826), .X(n868) );
  SEN_NR2_T_2 U746 ( .A1(n432), .A2(n842), .X(n660) );
  SEN_NR3_1 U747 ( .A1(n987), .A2(n986), .A3(n1053), .X(n435) );
  SEN_NR3_1 U748 ( .A1(n872), .A2(n871), .A3(n366), .X(n873) );
  SEN_NR3_1 U749 ( .A1(n901), .A2(n900), .A3(n1053), .X(n902) );
  SEN_INV_1 U750 ( .A(n718), .X(n901) );
  SEN_INV_1 U751 ( .A(n822), .X(n359) );
  SEN_INV_1 U752 ( .A(n739), .X(n883) );
  SEN_EN2_S_3 U753 ( .A1(n965), .A2(n966), .X(n969) );
  SEN_ND3_1 U754 ( .A1(n723), .A2(n779), .A3(n722), .X(n724) );
  SEN_ND3_T_2 U755 ( .A1(n717), .A2(n716), .A3(n715), .X(n973) );
  SEN_INV_6 U756 ( .A(n534), .X(n533) );
  SEN_INV_10 U757 ( .A(n544), .X(n361) );
  SEN_OAI21_S_0P5 U758 ( .A1(B[15]), .A2(A[15]), .B(n1057), .X(n844) );
  SEN_EO2_1 U759 ( .A1(n553), .A2(A[24]), .X(n729) );
  SEN_ND2_3 U760 ( .A1(n786), .A2(n557), .X(n781) );
  SEN_INV_1 U761 ( .A(A[2]), .X(n650) );
  SEN_OR2_1 U762 ( .A1(A[28]), .A2(B[28]), .X(n407) );
  SEN_INV_1 U763 ( .A(A[27]), .X(n753) );
  SEN_INV_0P8 U764 ( .A(A[30]), .X(n772) );
  SEN_OR2_1 U765 ( .A1(A[24]), .A2(B[24]), .X(n450) );
  SEN_INV_1 U766 ( .A(A[1]), .X(n645) );
  SEN_INV_0P8 U767 ( .A(A[19]), .X(n664) );
  SEN_INV_0P65 U768 ( .A(A[22]), .X(n707) );
  SEN_INV_1 U769 ( .A(A[11]), .X(n574) );
  SEN_INV_0P8 U770 ( .A(A[10]), .X(n561) );
  SEN_INV_0P8 U771 ( .A(A[8]), .X(n588) );
  SEN_INV_0P65 U772 ( .A(A[7]), .X(n627) );
  SEN_OR2_1 U773 ( .A1(A[10]), .A2(B[10]), .X(n438) );
  SEN_INV_1 U774 ( .A(A[28]), .X(n758) );
  SEN_INV_1 U775 ( .A(A[23]), .X(n721) );
  SEN_INV_1 U776 ( .A(A[13]), .X(n596) );
  SEN_INV_0P8 U777 ( .A(A[9]), .X(n567) );
  SEN_INV_1 U778 ( .A(A[16]), .X(n680) );
  SEN_INV_0P8 U779 ( .A(A[24]), .X(n728) );
  SEN_INV_0P65 U780 ( .A(A[18]), .X(n691) );
  SEN_INV_1 U781 ( .A(A[29]), .X(n766) );
  SEN_INV_0P8 U782 ( .A(A[15]), .X(n431) );
  SEN_INV_1 U783 ( .A(A[25]), .X(n734) );
  SEN_INV_0P8 U784 ( .A(A[3]), .X(n615) );
  SEN_INV_1 U785 ( .A(B[3]), .X(n620) );
  SEN_INV_1 U786 ( .A(B[6]), .X(n613) );
  SEN_INV_0P8 U787 ( .A(A[6]), .X(n608) );
  SEN_INV_1 U788 ( .A(B[7]), .X(n632) );
  SEN_MUXI2_S_3 U789 ( .D0(n542), .D1(n544), .S(n613), .X(n614) );
  SEN_INV_6 U790 ( .A(n781), .X(n544) );
  SEN_NR2_T_3 U791 ( .A1(n422), .A2(n545), .X(n1009) );
  SEN_MUXI2_S_2 U792 ( .D0(n361), .D1(n541), .S(B[20]), .X(n674) );
  SEN_MUXI2_S_2 U793 ( .D0(n543), .D1(n387), .S(B[2]), .X(n455) );
  SEN_ND3_T_2 U794 ( .A1(n612), .A2(n611), .A3(n610), .X(n945) );
  SEN_AOAI211_G_4 U795 ( .A1(n393), .A2(n750), .B(n749), .C(n748), .X(n859) );
  SEN_AOI21_2 U796 ( .A1(n532), .A2(n465), .B(n364), .X(n462) );
  SEN_OAI211_2 U797 ( .A1(n1036), .A2(n969), .B1(n968), .B2(n967), .X(Z[7]) );
  SEN_EO2_1 U798 ( .A1(n969), .A2(n963), .X(n964) );
  SEN_AOI21_S_1 U799 ( .A1(n532), .A2(n608), .B(n364), .X(n611) );
  SEN_NR3_G_1 U800 ( .A1(n1031), .A2(n388), .A3(n1053), .X(n1032) );
  SEN_NR2_T_1P5 U801 ( .A1(Z[24]), .A2(Z[19]), .X(n368) );
  SEN_NR3_T_3 U802 ( .A1(Z[23]), .A2(Z[12]), .A3(n369), .X(n514) );
  SEN_INV_2 U803 ( .A(n368), .X(n369) );
  SEN_OAI211_2 U804 ( .A1(n549), .A2(n919), .B1(n423), .B2(n424), .X(Z[12]) );
  SEN_ND3_T_2 U805 ( .A1(n514), .A2(n515), .A3(n503), .X(n508) );
  SEN_OAI211_3 U806 ( .A1(n895), .A2(n1044), .B1(n894), .B2(n893), .X(Z[23])
         );
  SEN_OAI21_3 U807 ( .A1(n391), .A2(n988), .B(n907), .X(n414) );
  SEN_EO2_2 U808 ( .A1(n874), .A2(n870), .X(n877) );
  SEN_INV_2 U809 ( .A(n373), .X(n432) );
  SEN_ND3_T_2 U810 ( .A1(n427), .A2(n428), .A3(n429), .X(n373) );
  SEN_BUF_6 U811 ( .A(INST[3]), .X(n370) );
  SEN_ND3_T_0P8 U812 ( .A1(n530), .A2(n531), .A3(n370), .X(n375) );
  SEN_ND2_4 U813 ( .A1(n531), .A2(n370), .X(n557) );
  SEN_INV_8 U814 ( .A(n370), .X(n1052) );
  SEN_ND2_T_4 U815 ( .A1(n370), .A2(n530), .X(n560) );
  SEN_ND2B_1 U816 ( .A(n531), .B(n370), .X(n790) );
  SEN_AOI21_S_1 U817 ( .A1(n1051), .A2(n1050), .B(n370), .X(n640) );
  SEN_INV_10 U818 ( .A(n371), .X(n372) );
  SEN_INV_4 U819 ( .A(n371), .X(n540) );
  SEN_INV_6 U820 ( .A(n371), .X(n539) );
  SEN_ND2_G_1 U821 ( .A1(n372), .A2(A[15]), .X(n427) );
  SEN_ND2_4 U822 ( .A1(n372), .A2(A[5]), .X(n461) );
  SEN_ND2_T_1P5 U823 ( .A1(n372), .A2(A[7]), .X(n631) );
  SEN_ND2_G_4 U824 ( .A1(n372), .A2(A[3]), .X(n619) );
  SEN_AOI21_T_2 U825 ( .A1(n372), .A2(A[20]), .B(n673), .X(n955) );
  SEN_ND2_G_1 U826 ( .A1(n372), .A2(A[10]), .X(n566) );
  SEN_ND2_G_1 U827 ( .A1(n372), .A2(A[9]), .X(n571) );
  SEN_ND2_G_1 U828 ( .A1(n372), .A2(A[17]), .X(n689) );
  SEN_ND2_G_1 U829 ( .A1(n372), .A2(A[18]), .X(n695) );
  SEN_ND2_G_1 U830 ( .A1(n372), .A2(A[22]), .X(n711) );
  SEN_ND2_G_1 U831 ( .A1(n372), .A2(A[21]), .X(n717) );
  SEN_ND2_G_1 U832 ( .A1(n372), .A2(A[24]), .X(n732) );
  SEN_ND2_G_1 U833 ( .A1(n372), .A2(A[30]), .X(n777) );
  SEN_AOI21_T_1 U834 ( .A1(n372), .A2(A[16]), .B(n683), .X(n987) );
  SEN_AOAI211_3 U835 ( .A1(n840), .A2(n858), .B(n374), .C(n487), .X(n486) );
  SEN_OAI211_1 U836 ( .A1(n374), .A2(n549), .B1(n844), .B2(n843), .X(n845) );
  SEN_INV_S_1 U837 ( .A(n374), .X(n841) );
  SEN_AO21_4 U838 ( .A1(n560), .A2(n638), .B(n1050), .X(n377) );
  SEN_OA21_2 U839 ( .A1(n562), .A2(n530), .B(n375), .X(n376) );
  SEN_ND2_4 U840 ( .A1(n966), .A2(n965), .X(n636) );
  SEN_INV_3 U841 ( .A(n636), .X(n379) );
  SEN_NR2_T_4 U842 ( .A1(n378), .A2(n379), .X(n654) );
  SEN_INV_3 U843 ( .A(n791), .X(n380) );
  SEN_ND2B_V1_6 U844 ( .A(n562), .B(n380), .X(n538) );
  SEN_EO2_2 U845 ( .A1(n554), .A2(A[4]), .X(n385) );
  SEN_ND2_G_1 U846 ( .A1(n533), .A2(n384), .X(n383) );
  SEN_ND2_G_1 U847 ( .A1(n536), .A2(n385), .X(n382) );
  SEN_ND3_T_2 U848 ( .A1(n382), .A2(n383), .A3(n779), .X(n381) );
  SEN_AOI21_T_3 U849 ( .A1(n539), .A2(A[4]), .B(n381), .X(n1020) );
  SEN_NR2_T_4 U850 ( .A1(n545), .A2(n386), .X(n1019) );
  SEN_MUXI2_S_4 U851 ( .D0(n361), .D1(n387), .S(B[4]), .X(n386) );
  SEN_EO2_2 U852 ( .A1(n1019), .A2(n1020), .X(n1022) );
  SEN_AN2_6 U853 ( .A1(n454), .A2(n557), .X(n542) );
  SEN_INV_10 U854 ( .A(n542), .X(n387) );
  SEN_INV_4 U855 ( .A(n542), .X(n541) );
  SEN_MUXI2_DG_2 U856 ( .D0(n361), .D1(n387), .S(B[5]), .X(n422) );
  SEN_MUXI2_DG_2 U857 ( .D0(n361), .D1(n387), .S(B[1]), .X(n643) );
  SEN_MUXI2_S_2 U858 ( .D0(n361), .D1(n387), .S(B[11]), .X(n578) );
  SEN_MUXI2_S_2 U859 ( .D0(n543), .D1(n387), .S(B[10]), .X(n558) );
  SEN_MUXI2_S_2 U860 ( .D0(n543), .D1(n387), .S(B[0]), .X(n639) );
  SEN_MUXI2_S_2 U861 ( .D0(n361), .D1(n387), .S(B[14]), .X(n606) );
  SEN_MUXI2_S_1 U862 ( .D0(n543), .D1(n387), .S(B[19]), .X(n668) );
  SEN_MUXI2_S_1 U863 ( .D0(n543), .D1(n387), .S(B[13]), .X(n600) );
  SEN_MUXI2_S_1 U864 ( .D0(n543), .D1(n387), .S(B[15]), .X(n594) );
  SEN_MUXI2_S_1 U865 ( .D0(n361), .D1(n387), .S(B[8]), .X(n587) );
  SEN_MUXI2_S_1 U866 ( .D0(n361), .D1(n387), .S(B[12]), .X(n584) );
  SEN_MUXI2_S_1 U867 ( .D0(n543), .D1(n387), .S(B[9]), .X(n572) );
  SEN_EO2_2 U868 ( .A1(n388), .A2(n1031), .X(n525) );
  SEN_NR2_T_4 U869 ( .A1(n390), .A2(n998), .X(n410) );
  SEN_ND2_T_4 U870 ( .A1(n390), .A2(n488), .X(n483) );
  SEN_EO2_S_0P5 U871 ( .A1(n997), .A2(n390), .X(n1006) );
  SEN_ND3_T_4 U872 ( .A1(n482), .A2(n483), .A3(n484), .X(n391) );
  SEN_NR2_T_3 U873 ( .A1(n391), .A2(n395), .X(n392) );
  SEN_EO2_1 U874 ( .A1(n988), .A2(n391), .X(n436) );
  SEN_OAI21_S_4 U875 ( .A1(n392), .A2(n396), .B(n397), .X(n393) );
  SEN_NR2_T_4 U876 ( .A1(n392), .A2(n879), .X(n970) );
  SEN_EO2_1 U877 ( .A1(n868), .A2(n394), .X(n399) );
  SEN_NR4_6 U878 ( .A1(Z[20]), .A2(Z[25]), .A3(n510), .A4(Z[27]), .X(n509) );
  SEN_ND3_T_1 U879 ( .A1(n703), .A2(n906), .A3(n699), .X(n395) );
  SEN_ND2_T_1P5 U880 ( .A1(n878), .A2(n880), .X(n396) );
  SEN_AOI21_S_1 U881 ( .A1(n996), .A2(n930), .B(n933), .X(n413) );
  SEN_ND2_G_1 U882 ( .A1(n928), .A2(n930), .X(n412) );
  SEN_AOI21_S_4 U883 ( .A1(n418), .A2(n924), .B(n828), .X(n419) );
  SEN_AOI21_3 U884 ( .A1(n414), .A2(n978), .B(n498), .X(n497) );
  SEN_AOI22_T_3 U885 ( .A1(n414), .A2(n415), .B1(n910), .B2(n909), .X(n951) );
  SEN_ND3_T_2 U886 ( .A1(n434), .A2(n433), .A3(n417), .X(Z[16]) );
  SEN_ND3_T_2 U887 ( .A1(n416), .A2(n499), .A3(n513), .X(n512) );
  SEN_EO2_1 U888 ( .A1(n920), .A2(n418), .X(n927) );
  SEN_OAI21_3 U889 ( .A1(n419), .A2(n919), .B(n829), .X(n839) );
  SEN_ND2_2 U890 ( .A1(n638), .A2(n789), .X(n1049) );
  SEN_ND2_G_1 U891 ( .A1(n1052), .A2(n529), .X(n420) );
  SEN_AN3B_1 U892 ( .B1(n918), .B2(n1010), .A(n917), .X(n425) );
  SEN_ND2_2 U893 ( .A1(n426), .A2(n367), .X(n423) );
  SEN_ND2_G_1 U894 ( .A1(n536), .A2(n430), .X(n429) );
  SEN_AOI21_S_1 U895 ( .A1(n533), .A2(n431), .B(n364), .X(n428) );
  SEN_ND2_2 U896 ( .A1(n436), .A2(n367), .X(n433) );
  SEN_AO21B_2 U897 ( .A1(n442), .A2(n367), .B(n437), .X(Z[10]) );
  SEN_EN2_3 U898 ( .A1(n527), .A2(n951), .X(n443) );
  SEN_OAI21_3 U899 ( .A1(n443), .A2(n444), .B(n445), .X(Z[19]) );
  SEN_OA21_2 U900 ( .A1(n970), .A2(n881), .B(n880), .X(n453) );
  SEN_EN2_3 U901 ( .A1(n884), .A2(n453), .X(n448) );
  SEN_MUXI2_S_4 U902 ( .D0(n1052), .D1(n529), .S(n530), .X(n454) );
  SEN_AOI21_3 U903 ( .A1(n1029), .A2(n525), .B(n389), .X(n1025) );
  SEN_NR3_G_1 U904 ( .A1(n1027), .A2(n1026), .A3(n1053), .X(n458) );
  SEN_EO2_S_0P5 U905 ( .A1(n1028), .A2(n1025), .X(n459) );
  SEN_ND2_G_1 U906 ( .A1(n459), .A2(n1058), .X(n456) );
  SEN_OAI211_1 U907 ( .A1(n1036), .A2(n1028), .B1(n456), .B2(n457), .X(Z[3])
         );
  SEN_NR2_T_3 U908 ( .A1(n930), .A2(n933), .X(n658) );
  SEN_ND3_T_4 U909 ( .A1(n461), .A2(n462), .A3(n463), .X(n1011) );
  SEN_ND2_4 U910 ( .A1(n536), .A2(n464), .X(n463) );
  SEN_EO2_2 U911 ( .A1(n1009), .A2(n1011), .X(n1015) );
  SEN_ND2_G_3 U912 ( .A1(n969), .A2(n636), .X(n477) );
  SEN_ND3_2 U913 ( .A1(n934), .A2(n635), .A3(n636), .X(n476) );
  SEN_ND4_1 U914 ( .A1(n1015), .A2(n635), .A3(n636), .A4(n942), .X(n475) );
  SEN_ND3_T_2 U915 ( .A1(n475), .A2(n476), .A3(n477), .X(n474) );
  SEN_OAI22_3 U916 ( .A1(n655), .A2(n938), .B1(n1022), .B2(n960), .X(n473) );
  SEN_AOI21_3 U917 ( .A1(n473), .A2(n654), .B(n474), .X(n467) );
  SEN_ND3_2 U918 ( .A1(n656), .A2(n928), .A3(n840), .X(n489) );
  SEN_OAI21_G_2 U919 ( .A1(n661), .A2(n838), .B(n486), .X(n485) );
  SEN_NR3_T_3 U920 ( .A1(n489), .A2(n658), .A3(n657), .X(n488) );
  SEN_NR2_1 U921 ( .A1(n924), .A2(n828), .X(n480) );
  SEN_NR2_2 U922 ( .A1(n658), .A2(n657), .X(n478) );
  SEN_AOI21_T_2 U923 ( .A1(n662), .A2(n919), .B(n485), .X(n484) );
  SEN_AOI22_T_2 U924 ( .A1(n478), .A2(n479), .B1(n662), .B2(n480), .X(n482) );
  SEN_NR4_3 U925 ( .A1(Z[3]), .A2(Z[2]), .A3(Z[1]), .A4(Z[0]), .X(n513) );
  SEN_INV_S_1 U926 ( .A(Z[8]), .X(n500) );
  SEN_NR3_T_2 U927 ( .A1(n512), .A2(Z[5]), .A3(Z[9]), .X(n511) );
  SEN_NR4_3 U928 ( .A1(Z[22]), .A2(Z[21]), .A3(Z[17]), .A4(Z[6]), .X(n503) );
  SEN_INV_S_1 U929 ( .A(Z[7]), .X(n515) );
  SEN_OR4B_4 U930 ( .B1(n508), .B2(Z[26]), .B3(Z[13]), .A(n509), .X(n506) );
  SEN_OA21_1 U931 ( .A1(n810), .A2(n549), .B(n808), .X(n517) );
  SEN_EN2_S_2 U932 ( .A1(n866), .A2(n859), .X(n518) );
  SEN_ND2_2 U933 ( .A1(n518), .A2(n367), .X(n865) );
  SEN_OA21_1 U934 ( .A1(n549), .A2(n905), .B(n903), .X(n519) );
  SEN_ND3_S_4 U935 ( .A1(n949), .A2(n522), .A3(n948), .X(Z[6]) );
  SEN_INV_2 U936 ( .A(n675), .X(n524) );
  SEN_EO2_5 U937 ( .A1(n523), .A2(n524), .X(n527) );
  SEN_AN2_S_3 U938 ( .A1(n530), .A2(n529), .X(n786) );
  SEN_AOI21_G_4 U939 ( .A1(n539), .A2(A[2]), .B(n653), .X(n1031) );
  SEN_NR2_T_3 U940 ( .A1(n690), .A2(n546), .X(n916) );
  SEN_AOI22_T_3 U941 ( .A1(n811), .A2(n812), .B1(n771), .B2(n770), .X(n803) );
  SEN_INV_5 U942 ( .A(n773), .X(n534) );
  SEN_EO2_1 U943 ( .A1(n554), .A2(A[7]), .X(n628) );
  SEN_NR2_T_4 U944 ( .A1(n560), .A2(n559), .X(n1046) );
  SEN_INV_3 U945 ( .A(n530), .X(n789) );
  SEN_EO2_1 U946 ( .A1(n554), .A2(A[1]), .X(n644) );
  SEN_INV_S_12 U947 ( .A(n534), .X(n532) );
  SEN_ND3_T_2 U948 ( .A1(n619), .A2(n618), .A3(n617), .X(n623) );
  SEN_ND2_T_1 U949 ( .A1(n536), .A2(n616), .X(n617) );
  SEN_INV_4 U950 ( .A(n635), .X(n960) );
  SEN_ND2_T_2 U951 ( .A1(n1052), .A2(n531), .X(n562) );
  SEN_ND2_2 U952 ( .A1(n932), .A2(n586), .X(n827) );
  SEN_ND2_G_4 U953 ( .A1(n999), .A2(n593), .X(n928) );
  SEN_NR2_T_2 U954 ( .A1(n559), .A2(n530), .X(n773) );
  SEN_ND2_T_1P5 U955 ( .A1(n621), .A2(n360), .X(n622) );
  SEN_NR2_T_3 U956 ( .A1(n578), .A2(n545), .X(n921) );
  SEN_NR2_S_5 U957 ( .A1(n854), .A2(n853), .X(n847) );
  SEN_ND3_T_2 U958 ( .A1(n571), .A2(n570), .A3(n569), .X(n992) );
  SEN_BUF_6 U959 ( .A(INST[1]), .X(n530) );
  SEN_ND2_S_4 U960 ( .A1(n1011), .A2(n624), .X(n942) );
  SEN_AOI31_0P5 U961 ( .A1(n1010), .A2(n965), .A3(n966), .B(n528), .X(n967) );
  SEN_NR2_T_4 U962 ( .A1(n660), .A2(n837), .X(n656) );
  SEN_AOI22_T_1P5 U963 ( .A1(n698), .A2(n527), .B1(n677), .B2(n959), .X(n703)
         );
  SEN_OAI211_3 U964 ( .A1(n959), .A2(n549), .B1(n958), .B2(n957), .X(Z[20]) );
  SEN_INV_2 U965 ( .A(n917), .X(n585) );
  SEN_NR2_S_5 U966 ( .A1(n661), .A2(n607), .X(n662) );
  SEN_ND2_G_3 U967 ( .A1(n945), .A2(n944), .X(n635) );
  SEN_EO2_2 U968 ( .A1(n634), .A2(n945), .X(n934) );
  SEN_EO2_2 U969 ( .A1(n554), .A2(A[6]), .X(n609) );
  SEN_AOI21_T_3 U970 ( .A1(n539), .A2(A[1]), .B(n648), .X(n1039) );
  SEN_INV_3 U971 ( .A(n1009), .X(n624) );
  SEN_AOI21_3 U972 ( .A1(n869), .A2(n868), .B(n867), .X(n870) );
  SEN_OAI211_3 U973 ( .A1(n877), .A2(n1044), .B1(n876), .B2(n875), .X(Z[26])
         );
  SEN_ND3_T_3 U974 ( .A1(n631), .A2(n630), .A3(n629), .X(n966) );
  SEN_ND2_T_1 U975 ( .A1(n536), .A2(n628), .X(n629) );
  SEN_INV_12 U976 ( .A(n544), .X(n543) );
  SEN_INV_AS_2 U977 ( .A(n1001), .X(n593) );
  SEN_EO2_5 U978 ( .A1(n1001), .A2(n999), .X(n998) );
  SEN_ND3_S_4 U979 ( .A1(n695), .A2(n694), .A3(n693), .X(n915) );
  SEN_MUXI2_S_1 U980 ( .D0(n543), .D1(n541), .S(B[24]), .X(n727) );
  SEN_MUXI2_S_1 U981 ( .D0(n361), .D1(n541), .S(B[23]), .X(n719) );
  SEN_ND2_G_1 U982 ( .A1(n535), .A2(n669), .X(n672) );
  SEN_INV_4 U983 ( .A(n538), .X(n535) );
  SEN_MUXI2_S_2 U984 ( .D0(n543), .D1(n541), .S(B[17]), .X(n684) );
  SEN_MUXI2_S_2 U985 ( .D0(n543), .D1(n541), .S(B[18]), .X(n690) );
  SEN_AOI21_S_2 U986 ( .A1(n1016), .A2(n1022), .B(n941), .X(n1007) );
  SEN_ND2_G_3 U987 ( .A1(n633), .A2(n360), .X(n965) );
  SEN_ND2_2 U988 ( .A1(n635), .A2(n939), .X(n655) );
  SEN_ND2_T_4 U989 ( .A1(n937), .A2(n936), .X(n1029) );
  SEN_EO2_1 U990 ( .A1(n961), .A2(n962), .X(n943) );
  SEN_EO2_2 U991 ( .A1(n986), .A2(n987), .X(n906) );
  SEN_ND3_T_2 U992 ( .A1(n689), .A2(n688), .A3(n687), .X(n981) );
  SEN_ND2_T_1 U993 ( .A1(n536), .A2(n602), .X(n603) );
  SEN_NR2_T_1P5 U994 ( .A1(n985), .A2(n914), .X(n699) );
  SEN_EO2_2 U995 ( .A1(n921), .A2(n922), .X(n924) );
  SEN_AOI21_T_3 U996 ( .A1(n539), .A2(A[13]), .B(n599), .X(n832) );
  SEN_AOI21_T_3 U997 ( .A1(n539), .A2(A[11]), .B(n577), .X(n922) );
  SEN_EO2_2 U998 ( .A1(n898), .A2(n897), .X(n899) );
  SEN_INV_2 U999 ( .A(n935), .X(n936) );
  SEN_NR2_2 U1000 ( .A1(n1039), .A2(n1038), .X(n935) );
  SEN_OAI21_S_3 U1001 ( .A1(n705), .A2(n704), .B(n703), .X(n878) );
  SEN_ND2_T_1 U1002 ( .A1(n533), .A2(n721), .X(n722) );
  SEN_ND2_T_1 U1003 ( .A1(n533), .A2(n650), .X(n651) );
  SEN_ND2_G_3 U1004 ( .A1(n533), .A2(n596), .X(n597) );
  SEN_EO2_2 U1005 ( .A1(n838), .A2(n839), .X(n830) );
  SEN_EO2_5 U1006 ( .A1(n931), .A2(n932), .X(n933) );
  SEN_ND3_3 U1007 ( .A1(n566), .A2(n565), .A3(n564), .X(n932) );
  SEN_ND2_T_1P5 U1008 ( .A1(n536), .A2(n595), .X(n598) );
  SEN_ND3_1 U1009 ( .A1(n682), .A2(n779), .A3(n681), .X(n683) );
  SEN_INV_2 U1010 ( .A(n1020), .X(n626) );
  SEN_ND2_G_3 U1011 ( .A1(n626), .A2(n625), .X(n940) );
  SEN_OAI211_3 U1012 ( .A1(n866), .A2(n549), .B1(n865), .B2(n864), .X(Z[27])
         );
  SEN_ND3_T_2 U1013 ( .A1(n598), .A2(n779), .A3(n597), .X(n599) );
  SEN_ND2_2 U1014 ( .A1(n614), .A2(n360), .X(n944) );
  SEN_INV_2 U1015 ( .A(n1019), .X(n625) );
  SEN_BUF_6 U1016 ( .A(INST[2]), .X(n531) );
  SEN_BUF_6 U1017 ( .A(INST[0]), .X(n529) );
  SEN_EO2_2 U1018 ( .A1(n959), .A2(n952), .X(n953) );
  SEN_OA21B_2 U1019 ( .A1(n951), .A2(n527), .B(n950), .X(n952) );
  SEN_EO2_2 U1020 ( .A1(n554), .A2(A[13]), .X(n595) );
  SEN_EO2_2 U1021 ( .A1(n810), .A2(n803), .X(n804) );
  SEN_ND2_2 U1022 ( .A1(n971), .A2(n367), .X(n976) );
  SEN_ND2_T_5 U1023 ( .A1(n529), .A2(n531), .X(n559) );
  SEN_INV_10 U1024 ( .A(n360), .X(n546) );
  SEN_INV_2 U1025 ( .A(n878), .X(n879) );
  SEN_INV_3 U1026 ( .A(n659), .X(n854) );
  SEN_ND3_T_3 U1027 ( .A1(n605), .A2(n604), .A3(n603), .X(n659) );
  SEN_NR2_T_1P5 U1028 ( .A1(n639), .A2(n545), .X(n1054) );
  SEN_EO2_2 U1029 ( .A1(n812), .A2(n811), .X(n813) );
  SEN_AOI21_T_1 U1030 ( .A1(n539), .A2(A[23]), .B(n724), .X(n890) );
  SEN_INV_S_8 U1031 ( .A(n538), .X(n536) );
  SEN_AOI21_S_2 U1032 ( .A1(n539), .A2(A[19]), .B(n667), .X(n912) );
  SEN_ND3_1 U1033 ( .A1(n666), .A2(n779), .A3(n665), .X(n667) );
  SEN_EO2_1 U1034 ( .A1(n554), .A2(A[19]), .X(n663) );
  SEN_EO2_2 U1035 ( .A1(n991), .A2(n992), .X(n996) );
  SEN_EO2_1 U1036 ( .A1(n977), .A2(n970), .X(n971) );
  SEN_NR2_T_3 U1037 ( .A1(n606), .A2(n545), .X(n853) );
  SEN_EO2_2 U1038 ( .A1(n853), .A2(n659), .X(n858) );
  SEN_ND3_T_2 U1039 ( .A1(n652), .A2(n779), .A3(n651), .X(n653) );
  SEN_EO2_1 U1040 ( .A1(n554), .A2(A[2]), .X(n649) );
  SEN_ND2_T_1 U1041 ( .A1(n536), .A2(n573), .X(n576) );
  SEN_ND3_T_2 U1042 ( .A1(n576), .A2(n779), .A3(n575), .X(n577) );
  SEN_EO2_2 U1043 ( .A1(n555), .A2(A[11]), .X(n573) );
  SEN_ND3_2 U1044 ( .A1(n647), .A2(n779), .A3(n646), .X(n648) );
  SEN_EO2_1 U1045 ( .A1(n858), .A2(n851), .X(n852) );
  SEN_OAI211_1 U1046 ( .A1(n1036), .A2(n996), .B1(n995), .B2(n994), .X(Z[9])
         );
  SEN_EO2_2 U1047 ( .A1(n831), .A2(n832), .X(n838) );
  SEN_OAI21_S_3 U1048 ( .A1(n1025), .A2(n1028), .B(n939), .X(n1016) );
  SEN_AOI21_2 U1049 ( .A1(n962), .A2(n961), .B(n960), .X(n963) );
  SEN_NR2_T_3 U1050 ( .A1(n558), .A2(n545), .X(n931) );
  SEN_INV_3 U1051 ( .A(n623), .X(n1027) );
  SEN_NR3_G_1 U1052 ( .A1(n854), .A2(n853), .A3(n366), .X(n855) );
  SEN_ND3_T_0P8 U1053 ( .A1(n859), .A2(n860), .A3(n823), .X(n764) );
  SEN_NR3_G_1 U1054 ( .A1(n1039), .A2(n1038), .A3(n1053), .X(n1040) );
  SEN_OAI31_G_1 U1055 ( .A1(n1020), .A2(n526), .A3(n1053), .B(n1018), .X(n1021) );
  SEN_NR2_1 U1056 ( .A1(n791), .A2(n790), .X(n1010) );
  SEN_NR3_G_1 U1057 ( .A1(n790), .A2(n1050), .A3(n530), .X(n1057) );
  SEN_EO2_S_0P5 U1058 ( .A1(n553), .A2(A[18]), .X(n692) );
  SEN_AOI21_S_1 U1059 ( .A1(n539), .A2(A[25]), .B(n737), .X(n826) );
  SEN_OAI21_S_0P5 U1060 ( .A1(n534), .A2(n553), .B(n779), .X(n780) );
  SEN_OAI211_1 U1061 ( .A1(n802), .A2(n799), .B1(n796), .B2(n784), .X(n783) );
  SEN_OAI21_G_1 U1062 ( .A1(n549), .A2(n796), .B(n795), .X(n797) );
  SEN_ND2_G_1 U1063 ( .A1(n536), .A2(n774), .X(n775) );
  SEN_ND2_G_1 U1064 ( .A1(n535), .A2(n757), .X(n760) );
  SEN_ND2_G_1 U1065 ( .A1(n532), .A2(n766), .X(n767) );
  SEN_ND2_G_1 U1066 ( .A1(n535), .A2(n765), .X(n768) );
  SEN_INV_S_1 U1067 ( .A(n360), .X(n547) );
  SEN_ND2_G_1 U1068 ( .A1(n990), .A2(n367), .X(n995) );
  SEN_ND2_G_1 U1069 ( .A1(n1008), .A2(n367), .X(n1014) );
  SEN_OAI211_1 U1070 ( .A1(n1045), .A2(n1044), .B1(n1043), .B2(n1042), .X(Z[1]) );
  SEN_OAI211_1 U1071 ( .A1(n1036), .A2(n1035), .B1(n1034), .B2(n1033), .X(Z[2]) );
  SEN_ND2_G_1 U1072 ( .A1(n1030), .A2(n1058), .X(n1034) );
  SEN_OAI21_G_1 U1073 ( .A1(n1006), .A2(n1044), .B(n1005), .X(Z[8]) );
  SEN_OAI21_G_1 U1074 ( .A1(n1002), .A2(n1001), .B(n1000), .X(n1003) );
  SEN_ND2_G_1 U1075 ( .A1(n999), .A2(n1010), .X(n1002) );
  SEN_NR2_1 U1076 ( .A1(n998), .A2(n549), .X(n1004) );
  SEN_ND2_G_1 U1077 ( .A1(n924), .A2(n548), .X(n925) );
  SEN_ND2_G_1 U1078 ( .A1(n535), .A2(n752), .X(n755) );
  SEN_ND2_G_1 U1079 ( .A1(n535), .A2(n733), .X(n736) );
  SEN_ND2_G_1 U1080 ( .A1(n532), .A2(n742), .X(n743) );
  SEN_ND2_G_1 U1081 ( .A1(n535), .A2(n741), .X(n744) );
  SEN_ND2_G_1 U1082 ( .A1(n979), .A2(n367), .X(n984) );
  SEN_ND2_G_1 U1083 ( .A1(n961), .A2(n548), .X(n948) );
  SEN_ND2_G_1 U1084 ( .A1(n943), .A2(n367), .X(n949) );
  SEN_ND2_G_1 U1085 ( .A1(n964), .A2(n367), .X(n968) );
  SEN_ND2_G_1 U1086 ( .A1(n535), .A2(n729), .X(n730) );
  SEN_ND2_G_1 U1087 ( .A1(n913), .A2(n908), .X(n910) );
  SEN_ND2_G_1 U1088 ( .A1(n535), .A2(n714), .X(n715) );
  SEN_ND2_G_1 U1089 ( .A1(n535), .A2(n708), .X(n709) );
  SEN_NR2_1 U1090 ( .A1(n702), .A2(n907), .X(n704) );
  SEN_OAI211_1 U1091 ( .A1(n914), .A2(n913), .B1(n698), .B2(n908), .X(n705) );
  SEN_ND2_G_1 U1092 ( .A1(n697), .A2(n915), .X(n908) );
  SEN_ND2_G_1 U1093 ( .A1(n696), .A2(n981), .X(n913) );
  SEN_ND2_G_1 U1094 ( .A1(n535), .A2(n692), .X(n693) );
  SEN_ND2_G_1 U1095 ( .A1(n535), .A2(n686), .X(n687) );
  SEN_ND2_G_1 U1096 ( .A1(n533), .A2(n680), .X(n681) );
  SEN_ND2_G_1 U1097 ( .A1(n535), .A2(n679), .X(n682) );
  SEN_ND2_G_1 U1098 ( .A1(n533), .A2(n670), .X(n671) );
  SEN_NR2_1 U1099 ( .A1(n912), .A2(n911), .X(n950) );
  SEN_ND2_G_1 U1100 ( .A1(n533), .A2(n664), .X(n665) );
  SEN_ND2_G_1 U1101 ( .A1(n536), .A2(n663), .X(n666) );
  SEN_ND2_G_1 U1102 ( .A1(n536), .A2(n649), .X(n652) );
  SEN_ND2_G_1 U1103 ( .A1(n533), .A2(n645), .X(n646) );
  SEN_ND2_G_1 U1104 ( .A1(n536), .A2(n644), .X(n647) );
  SEN_OAI21_G_1 U1105 ( .A1(n639), .A2(n1047), .B(n640), .X(n642) );
  SEN_ND2_G_1 U1106 ( .A1(n540), .A2(A[14]), .X(n605) );
  SEN_ND2_G_1 U1107 ( .A1(n536), .A2(n589), .X(n590) );
  SEN_ND2_G_1 U1108 ( .A1(n536), .A2(n580), .X(n581) );
  SEN_ND2_G_1 U1109 ( .A1(n540), .A2(A[12]), .X(n583) );
  SEN_ND2_G_1 U1110 ( .A1(n533), .A2(n574), .X(n575) );
  SEN_ND2_G_1 U1111 ( .A1(n537), .A2(n568), .X(n569) );
  SEN_ND2_G_1 U1112 ( .A1(n535), .A2(n563), .X(n564) );
  SEN_ND2_G_1 U1113 ( .A1(n535), .A2(n720), .X(n723) );
  SEN_AOI21_S_1 U1114 ( .A1(n539), .A2(n553), .B(n780), .X(n793) );
  SEN_AOI21_S_1 U1115 ( .A1(n532), .A2(n772), .B(n364), .X(n776) );
  SEN_AOI21_S_1 U1116 ( .A1(n539), .A2(A[28]), .B(n761), .X(n822) );
  SEN_EO2_S_0P5 U1117 ( .A1(n553), .A2(A[28]), .X(n757) );
  SEN_AOI21_S_1 U1118 ( .A1(n539), .A2(A[29]), .B(n769), .X(n815) );
  SEN_AN3B_1 U1119 ( .B1(n992), .B2(n1010), .A(n991), .X(n993) );
  SEN_EN2_0P5 U1120 ( .A1(n1041), .A2(n1037), .X(n1045) );
  SEN_AOI21_S_1 U1121 ( .A1(n1022), .A2(n548), .B(n1021), .X(n1023) );
  SEN_EO2_S_0P5 U1122 ( .A1(n1017), .A2(n1016), .X(n1024) );
  SEN_INV_S_1 U1123 ( .A(n1022), .X(n1017) );
  SEN_AOI21_S_1 U1124 ( .A1(n539), .A2(A[27]), .B(n756), .X(n862) );
  SEN_EO2_S_0P5 U1125 ( .A1(n553), .A2(A[27]), .X(n752) );
  SEN_MUXI2_S_1 U1126 ( .D0(n543), .D1(n541), .S(B[27]), .X(n751) );
  SEN_EO2_S_0P5 U1127 ( .A1(n554), .A2(A[25]), .X(n733) );
  SEN_MUXI2_S_1 U1128 ( .D0(n361), .D1(n541), .S(B[25]), .X(n738) );
  SEN_AOI21_S_1 U1129 ( .A1(n539), .A2(A[26]), .B(n745), .X(n872) );
  SEN_EO2_S_0P5 U1130 ( .A1(n553), .A2(A[26]), .X(n741) );
  SEN_MUXI2_S_1 U1131 ( .D0(n361), .D1(n541), .S(B[26]), .X(n740) );
  SEN_AN3B_1 U1132 ( .B1(n981), .B2(n1010), .A(n980), .X(n982) );
  SEN_ND3_S_0P5 U1133 ( .A1(n945), .A2(n944), .A3(n1010), .X(n946) );
  SEN_AN3B_1 U1134 ( .B1(n973), .B2(n1010), .A(n972), .X(n974) );
  SEN_INV_S_1 U1135 ( .A(n934), .X(n961) );
  SEN_INV_S_1 U1136 ( .A(n940), .X(n941) );
  SEN_AOI21_S_1 U1137 ( .A1(n532), .A2(n728), .B(n365), .X(n731) );
  SEN_EO2_S_0P5 U1138 ( .A1(n553), .A2(A[21]), .X(n714) );
  SEN_AOI21_S_1 U1139 ( .A1(n532), .A2(n713), .B(n365), .X(n716) );
  SEN_MUXI2_S_1 U1140 ( .D0(n543), .D1(n541), .S(B[21]), .X(n712) );
  SEN_EO2_S_0P5 U1141 ( .A1(n553), .A2(A[22]), .X(n708) );
  SEN_AOI21_S_1 U1142 ( .A1(n532), .A2(n707), .B(n365), .X(n710) );
  SEN_MUXI2_S_1 U1143 ( .D0(n361), .D1(n541), .S(B[22]), .X(n706) );
  SEN_INV_S_1 U1144 ( .A(n970), .X(n887) );
  SEN_AOI21_S_1 U1145 ( .A1(n532), .A2(n691), .B(n364), .X(n694) );
  SEN_EO2_S_0P5 U1146 ( .A1(n554), .A2(A[17]), .X(n686) );
  SEN_AOI21_S_1 U1147 ( .A1(n532), .A2(n685), .B(n364), .X(n688) );
  SEN_EO2_S_0P5 U1148 ( .A1(n554), .A2(A[16]), .X(n679) );
  SEN_MUXI2_S_1 U1149 ( .D0(n543), .D1(n541), .S(B[16]), .X(n678) );
  SEN_INV_S_1 U1150 ( .A(n912), .X(n675) );
  SEN_EO2_S_0P5 U1151 ( .A1(n554), .A2(A[20]), .X(n669) );
  SEN_AOI22_1 U1152 ( .A1(n540), .A2(A[0]), .B1(n535), .B2(n637), .X(n1048) );
  SEN_EO2_S_0P5 U1153 ( .A1(n554), .A2(A[0]), .X(n637) );
  SEN_MUXI2_S_1 U1154 ( .D0(n542), .D1(n544), .S(n632), .X(n633) );
  SEN_AOI21_S_1 U1155 ( .A1(n532), .A2(n627), .B(n363), .X(n630) );
  SEN_MUXI2_S_1 U1156 ( .D0(n542), .D1(n544), .S(n620), .X(n621) );
  SEN_AOI21_S_1 U1157 ( .A1(n532), .A2(n615), .B(n365), .X(n618) );
  SEN_AOI21_S_1 U1158 ( .A1(n532), .A2(n601), .B(n365), .X(n604) );
  SEN_EO2_S_0P5 U1159 ( .A1(n555), .A2(A[8]), .X(n589) );
  SEN_AOI21_S_1 U1160 ( .A1(n532), .A2(n579), .B(n365), .X(n582) );
  SEN_INV_S_1 U1161 ( .A(n538), .X(n537) );
  SEN_AOI21_S_1 U1162 ( .A1(n533), .A2(n567), .B(n365), .X(n570) );
  SEN_EO2_S_0P5 U1163 ( .A1(n553), .A2(A[10]), .X(n563) );
  SEN_AOI21_S_1 U1164 ( .A1(n532), .A2(n561), .B(n364), .X(n565) );
  SEN_OA21_1 U1165 ( .A1(B[7]), .A2(A[7]), .B(n1057), .X(n528) );
  SEN_TIE0_1 U1166 ( .X(FLAGS[3]) );
endmodule

