
module Alu ( Z, A, B, INST, SEL );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  input SEL;
  wire   n216, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388;

  SEN_NR2_T_2 U263 ( .A1(n646), .A2(n645), .X(n652) );
  SEN_ND2_S_3 U264 ( .A1(n1366), .A2(n1315), .X(n1264) );
  SEN_NR2_S_0P65 U265 ( .A1(n467), .A2(n271), .X(n456) );
  SEN_NR2B_V1_1 U266 ( .A(n809), .B(n832), .X(n433) );
  SEN_AOI21B_3 U267 ( .A1(n811), .A2(n810), .B(n809), .X(n817) );
  SEN_AN4B_1 U268 ( .B1(n918), .B2(n988), .B3(n483), .A(n482), .X(n517) );
  SEN_AOAI211_0P75 U269 ( .A1(n638), .A2(n656), .B(n488), .C(n487), .X(n502)
         );
  SEN_AOI211_G_1 U270 ( .A1(n503), .A2(n502), .B1(n501), .B2(n500), .X(n504)
         );
  SEN_ND2_G_0P65 U271 ( .A1(n414), .A2(n272), .X(n1245) );
  SEN_BUF_1P5 U272 ( .A(n592), .X(n256) );
  SEN_AOAI211_1 U273 ( .A1(n428), .A2(n427), .B(n426), .C(n425), .X(n432) );
  SEN_AOAI211_G_3 U274 ( .A1(n652), .A2(n651), .B(n650), .C(n649), .X(n301) );
  SEN_ND2_S_0P8 U275 ( .A1(n421), .A2(n1293), .X(n1273) );
  SEN_ND2B_V1DG_1 U276 ( .A(n669), .B(n668), .X(n670) );
  SEN_ND2_G_0P65 U277 ( .A1(n674), .A2(n673), .X(Z[5]) );
  SEN_AN2_S_0P5 U278 ( .A1(n332), .A2(n1381), .X(n235) );
  SEN_NR2B_V1_4 U279 ( .A(n235), .B(n1330), .X(n252) );
  SEN_INV_6 U280 ( .A(n1297), .X(n1330) );
  SEN_MUXI2_S_4 U281 ( .D0(n1300), .D1(n1299), .S(n400), .X(n1301) );
  SEN_OR2_1P5 U282 ( .A1(n379), .A2(n352), .X(n753) );
  SEN_BUF_S_4 U283 ( .A(B[8]), .X(n352) );
  SEN_ND2_T_2 U284 ( .A1(n819), .A2(n818), .X(n787) );
  SEN_ND2_3 U285 ( .A1(n779), .A2(n258), .X(n819) );
  SEN_BUF_S_3 U286 ( .A(A[2]), .X(n373) );
  SEN_ND2_G_1 U287 ( .A1(n626), .A2(n625), .X(n646) );
  SEN_ND2_S_0P5 U288 ( .A1(n372), .A2(n345), .X(n626) );
  SEN_MUXI2_DG_2 U289 ( .D0(n902), .D1(n1379), .S(n357), .X(n903) );
  SEN_ND3_S_2 U290 ( .A1(n291), .A2(n292), .A3(n406), .X(n902) );
  SEN_ND2_T_1 U291 ( .A1(n933), .A2(n900), .X(n906) );
  SEN_AOAI211_G_1 U292 ( .A1(n338), .A2(n1303), .B(n1302), .C(n1301), .X(Z[29]) );
  SEN_ND2B_1 U293 ( .A(n782), .B(n258), .X(n783) );
  SEN_INV_1P25 U294 ( .A(n257), .X(n258) );
  SEN_ND2_0P8 U295 ( .A1(n752), .A2(n751), .X(n782) );
  SEN_AN2_S_1 U296 ( .A1(n975), .A2(n974), .X(n981) );
  SEN_INV_S_3 U297 ( .A(n1065), .X(n285) );
  SEN_INV_1 U298 ( .A(n404), .X(n403) );
  SEN_OAI21_G_2 U299 ( .A1(n1295), .A2(n369), .B(n254), .X(n1300) );
  SEN_ND2_T_4 U300 ( .A1(n251), .A2(n252), .X(n1299) );
  SEN_ND2B_V1_3 U301 ( .A(n400), .B(n1330), .X(n1382) );
  SEN_INV_0P8 U302 ( .A(n1344), .X(n1283) );
  SEN_OAI21_3 U303 ( .A1(n1285), .A2(n1284), .B(n1305), .X(n1289) );
  SEN_ND2_T_4 U304 ( .A1(n301), .A2(n308), .X(n675) );
  SEN_AOAI211_0P5 U305 ( .A1(n1386), .A2(A[31]), .B(n1385), .C(n370), .X(n1387) );
  SEN_ND2_S_1P5 U306 ( .A1(n1388), .A2(n1387), .X(Z[31]) );
  SEN_ND2_T_0P5 U307 ( .A1(n1212), .A2(n1211), .X(n1213) );
  SEN_ND2_T_1 U308 ( .A1(n1261), .A2(n1260), .X(n323) );
  SEN_NR2B_V1_1 U309 ( .A(n1261), .B(n1238), .X(n524) );
  SEN_ND2B_V1_1 U310 ( .A(n398), .B(n367), .X(n1261) );
  SEN_ND2_G_1 U311 ( .A1(n463), .A2(n534), .X(n467) );
  SEN_ND2_T_1 U312 ( .A1(n329), .A2(n453), .X(n463) );
  SEN_INV_1 U313 ( .A(n1036), .X(n1037) );
  SEN_ND2B_1 U314 ( .A(n1039), .B(n1038), .X(n1040) );
  SEN_OAI21_S_2 U315 ( .A1(n1367), .A2(n323), .B(n1365), .X(n1368) );
  SEN_OAI22_T_1P5 U316 ( .A1(n1369), .A2(n402), .B1(n1368), .B2(n409), .X(
        n1386) );
  SEN_AN2_3 U317 ( .A1(n1378), .A2(n1377), .X(n253) );
  SEN_OAI21_T_0P5 U318 ( .A1(n1293), .A2(n417), .B(n1294), .X(n1270) );
  SEN_INV_S_6 U319 ( .A(n1244), .X(n1293) );
  SEN_INV_0P65 U320 ( .A(n408), .X(n407) );
  SEN_MUXI2_DG_1 U321 ( .D0(n1153), .D1(n1152), .S(n394), .X(n1154) );
  SEN_ND2_T_1 U322 ( .A1(n327), .A2(n1147), .X(n1153) );
  SEN_ND2_T_0P5 U323 ( .A1(n283), .A2(n284), .X(n899) );
  SEN_NR2_T_4 U324 ( .A1(n319), .A2(n1343), .X(n1354) );
  SEN_ND2_T_1 U325 ( .A1(n1249), .A2(n1248), .X(n1254) );
  SEN_ND3_T_1P5 U326 ( .A1(n1336), .A2(n1335), .A3(n1334), .X(Z[30]) );
  SEN_NR2B_V1_1 U327 ( .A(n633), .B(n486), .X(n427) );
  SEN_ND2B_V1_1 U328 ( .A(n374), .B(n347), .X(n633) );
  SEN_ND2_0P65 U329 ( .A1(n1063), .A2(n1195), .X(n1140) );
  SEN_BUF_S_1 U330 ( .A(n422), .X(n420) );
  SEN_ND2B_S_1 U331 ( .A(n1208), .B(n420), .X(n1230) );
  SEN_OAI21_G_0P5 U332 ( .A1(n791), .A2(n410), .B(n788), .X(n794) );
  SEN_ND3_S_2 U333 ( .A1(n304), .A2(n305), .A3(n406), .X(n1327) );
  SEN_OR2_1P5 U334 ( .A1(n1321), .A2(n242), .X(n304) );
  SEN_ND2B_S_8 U335 ( .A(n1296), .B(n420), .X(n1297) );
  SEN_OR3B_4 U336 ( .B1(n398), .B2(n399), .A(n1293), .X(n1296) );
  SEN_ND2_S_4 U337 ( .A1(n663), .A2(n306), .X(n307) );
  SEN_AOAI211_4 U338 ( .A1(n661), .A2(n660), .B(n659), .C(n658), .X(n663) );
  SEN_OAI21_S_3 U339 ( .A1(n1287), .A2(n1286), .B(n1316), .X(n1291) );
  SEN_INV_3 U340 ( .A(n1264), .X(n1287) );
  SEN_INV_S_1 U341 ( .A(n1292), .X(n1295) );
  SEN_OAI21_2 U342 ( .A1(n330), .A2(n1166), .B(n1165), .X(n1187) );
  SEN_MUXI2_S_1 U343 ( .D0(n539), .D1(n538), .S(n340), .X(n546) );
  SEN_MUXI2_D_1 U344 ( .D0(n541), .D1(n537), .S(n341), .X(n538) );
  SEN_ND2_T_2 U345 ( .A1(n758), .A2(n757), .X(n775) );
  SEN_ND2B_1 U346 ( .A(n379), .B(n352), .X(n757) );
  SEN_INV_0P65 U347 ( .A(n405), .X(n236) );
  SEN_INV_0P65 U348 ( .A(n405), .X(n243) );
  SEN_INV_S_1P5 U349 ( .A(n1344), .X(n318) );
  SEN_NR2B_V1DG_1 U350 ( .A(n988), .B(n928), .X(n458) );
  SEN_ND2_G_1 U351 ( .A1(n989), .A2(n988), .X(n990) );
  SEN_INV_S_3 U352 ( .A(n1023), .X(n986) );
  SEN_ND2B_V1_1 U353 ( .A(n357), .B(n386), .X(n1023) );
  SEN_OAI211_4 U354 ( .A1(n1382), .A2(n401), .B1(n250), .B2(n269), .X(n1383)
         );
  SEN_AOI211_2 U355 ( .A1(n413), .A2(n1095), .B1(n1094), .B2(n408), .X(n1099)
         );
  SEN_NR2_0P65 U356 ( .A1(n1093), .A2(n236), .X(n1094) );
  SEN_ND2B_2 U357 ( .A(n976), .B(n1016), .X(n980) );
  SEN_AOAI211_3 U358 ( .A1(n915), .A2(n261), .B(n914), .C(n259), .X(n976) );
  SEN_AOI21B_1 U359 ( .A1(n753), .A2(n734), .B(n751), .X(n328) );
  SEN_ND2_0P8 U360 ( .A1(n752), .A2(n786), .X(n734) );
  SEN_ND2B_V1_2 U361 ( .A(n383), .B(n355), .X(n867) );
  SEN_BUF_6 U362 ( .A(A[12]), .X(n383) );
  SEN_ND2_4 U363 ( .A1(n1369), .A2(n404), .X(n1371) );
  SEN_OAI21_5 U364 ( .A1(n365), .A2(n395), .B(n1185), .X(n1344) );
  SEN_AOAI211_4 U365 ( .A1(n1164), .A2(n1163), .B(n1162), .C(n1161), .X(n1185)
         );
  SEN_AO2BB2_4 U366 ( .A1(n360), .A2(n389), .B1(n1021), .B2(n1072), .X(n1065)
         );
  SEN_AOAI211_G_3 U367 ( .A1(n980), .A2(n981), .B(n979), .C(n978), .X(n1021)
         );
  SEN_BUF_S_3 U368 ( .A(A[14]), .X(n385) );
  SEN_AOI211_3 U369 ( .A1(n1283), .A2(n1310), .B1(n1282), .B2(n1307), .X(n1285) );
  SEN_ND2_T_2 U370 ( .A1(n311), .A2(n1281), .X(n1224) );
  SEN_ND2_1P5 U371 ( .A1(n1310), .A2(n1309), .X(n311) );
  SEN_OR3B_4 U372 ( .B1(n374), .B2(n375), .A(n644), .X(n667) );
  SEN_INV_S_4 U373 ( .A(n599), .X(n644) );
  SEN_MUXI2_S_2 U374 ( .D0(n1275), .D1(n1274), .S(n399), .X(n1276) );
  SEN_OAI21B_1 U375 ( .A1(n986), .A2(n928), .B(n507), .X(n511) );
  SEN_INV_S_2 U376 ( .A(n1228), .X(n1207) );
  SEN_AOI21B_4 U377 ( .A1(n1355), .A2(n1354), .B(n277), .X(n1369) );
  SEN_ND2_S_0P5 U378 ( .A1(n812), .A2(n816), .X(n715) );
  SEN_ND2B_1 U379 ( .A(n350), .B(n377), .X(n812) );
  SEN_NR2_G_2 U380 ( .A1(n654), .A2(n653), .X(n661) );
  SEN_INV_0P65 U381 ( .A(n656), .X(n653) );
  SEN_ND2_2 U382 ( .A1(n631), .A2(n630), .X(n654) );
  SEN_ND2_2 U383 ( .A1(n1344), .A2(n1280), .X(n1309) );
  SEN_AN2_2 U384 ( .A1(n756), .A2(n755), .X(n337) );
  SEN_ND2_0P5 U385 ( .A1(n755), .A2(n777), .X(n719) );
  SEN_ND2B_V1DG_1 U386 ( .A(n351), .B(n378), .X(n755) );
  SEN_AO21B_2 U387 ( .A1(n657), .A2(n656), .B(n655), .X(n659) );
  SEN_ND2B_V1_1 U388 ( .A(n358), .B(n387), .X(n1024) );
  SEN_BUF_AS_3 U389 ( .A(B[16]), .X(n358) );
  SEN_INV_S_1 U390 ( .A(n1273), .X(n1250) );
  SEN_ND2_2 U391 ( .A1(n776), .A2(n775), .X(n807) );
  SEN_INV_S_1 U392 ( .A(n1230), .X(n1209) );
  SEN_ND2_S_4 U393 ( .A1(n1260), .A2(n1261), .X(n1366) );
  SEN_OAI21_T_6 U394 ( .A1(n325), .A2(n1238), .B(n1237), .X(n1260) );
  SEN_OR3B_4 U395 ( .B1(n394), .B2(n395), .A(n1202), .X(n1208) );
  SEN_ND2_S_1 U396 ( .A1(n1271), .A2(n1249), .X(n1275) );
  SEN_MUXI2_S_1 U397 ( .D0(n1232), .D1(n1231), .S(n397), .X(n1233) );
  SEN_OAI221_1 U398 ( .A1(n266), .A2(n1240), .B1(n1230), .B2(n396), .C(n269), 
        .X(n1231) );
  SEN_INV_S_4 U399 ( .A(n528), .X(n1267) );
  SEN_ND2_S_3 U400 ( .A1(n1316), .A2(n1318), .X(n528) );
  SEN_MUXI2_DG_1 U401 ( .D0(n1375), .D1(n1333), .S(n401), .X(n1335) );
  SEN_INV_S_3 U402 ( .A(n1375), .X(n1376) );
  SEN_ND2_S_4 U403 ( .A1(n254), .A2(n1328), .X(n1375) );
  SEN_AO21B_1 U404 ( .A1(n1315), .A2(n1237), .B(n245), .X(n444) );
  SEN_INV_1 U405 ( .A(n239), .X(n259) );
  SEN_BUF_1P5 U406 ( .A(n919), .X(n260) );
  SEN_ND2B_V1_2 U407 ( .A(n816), .B(n817), .X(n1060) );
  SEN_OR2_2 U408 ( .A1(n278), .A2(n279), .X(n1095) );
  SEN_ND3_S_0P5 U409 ( .A1(n655), .A2(n699), .A3(n806), .X(n496) );
  SEN_ND2_T_1 U410 ( .A1(n443), .A2(n334), .X(n450) );
  SEN_ND2_G_1 U411 ( .A1(n913), .A2(n912), .X(n914) );
  SEN_OR2_2 U412 ( .A1(n273), .A2(n274), .X(n648) );
  SEN_ND2_3 U413 ( .A1(n676), .A2(n675), .X(n697) );
  SEN_OR3B_1 U414 ( .B1(n378), .B2(n379), .A(n733), .X(n743) );
  SEN_ND3_T_3 U415 ( .A1(n1060), .A2(n1059), .A3(n247), .X(n1195) );
  SEN_INV_0P65 U416 ( .A(n521), .X(n1221) );
  SEN_AOAI211_0P75 U417 ( .A1(n889), .A2(n293), .B(n888), .C(n259), .X(n898)
         );
  SEN_NR2_T_0P5 U418 ( .A1(n1018), .A2(n885), .X(n889) );
  SEN_OR3B_1 U419 ( .B1(n388), .B2(n389), .A(n1013), .X(n1014) );
  SEN_INV_S_2 U420 ( .A(n1224), .X(n1259) );
  SEN_OAI211_1 U421 ( .A1(n1246), .A2(n402), .B1(n407), .B2(n1245), .X(n1251)
         );
  SEN_ND4_2 U422 ( .A1(n1311), .A2(n1310), .A3(n1338), .A4(n1309), .X(n1313)
         );
  SEN_INV_1P25 U423 ( .A(n404), .X(n402) );
  SEN_MUXI2_D_1 U424 ( .D0(n742), .D1(n266), .S(n353), .X(n745) );
  SEN_AN2_S_2 U425 ( .A1(n1362), .A2(n449), .X(n329) );
  SEN_AO21_1 U426 ( .A1(n776), .A2(n337), .B(n778), .X(n813) );
  SEN_OAI21_3 U427 ( .A1(n350), .A2(n377), .B(n697), .X(n828) );
  SEN_ND2_G_1 U428 ( .A1(n814), .A2(n813), .X(n808) );
  SEN_ND2_0P5 U429 ( .A1(n718), .A2(n820), .X(n786) );
  SEN_AN2_1 U430 ( .A1(n1052), .A2(n1059), .X(n275) );
  SEN_BUF_1P5 U431 ( .A(n943), .X(n261) );
  SEN_OAI21_2 U432 ( .A1(n299), .A2(n1056), .B(n1028), .X(n1051) );
  SEN_NR2_G_2 U433 ( .A1(n286), .A2(n1064), .X(n1078) );
  SEN_ND2B_3 U434 ( .A(n392), .B(n363), .X(n1191) );
  SEN_AOAI211_1 U435 ( .A1(n1357), .A2(n536), .B(n535), .C(n534), .X(n541) );
  SEN_BUF_1P5 U436 ( .A(INST[0]), .X(n340) );
  SEN_BUF_S_1 U437 ( .A(INST[1]), .X(n341) );
  SEN_INV_S_0P5 U438 ( .A(n341), .X(n559) );
  SEN_BUF_S_2 U439 ( .A(n632), .X(n324) );
  SEN_ND2_S_1 U440 ( .A1(n812), .A2(n699), .X(n683) );
  SEN_INV_S_3 U441 ( .A(n701), .X(n733) );
  SEN_ND2_G_0P65 U442 ( .A1(n739), .A2(n738), .X(n741) );
  SEN_OAI21_S_2 U443 ( .A1(n848), .A2(n921), .B(n1053), .X(n850) );
  SEN_AO21B_1 U444 ( .A1(n847), .A2(n911), .B(n944), .X(n852) );
  SEN_BUF_S_2 U445 ( .A(B[15]), .X(n357) );
  SEN_BUF_S_1 U446 ( .A(n1058), .X(n255) );
  SEN_INV_S_0P5 U447 ( .A(n1170), .X(n1063) );
  SEN_OAI211_1 U448 ( .A1(n1309), .A2(n243), .B1(n407), .B2(n1204), .X(n1210)
         );
  SEN_BUF_S_3 U449 ( .A(A[1]), .X(n372) );
  SEN_BUF_4 U450 ( .A(A[3]), .X(n374) );
  SEN_BUF_2 U451 ( .A(A[4]), .X(n375) );
  SEN_BUF_1P5 U452 ( .A(B[4]), .X(n348) );
  SEN_BUF_S_4 U453 ( .A(A[7]), .X(n378) );
  SEN_BUF_S_3 U454 ( .A(B[12]), .X(n355) );
  SEN_OR2_DG_1 U455 ( .A1(n893), .A2(n402), .X(n283) );
  SEN_BUF_S_4 U456 ( .A(A[15]), .X(n386) );
  SEN_BUF_1P5 U457 ( .A(A[16]), .X(n387) );
  SEN_MUXI2_D_1 U458 ( .D0(n958), .D1(n963), .S(n359), .X(n959) );
  SEN_BUF_1P5 U459 ( .A(A[17]), .X(n388) );
  SEN_BUF_1P5 U460 ( .A(B[17]), .X(n359) );
  SEN_BUF_S_1 U461 ( .A(A[18]), .X(n389) );
  SEN_BUF_1P5 U462 ( .A(A[20]), .X(n391) );
  SEN_MUXI2_S_0P5 U463 ( .D0(n1210), .D1(n1379), .S(n366), .X(n1211) );
  SEN_ND2_2 U464 ( .A1(n1298), .A2(n1302), .X(n251) );
  SEN_ND2B_S_1 U465 ( .A(n745), .B(n744), .X(n746) );
  SEN_ND2_S_1 U466 ( .A1(n1107), .A2(n1106), .X(Z[21]) );
  SEN_ND2_S_0P5 U467 ( .A1(n1151), .A2(n1150), .X(n1152) );
  SEN_ND3_S_0P5 U468 ( .A1(n1235), .A2(n1234), .A3(n1233), .X(Z[26]) );
  SEN_MUXI2_DG_3 U469 ( .D0(n1254), .D1(n1253), .S(n398), .X(n1255) );
  SEN_AOAI211_3 U470 ( .A1(n1259), .A2(n1346), .B(n1304), .C(n1306), .X(n1263)
         );
  SEN_INV_S_2 U471 ( .A(n1263), .X(n1266) );
  SEN_OAI211_2 U472 ( .A1(n1263), .A2(n242), .B1(n1262), .B2(n407), .X(n1269)
         );
  SEN_MUXI2_S_1 U473 ( .D0(n1146), .D1(n1149), .S(n364), .X(n1147) );
  SEN_MUXI2_DG_1 U474 ( .D0(n546), .D1(n545), .S(n342), .X(n566) );
  SEN_AOI221_0P5 U475 ( .A1(B[22]), .A2(n393), .B1(n1136), .B2(n1135), .C(
        n1134), .X(n237) );
  SEN_NR3B_4 U476 ( .A(n1135), .B1(n1133), .B2(n1132), .X(n1134) );
  SEN_AOAI211_1 U477 ( .A1(n1114), .A2(n1113), .B(n1132), .C(n1112), .X(n1136)
         );
  SEN_OAI21_G_0P5 U478 ( .A1(n996), .A2(n1027), .B(n995), .X(n998) );
  SEN_OAI21_0P75 U479 ( .A1(n1219), .A2(n236), .B(n1201), .X(n1205) );
  SEN_MUXI2_S_0P5 U480 ( .D0(n1205), .D1(n1210), .S(n366), .X(n1206) );
  SEN_AN3B_0P5 U481 ( .B1(n1072), .B2(n1017), .A(n238), .X(n1019) );
  SEN_NR3_T_0P5 U482 ( .A1(n864), .A2(n1067), .A3(n238), .X(n865) );
  SEN_INV_S_0P5 U483 ( .A(n238), .X(n293) );
  SEN_NR2_S_0P65 U484 ( .A1(n829), .A2(n828), .X(n238) );
  SEN_MUXI2_S_0P5 U485 ( .D0(n1003), .D1(n1002), .S(n1001), .X(n1012) );
  SEN_OAI22_T_0P5 U486 ( .A1(n242), .A2(n997), .B1(n998), .B2(n410), .X(n1003)
         );
  SEN_BUF_1P5 U487 ( .A(n244), .X(n405) );
  SEN_INV_S_0P5 U488 ( .A(n405), .X(n242) );
  SEN_AN2_S_0P5 U489 ( .A1(n385), .A2(B[14]), .X(n239) );
  SEN_BUF_S_1 U490 ( .A(n244), .X(n404) );
  SEN_AN2_1 U491 ( .A1(n309), .A2(n310), .X(n240) );
  SEN_INV_2 U492 ( .A(n1309), .X(n1219) );
  SEN_ND2_4 U493 ( .A1(n817), .A2(n815), .X(n1059) );
  SEN_OAI21_G_1 U494 ( .A1(n1029), .A2(n1051), .B(n255), .X(n1031) );
  SEN_NR3_T_0P65 U495 ( .A1(n1026), .A2(n1054), .A3(n1025), .X(n1029) );
  SEN_INV_1 U496 ( .A(n854), .X(n855) );
  SEN_ND2_0P5 U497 ( .A1(n863), .A2(n862), .X(Z[13]) );
  SEN_INV_S_1 U498 ( .A(n413), .X(n411) );
  SEN_ND2_S_0P65 U499 ( .A1(n389), .A2(n360), .X(n1071) );
  SEN_NR2B_V1_4 U500 ( .A(n1071), .B(n285), .X(n286) );
  SEN_ND2_S_0P8 U501 ( .A1(n1242), .A2(n1241), .X(n1247) );
  SEN_AOAI211_1 U502 ( .A1(n338), .A2(n1256), .B(n1258), .C(n1255), .X(Z[27])
         );
  SEN_BUF_1 U503 ( .A(n1065), .X(n241) );
  SEN_ND2_S_0P65 U504 ( .A1(n351), .A2(n378), .X(n752) );
  SEN_AOAI211_0P75 U505 ( .A1(n338), .A2(n908), .B(n910), .C(n907), .X(Z[15])
         );
  SEN_MUXI2_DG_1 U506 ( .D0(n906), .D1(n905), .S(n386), .X(n907) );
  SEN_NR2_1 U507 ( .A1(n1091), .A2(n1171), .X(n278) );
  SEN_OAI22_S_1 U508 ( .A1(n1092), .A2(n402), .B1(n1095), .B2(n409), .X(n1105)
         );
  SEN_AOAI211_G_4 U509 ( .A1(n263), .A2(n921), .B(n920), .C(n260), .X(n987) );
  SEN_INV_1 U510 ( .A(n1194), .X(n1196) );
  SEN_NR2_S_0P65 U511 ( .A1(n374), .A2(n347), .X(n273) );
  SEN_ND3_T_2 U512 ( .A1(n473), .A2(n472), .A3(n471), .X(n537) );
  SEN_ND2B_V1DG_1 U513 ( .A(n858), .B(n857), .X(n859) );
  SEN_NR3_T_0P5 U514 ( .A1(n1069), .A2(n1068), .A3(n1067), .X(n1076) );
  SEN_INV_S_1P5 U515 ( .A(n302), .X(n303) );
  SEN_INV_S_0P5 U516 ( .A(n1000), .X(n997) );
  SEN_OAI21_G_0P5 U517 ( .A1(n982), .A2(n248), .B(n1072), .X(n1000) );
  SEN_ND2_T_0P5 U518 ( .A1(n819), .A2(n246), .X(n824) );
  SEN_AN2_DG_1 U519 ( .A1(n820), .A2(n818), .X(n246) );
  SEN_AOAI211_0P75 U520 ( .A1(n1366), .A2(n1360), .B(n1356), .C(n1361), .X(
        n1322) );
  SEN_MUXI2_DG_3 U521 ( .D0(n1327), .D1(n1326), .S(n1325), .X(n1336) );
  SEN_BUF_S_4 U522 ( .A(A[8]), .X(n379) );
  SEN_OR2_2 U523 ( .A1(n320), .A2(n321), .X(n779) );
  SEN_OR3B_2 U524 ( .B1(n390), .B2(n391), .A(n1088), .X(n1100) );
  SEN_OAI22_1 U525 ( .A1(n954), .A2(n236), .B1(n956), .B2(n410), .X(n958) );
  SEN_AOAI211_1 U526 ( .A1(n338), .A2(n970), .B(n969), .C(n968), .X(Z[17]) );
  SEN_BUF_1P5 U527 ( .A(A[28]), .X(n399) );
  SEN_INV_0P5 U528 ( .A(n467), .X(n469) );
  SEN_ND2B_1 U529 ( .A(n1102), .B(n1101), .X(n1103) );
  SEN_MUXI2_S_2 U530 ( .D0(n1104), .D1(n1103), .S(n392), .X(n1107) );
  SEN_ND2_0P5 U531 ( .A1(n383), .A2(n355), .X(n944) );
  SEN_ND3_S_4 U532 ( .A1(n287), .A2(n288), .A3(n406), .X(n963) );
  SEN_OR2_1 U533 ( .A1(n957), .A2(n402), .X(n287) );
  SEN_OR2_1 U534 ( .A1(n276), .A2(n411), .X(n288) );
  SEN_INV_4 U535 ( .A(n1368), .X(n1373) );
  SEN_INV_0P65 U536 ( .A(n414), .X(n410) );
  SEN_BUF_1 U537 ( .A(n416), .X(n414) );
  SEN_NR2B_V1_1 U538 ( .A(n1052), .B(n832), .X(n475) );
  SEN_ND2_S_0P8 U539 ( .A1(n1053), .A2(n867), .X(n832) );
  SEN_AOAI211_1 U540 ( .A1(n532), .A2(n531), .B(n530), .C(n529), .X(n536) );
  SEN_AOAI211_1 U541 ( .A1(n527), .A2(n526), .B(n525), .C(n524), .X(n532) );
  SEN_ND2B_V1DG_1 U542 ( .A(B[26]), .B(n397), .X(n1237) );
  SEN_NR2_S_1 U543 ( .A1(n1221), .A2(n522), .X(n441) );
  SEN_INV_0P65 U544 ( .A(n569), .X(n587) );
  SEN_ND2_S_1 U545 ( .A1(n371), .A2(n344), .X(n569) );
  SEN_INV_3 U546 ( .A(n808), .X(n810) );
  SEN_INV_S_1P5 U547 ( .A(n647), .X(n645) );
  SEN_ND2_0P65 U548 ( .A1(n347), .A2(n374), .X(n647) );
  SEN_MUXI2_D_1 U549 ( .D0(n1105), .D1(n1096), .S(n363), .X(n1097) );
  SEN_ND2_G_1 U550 ( .A1(n877), .A2(n853), .X(n860) );
  SEN_MUXI2_S_1 U551 ( .D0(n1247), .D1(n1251), .S(n367), .X(n1248) );
  SEN_INV_1 U552 ( .A(n1322), .X(n1320) );
  SEN_OAI22_S_1 U553 ( .A1(n1323), .A2(n242), .B1(n1322), .B2(n409), .X(n1326)
         );
  SEN_MUXI2_DG_1 U554 ( .D0(n1298), .D1(n1292), .S(n400), .X(n1303) );
  SEN_OAI211_1 U555 ( .A1(n1273), .A2(n398), .B1(n269), .B2(n1272), .X(n1274)
         );
  SEN_OAI221_1 U556 ( .A1(n606), .A2(n403), .B1(n605), .B2(n410), .C(n406), 
        .X(n608) );
  SEN_INV_0P65 U557 ( .A(n408), .X(n406) );
  SEN_MUXI2_D_1 U558 ( .D0(n544), .D1(n543), .S(n542), .X(n545) );
  SEN_ND2_T_0P5 U559 ( .A1(n658), .A2(n655), .X(n486) );
  SEN_ND2B_V1DG_1 U560 ( .A(n348), .B(n375), .X(n658) );
  SEN_ND2_2 U561 ( .A1(n568), .A2(n494), .X(n660) );
  SEN_ND2B_V1_1 U562 ( .A(n371), .B(n344), .X(n568) );
  SEN_OAI22_S_1 U563 ( .A1(n1030), .A2(n402), .B1(n1031), .B2(n410), .X(n1042)
         );
  SEN_OAI221_2 U564 ( .A1(n1033), .A2(n403), .B1(n1032), .B2(n410), .C(n406), 
        .X(n1036) );
  SEN_INV_0P8 U565 ( .A(n1031), .X(n1032) );
  SEN_AO2BB2_4 U566 ( .A1(n348), .A2(n375), .B1(n648), .B2(n647), .X(n650) );
  SEN_ND2_4 U567 ( .A1(n784), .A2(n783), .X(n826) );
  SEN_INV_S_4 U568 ( .A(n787), .X(n784) );
  SEN_OAI22_T_0P5 U569 ( .A1(n849), .A2(n243), .B1(n850), .B2(n410), .X(n861)
         );
  SEN_ND2_G_1 U570 ( .A1(n255), .A2(n1028), .X(n1001) );
  SEN_MUXI2_D_1 U571 ( .D0(n855), .D1(n266), .S(n356), .X(n858) );
  SEN_OAI21_G_2 U572 ( .A1(n736), .A2(n735), .B(n756), .X(n737) );
  SEN_INV_1P5 U573 ( .A(n719), .X(n736) );
  SEN_MUXI2_S_1 U574 ( .D0(n1149), .D1(n1379), .S(n364), .X(n1150) );
  SEN_ND2_S_1P5 U575 ( .A1(n1098), .A2(n1097), .X(n1104) );
  SEN_ND2_T_2 U576 ( .A1(n699), .A2(n698), .X(n816) );
  SEN_ND2B_1 U577 ( .A(n377), .B(n350), .X(n699) );
  SEN_MUXI2_DG_0P75 U578 ( .D0(n1099), .D1(n266), .S(n363), .X(n1102) );
  SEN_OR2_5 U579 ( .A1(n313), .A2(n314), .X(n1298) );
  SEN_ND2_S_1 U580 ( .A1(n630), .A2(n660), .X(n601) );
  SEN_OAI221_1 U581 ( .A1(n793), .A2(n403), .B1(n792), .B2(n410), .C(n406), 
        .X(n797) );
  SEN_INV_S_1 U582 ( .A(n791), .X(n792) );
  SEN_ND2B_V1_1 U583 ( .A(n354), .B(n382), .X(n1052) );
  SEN_ND2_G_1 U584 ( .A1(n1192), .A2(n1194), .X(n1170) );
  SEN_ND2_T_1 U585 ( .A1(n904), .A2(n903), .X(n905) );
  SEN_ND2_2 U586 ( .A1(n965), .A2(n964), .X(n966) );
  SEN_MUXI2_S_3 U587 ( .D0(n963), .D1(n1379), .S(n359), .X(n964) );
  SEN_MUXI2_S_3 U588 ( .D0(n1041), .D1(n1040), .S(n390), .X(n1044) );
  SEN_MUXI2_S_1 U589 ( .D0(n1042), .D1(n1036), .S(n361), .X(n1034) );
  SEN_AOAI211_G_2 U590 ( .A1(n1344), .A2(n1345), .B(n1341), .C(n1346), .X(
        n1246) );
  SEN_ND2B_S_0P5 U591 ( .A(n401), .B(B[30]), .X(n1357) );
  SEN_BUF_S_1 U592 ( .A(A[30]), .X(n401) );
  SEN_ND2B_V1_1 U593 ( .A(n402), .B(n1246), .X(n1241) );
  SEN_INV_S_4 U594 ( .A(n1014), .X(n1088) );
  SEN_ND2_S_3 U595 ( .A1(n918), .A2(n917), .X(n920) );
  SEN_ND2B_1 U596 ( .A(n384), .B(n356), .X(n917) );
  SEN_NR2_S_0P5 U597 ( .A1(n678), .A2(n683), .X(n425) );
  SEN_NR2B_V1_2 U598 ( .A(n677), .B(n683), .X(n487) );
  SEN_INV_1 U599 ( .A(n1033), .X(n1030) );
  SEN_OAI21_0P75 U600 ( .A1(n1022), .A2(n241), .B(n1071), .X(n1033) );
  SEN_ND2_2 U601 ( .A1(n633), .A2(n324), .X(n657) );
  SEN_ND2B_V1_1 U602 ( .A(n345), .B(n372), .X(n630) );
  SEN_OAI22_0P5 U603 ( .A1(n702), .A2(n243), .B1(n715), .B2(n409), .X(n705) );
  SEN_ND2_G_1 U604 ( .A1(n806), .A2(n715), .X(n777) );
  SEN_AOI211_G_1 U605 ( .A1(n1108), .A2(n1110), .B1(n467), .B2(n466), .X(n468)
         );
  SEN_ND2B_S_0P5 U606 ( .A(B[22]), .B(n393), .X(n1138) );
  SEN_ND2B_V1_2 U607 ( .A(n368), .B(n399), .X(n1316) );
  SEN_OR3B_2 U608 ( .B1(n392), .B2(n393), .A(n1142), .X(n1143) );
  SEN_BUF_S_1 U609 ( .A(B[23]), .X(n364) );
  SEN_INV_S_0P5 U610 ( .A(n1329), .X(n1379) );
  SEN_BUF_S_4 U611 ( .A(B[9]), .X(n353) );
  SEN_NR2_S_2 U612 ( .A1(n1289), .A2(n403), .X(n313) );
  SEN_INV_S_0P5 U613 ( .A(n510), .X(n505) );
  SEN_NR2_S_0P5 U614 ( .A1(n485), .A2(n484), .X(n503) );
  SEN_AOAI211_1 U615 ( .A1(n512), .A2(n511), .B(n510), .C(n509), .X(n514) );
  SEN_ND2_S_0P5 U616 ( .A1(n1167), .A2(n1168), .X(n1188) );
  SEN_INV_1 U617 ( .A(n333), .X(n334) );
  SEN_ND2_G_1 U618 ( .A1(n444), .A2(n442), .X(n333) );
  SEN_ND2_S_0P5 U619 ( .A1(n354), .A2(n382), .X(n1066) );
  SEN_INV_S_0P5 U620 ( .A(n822), .X(n823) );
  SEN_ND2B_S_1 U621 ( .A(n353), .B(n380), .X(n776) );
  SEN_ND2B_V1DG_1 U622 ( .A(B[10]), .B(n381), .X(n814) );
  SEN_ND2_G_1 U623 ( .A1(n805), .A2(n807), .X(n778) );
  SEN_OR2_1 U624 ( .A1(n383), .A2(n355), .X(n911) );
  SEN_ND2B_S_1 U625 ( .A(n355), .B(n383), .X(n1053) );
  SEN_INV_S_0P5 U626 ( .A(n1168), .X(n1139) );
  SEN_ND2B_1 U627 ( .A(n399), .B(n368), .X(n1318) );
  SEN_INV_S_0P5 U628 ( .A(n340), .X(n551) );
  SEN_INV_S_0P5 U629 ( .A(n1110), .X(n279) );
  SEN_BUF_S_1 U630 ( .A(B[25]), .X(n366) );
  SEN_BUF_S_1 U631 ( .A(n1260), .X(n272) );
  SEN_BUF_AS_0P5 U632 ( .A(n422), .X(n419) );
  SEN_INV_0P65 U633 ( .A(n1370), .X(n408) );
  SEN_BUF_S_4 U634 ( .A(A[9]), .X(n380) );
  SEN_INV_S_1 U635 ( .A(n741), .X(n742) );
  SEN_BUF_S_2 U636 ( .A(B[21]), .X(n363) );
  SEN_BUF_S_1 U637 ( .A(A[23]), .X(n394) );
  SEN_NR2_S_0P5 U638 ( .A1(n1148), .A2(n1332), .X(n1151) );
  SEN_INV_0P5 U639 ( .A(n1158), .X(n1148) );
  SEN_BUF_S_1 U640 ( .A(A[24]), .X(n395) );
  SEN_BUF_S_1 U641 ( .A(B[24]), .X(n365) );
  SEN_ND2_2 U642 ( .A1(n316), .A2(n1290), .X(n1292) );
  SEN_ND2_2 U643 ( .A1(n405), .A2(n1289), .X(n1290) );
  SEN_BUF_S_1 U644 ( .A(A[29]), .X(n400) );
  SEN_NR2_0P65 U645 ( .A1(n474), .A2(n762), .X(n478) );
  SEN_ND2_S_0P5 U646 ( .A1(n495), .A2(n655), .X(n488) );
  SEN_NR2B_V1_1 U647 ( .A(n755), .B(n489), .X(n493) );
  SEN_INV_S_0P5 U648 ( .A(n776), .X(n474) );
  SEN_NR2_S_0P5 U649 ( .A1(n445), .A2(n1358), .X(n442) );
  SEN_ND3_1 U650 ( .A1(n450), .A2(n448), .A3(n447), .X(n449) );
  SEN_OAI21_0P75 U651 ( .A1(n520), .A2(n1188), .B(n519), .X(n527) );
  SEN_ND2B_V1DG_1 U652 ( .A(n381), .B(n780), .X(n818) );
  SEN_ND2_0P5 U653 ( .A1(n717), .A2(n716), .X(n820) );
  SEN_ND2_S_0P5 U654 ( .A1(n910), .A2(n909), .X(n974) );
  SEN_ND2_S_0P5 U655 ( .A1(n1016), .A2(n1015), .X(n1070) );
  SEN_ND2_G_1 U656 ( .A1(n255), .A2(n1051), .X(n1194) );
  SEN_ND2B_S_0P5 U657 ( .A(n390), .B(n361), .X(n1192) );
  SEN_AOAI211_0P5 U658 ( .A1(n439), .A2(n438), .B(n437), .C(n952), .X(n459) );
  SEN_AOAI211_0P5 U659 ( .A1(n436), .A2(n435), .B(n434), .C(n433), .X(n439) );
  SEN_ND2_S_0P5 U660 ( .A1(n373), .A2(n346), .X(n625) );
  SEN_ND2B_V1DG_1 U661 ( .A(n375), .B(n348), .X(n655) );
  SEN_ND2B_V1DG_1 U662 ( .A(n347), .B(n374), .X(n656) );
  SEN_AO21B_1 U663 ( .A1(n598), .A2(n588), .B(n587), .X(n651) );
  SEN_INV_S_0P5 U664 ( .A(n495), .X(n678) );
  SEN_INV_0P8 U665 ( .A(n781), .X(n257) );
  SEN_ND2B_V1DG_1 U666 ( .A(n381), .B(B[10]), .X(n805) );
  SEN_INV_S_1P5 U667 ( .A(n790), .X(n846) );
  SEN_INV_S_0P5 U668 ( .A(n944), .X(n1067) );
  SEN_AOI31_1 U669 ( .A1(n827), .A2(n826), .A3(n825), .B(n829), .X(n1073) );
  SEN_ND2_T_0P5 U670 ( .A1(n356), .A2(n384), .X(n943) );
  SEN_OR2_DG_1 U671 ( .A1(n387), .A2(n358), .X(n975) );
  SEN_NR2_T_1 U672 ( .A1(n991), .A2(n990), .X(n994) );
  SEN_INV_S_0P5 U673 ( .A(n995), .X(n1056) );
  SEN_ND2_0P65 U674 ( .A1(n1053), .A2(n275), .X(n1025) );
  SEN_ND2_G_1 U675 ( .A1(n942), .A2(n944), .X(n1018) );
  SEN_ND2B_S_2 U676 ( .A(n391), .B(n362), .X(n1193) );
  SEN_ND2B_S_1 U677 ( .A(n361), .B(n390), .X(n1109) );
  SEN_ND2B_V1DG_1 U678 ( .A(n362), .B(n391), .X(n1110) );
  SEN_ND2B_1 U679 ( .A(n393), .B(B[22]), .X(n1168) );
  SEN_INV_S_0P5 U680 ( .A(n1193), .X(n1171) );
  SEN_ND2B_S_0P5 U681 ( .A(B[30]), .B(n401), .X(n1362) );
  SEN_BUF_S_3 U682 ( .A(A[0]), .X(n371) );
  SEN_BUF_1P5 U683 ( .A(B[0]), .X(n344) );
  SEN_BUF_1P5 U684 ( .A(B[1]), .X(n345) );
  SEN_ND2B_V1DG_1 U685 ( .A(n373), .B(n346), .X(n632) );
  SEN_ND2_1P5 U686 ( .A1(n307), .A2(n677), .X(n698) );
  SEN_INV_S_0P5 U687 ( .A(n678), .X(n306) );
  SEN_BUF_S_3 U688 ( .A(B[7]), .X(n351) );
  SEN_INV_S_3 U689 ( .A(n743), .X(n789) );
  SEN_INV_S_0P5 U690 ( .A(B[10]), .X(n780) );
  SEN_ND2_0P8 U691 ( .A1(n814), .A2(n805), .X(n762) );
  SEN_OAI221_1 U692 ( .A1(n852), .A2(n402), .B1(n851), .B2(n411), .C(n406), 
        .X(n854) );
  SEN_INV_S_0P5 U693 ( .A(n850), .X(n851) );
  SEN_INV_S_0P5 U694 ( .A(B[14]), .X(n886) );
  SEN_ND2_S_0P5 U695 ( .A1(n260), .A2(n918), .X(n490) );
  SEN_NR2_S_1 U696 ( .A1(n985), .A2(n949), .X(n953) );
  SEN_INV_S_0P5 U697 ( .A(n1081), .X(n1091) );
  SEN_ND2_T_0P5 U698 ( .A1(n1109), .A2(n1140), .X(n1081) );
  SEN_OAI21_0P75 U699 ( .A1(n1090), .A2(n1089), .B(n1113), .X(n1093) );
  SEN_INV_S_2 U700 ( .A(n1100), .X(n1142) );
  SEN_ND2B_S_0P5 U701 ( .A(n1100), .B(n420), .X(n1125) );
  SEN_ND2_S_0P5 U702 ( .A1(n1237), .A2(n523), .X(n522) );
  SEN_ND2_S_0P5 U703 ( .A1(n1362), .A2(n1357), .X(n1324) );
  SEN_AOI211_0P5 U704 ( .A1(n1341), .A2(n1346), .B1(n1340), .B2(n1339), .X(
        n1355) );
  SEN_BUF_S_1 U705 ( .A(INST[2]), .X(n342) );
  SEN_BUF_S_3 U706 ( .A(B[2]), .X(n346) );
  SEN_BUF_S_2 U707 ( .A(B[3]), .X(n347) );
  SEN_BUF_S_1 U708 ( .A(B[5]), .X(n349) );
  SEN_BUF_1P5 U709 ( .A(A[5]), .X(n376) );
  SEN_BUF_1P5 U710 ( .A(A[6]), .X(n377) );
  SEN_BUF_S_1 U711 ( .A(B[6]), .X(n350) );
  SEN_MUXI2_S_0P5 U712 ( .D0(n705), .D1(n708), .S(n351), .X(n706) );
  SEN_BUF_1P5 U713 ( .A(A[10]), .X(n381) );
  SEN_BUF_S_1 U714 ( .A(A[11]), .X(n382) );
  SEN_BUF_S_1 U715 ( .A(B[11]), .X(n354) );
  SEN_BUF_S_3 U716 ( .A(B[13]), .X(n356) );
  SEN_BUF_S_4 U717 ( .A(A[13]), .X(n384) );
  SEN_ND2B_S_0P5 U718 ( .A(n412), .B(n926), .X(n924) );
  SEN_OAI22_S_0P5 U719 ( .A1(n242), .A2(n927), .B1(n926), .B2(n410), .X(n930)
         );
  SEN_INV_S_0P5 U720 ( .A(n925), .X(n927) );
  SEN_BUF_S_1 U721 ( .A(B[18]), .X(n360) );
  SEN_BUF_S_1 U722 ( .A(B[19]), .X(n361) );
  SEN_BUF_S_1 U723 ( .A(A[19]), .X(n390) );
  SEN_BUF_1P5 U724 ( .A(B[20]), .X(n362) );
  SEN_BUF_S_2 U725 ( .A(A[21]), .X(n392) );
  SEN_BUF_S_1 U726 ( .A(A[22]), .X(n393) );
  SEN_ND3_S_0P5 U727 ( .A1(n1117), .A2(n1116), .A3(n406), .X(n1122) );
  SEN_BUF_S_1 U728 ( .A(A[25]), .X(n396) );
  SEN_ND2_S_0P65 U729 ( .A1(n1207), .A2(n1206), .X(n1214) );
  SEN_ND2_S_0P5 U730 ( .A1(n415), .A2(n1236), .X(n1223) );
  SEN_OAI22_0P75 U731 ( .A1(n1236), .A2(n410), .B1(n1259), .B2(n242), .X(n1226) );
  SEN_BUF_S_1 U732 ( .A(A[26]), .X(n397) );
  SEN_BUF_S_3 U733 ( .A(A[27]), .X(n398) );
  SEN_OAI21_2 U734 ( .A1(n242), .A2(n1266), .B(n1265), .X(n1268) );
  SEN_BUF_S_1 U735 ( .A(B[28]), .X(n368) );
  SEN_OR3B_0P5 U736 ( .B1(n1332), .B2(n1331), .A(n1382), .X(n1333) );
  SEN_ND3_S_0P5 U737 ( .A1(n643), .A2(n642), .A3(n641), .X(Z[4]) );
  SEN_ND2_S_0P5 U738 ( .A1(n348), .A2(n267), .X(n641) );
  SEN_AOAI211_0P5 U739 ( .A1(n380), .A2(n748), .B(n267), .C(n353), .X(n749) );
  SEN_ND2_S_0P5 U740 ( .A1(n386), .A2(n899), .X(n908) );
  SEN_MUXI2_D_1 U741 ( .D0(n967), .D1(n966), .S(n388), .X(n968) );
  SEN_ND3_S_0P5 U742 ( .A1(n1184), .A2(n1183), .A3(n1182), .X(Z[24]) );
  SEN_ND2_T_2 U743 ( .A1(n1077), .A2(n1078), .X(n1133) );
  SEN_MUXI2_S_0P5 U744 ( .D0(n1227), .D1(n1226), .S(n1225), .X(n1235) );
  SEN_BUF_S_1 U745 ( .A(B[29]), .X(n369) );
  SEN_INV_0P65 U746 ( .A(n601), .X(n498) );
  SEN_BUF_S_1 U747 ( .A(B[27]), .X(n367) );
  SEN_AN2_S_0P5 U748 ( .A1(n335), .A2(n336), .X(n244) );
  SEN_AN2_S_0P5 U749 ( .A1(n1267), .A2(n1261), .X(n245) );
  SEN_INV_1P25 U750 ( .A(n628), .X(n274) );
  SEN_BUF_S_1 U751 ( .A(INST[3]), .X(n343) );
  SEN_INV_S_0P5 U752 ( .A(n343), .X(n565) );
  SEN_AN2_S_0P5 U753 ( .A1(n1062), .A2(n1061), .X(n247) );
  SEN_ND2B_V1DG_1 U754 ( .A(n385), .B(B[14]), .X(n918) );
  SEN_INV_S_0P5 U755 ( .A(n663), .X(n679) );
  SEN_AOI21B_0P5 U756 ( .A1(n244), .A2(n328), .B(n407), .X(n739) );
  SEN_AOAI211_0P5 U757 ( .A1(n981), .A2(n980), .B(n979), .C(n978), .X(n248) );
  SEN_AO31_2 U758 ( .A1(n827), .A2(n826), .A3(n825), .B(n829), .X(n249) );
  SEN_AN2_S_4 U759 ( .A1(n297), .A2(n298), .X(n250) );
  SEN_ND2_2 U760 ( .A1(n1380), .A2(n296), .X(n297) );
  SEN_OR3B_2 U761 ( .B1(n373), .B2(n371), .A(n598), .X(n599) );
  SEN_OR3B_2 U762 ( .B1(n380), .B2(n381), .A(n789), .X(n790) );
  SEN_OAI211_0P5 U763 ( .A1(n925), .A2(n402), .B1(n924), .B2(n407), .X(n931)
         );
  SEN_MUXI2_DG_3 U764 ( .D0(n1386), .D1(n1380), .S(n370), .X(n1378) );
  SEN_ND2_0P8 U765 ( .A1(n960), .A2(n959), .X(n967) );
  SEN_AN2_S_4 U766 ( .A1(n331), .A2(n1294), .X(n254) );
  SEN_ND2_4 U767 ( .A1(n1200), .A2(n1199), .X(n1203) );
  SEN_OR4B_4 U768 ( .B1(n1198), .B2(n1197), .B3(n1196), .A(n1195), .X(n1199)
         );
  SEN_INV_0P65 U769 ( .A(n911), .X(n915) );
  SEN_INV_S_0P5 U770 ( .A(n1270), .X(n1249) );
  SEN_ND3_T_2 U771 ( .A1(n1074), .A2(n249), .A3(n303), .X(n1077) );
  SEN_AOI211_G_2 U772 ( .A1(n499), .A2(n498), .B1(n497), .B2(n496), .X(n500)
         );
  SEN_NR2_T_2 U773 ( .A1(n987), .A2(n986), .X(n991) );
  SEN_ND2_T_2 U774 ( .A1(n1376), .A2(n253), .X(n1384) );
  SEN_AN3B_1 U775 ( .B1(n263), .B2(n1052), .A(n490), .X(n491) );
  SEN_ND2B_V1DG_1 U776 ( .A(n352), .B(n379), .X(n756) );
  SEN_ND3_T_0P5 U777 ( .A1(n944), .A2(n261), .A3(n942), .X(n973) );
  SEN_ND2_T_0P5 U778 ( .A1(n357), .A2(n386), .X(n1016) );
  SEN_INV_S_2 U779 ( .A(n864), .X(n942) );
  SEN_ND2B_1 U780 ( .A(n349), .B(n376), .X(n677) );
  SEN_NR2B_V1_1 U781 ( .A(n758), .B(n762), .X(n435) );
  SEN_ND2B_V1DG_1 U782 ( .A(n380), .B(n353), .X(n758) );
  SEN_ND2B_V1DG_1 U783 ( .A(n1073), .B(n1066), .X(n864) );
  SEN_ND2_T_1 U784 ( .A1(n631), .A2(n324), .X(n592) );
  SEN_AOAI211_3 U785 ( .A1(n1314), .A2(n1313), .B(n1337), .C(n1352), .X(n1321)
         );
  SEN_ND3_T_2 U786 ( .A1(n1278), .A2(n1277), .A3(n1276), .X(Z[28]) );
  SEN_ND2B_V1DG_2 U787 ( .A(n412), .B(n1291), .X(n1288) );
  SEN_ND2B_V1DG_1 U788 ( .A(n387), .B(n358), .X(n989) );
  SEN_ND2B_V1DG_1 U789 ( .A(n385), .B(n886), .X(n913) );
  SEN_INV_S_4 U790 ( .A(n667), .X(n700) );
  SEN_ND2_2 U791 ( .A1(n1251), .A2(n1258), .X(n309) );
  SEN_INV_S_2 U792 ( .A(n922), .X(n262) );
  SEN_INV_4 U793 ( .A(n262), .X(n263) );
  SEN_AOAI211_0P75 U794 ( .A1(n390), .A2(n1042), .B(n267), .C(n361), .X(n1043)
         );
  SEN_ND2_S_0P5 U795 ( .A1(n261), .A2(n259), .X(n1068) );
  SEN_INV_S_0P5 U796 ( .A(n339), .X(n264) );
  SEN_INV_S_0P5 U797 ( .A(n1329), .X(n265) );
  SEN_INV_S_0P5 U798 ( .A(n265), .X(n266) );
  SEN_AN2_S_0P5 U799 ( .A1(n547), .A2(n551), .X(n335) );
  SEN_INV_S_0P5 U800 ( .A(n338), .X(n267) );
  SEN_INV_S_0P5 U801 ( .A(n1381), .X(n268) );
  SEN_INV_S_0P5 U802 ( .A(n268), .X(n269) );
  SEN_OAI211_4 U803 ( .A1(n1373), .A2(n411), .B1(n1371), .B2(n407), .X(n1380)
         );
  SEN_MUXI2_D_1 U804 ( .D0(n551), .D1(n559), .S(n540), .X(n543) );
  SEN_NR2_S_0P5 U805 ( .A1(n455), .A2(n454), .X(n270) );
  SEN_INV_S_0P5 U806 ( .A(n270), .X(n271) );
  SEN_OA21_2 U807 ( .A1(n994), .A2(n993), .B(n992), .X(n299) );
  SEN_AO21B_6 U808 ( .A1(n824), .A2(n312), .B(n823), .X(n829) );
  SEN_ND2_2 U809 ( .A1(n1296), .A2(n421), .X(n331) );
  SEN_INV_0P65 U810 ( .A(n1321), .X(n1323) );
  SEN_AN4B_1 U811 ( .B1(n1191), .B2(n505), .B3(n1193), .A(n504), .X(n516) );
  SEN_INV_1 U812 ( .A(n541), .X(n542) );
  SEN_INV_1 U813 ( .A(n830), .X(n848) );
  SEN_AOA211_DG_1 U814 ( .A1(n953), .A2(n952), .B(n951), .C(n1024), .X(n276)
         );
  SEN_AOA211_DG_1 U815 ( .A1(n1353), .A2(n1352), .B(n1351), .C(n1350), .X(n277) );
  SEN_OR2_DG_1 U816 ( .A1(n328), .A2(n402), .X(n280) );
  SEN_OR2_1 U817 ( .A1(n737), .A2(n409), .X(n281) );
  SEN_ND2_2 U818 ( .A1(n280), .A2(n281), .X(n748) );
  SEN_INV_S_0P5 U819 ( .A(n414), .X(n409) );
  SEN_MUXI2_DG_3 U820 ( .D0(n1269), .D1(n1268), .S(n1267), .X(n1278) );
  SEN_BUF_1 U821 ( .A(n1185), .X(n282) );
  SEN_MUXI2_DG_3 U822 ( .D0(n1384), .D1(n1383), .S(A[31]), .X(n1388) );
  SEN_OR2_1 U823 ( .A1(n896), .A2(n409), .X(n284) );
  SEN_AOAI211_1 U824 ( .A1(n892), .A2(n263), .B(n891), .C(n260), .X(n896) );
  SEN_AOAI211_1 U825 ( .A1(n947), .A2(n293), .B(n946), .C(n1015), .X(n957) );
  SEN_ND2_S_0P5 U826 ( .A1(n812), .A2(n814), .X(n289) );
  SEN_ND2_S_0P5 U827 ( .A1(n813), .A2(n290), .X(n815) );
  SEN_INV_S_0P5 U828 ( .A(n289), .X(n290) );
  SEN_OR2_DG_1 U829 ( .A1(n898), .A2(n403), .X(n291) );
  SEN_OR2_1 U830 ( .A1(n897), .A2(n411), .X(n292) );
  SEN_MUXI2_S_1 U831 ( .D0(n899), .D1(n902), .S(n357), .X(n900) );
  SEN_OR2_2 U832 ( .A1(n829), .A2(n828), .X(n1074) );
  SEN_INV_S_1P5 U833 ( .A(n372), .X(n598) );
  SEN_ND2_G_1 U834 ( .A1(n415), .A2(n737), .X(n738) );
  SEN_INV_S_0P5 U835 ( .A(n518), .X(n1179) );
  SEN_OAI21_S_0P5 U836 ( .A1(n994), .A2(n993), .B(n992), .X(n1027) );
  SEN_NR2_G_1 U837 ( .A1(n1055), .A2(n1054), .X(n1062) );
  SEN_AOI211_G_2 U838 ( .A1(n470), .A2(n469), .B1(n468), .B2(n535), .X(n471)
         );
  SEN_INV_S_1 U839 ( .A(n1288), .X(n315) );
  SEN_OR2_2P5 U840 ( .A1(n315), .A2(n408), .X(n314) );
  SEN_INV_1 U841 ( .A(n1175), .X(n1176) );
  SEN_OAI21_S_0P5 U842 ( .A1(n1178), .A2(n243), .B(n1177), .X(n1180) );
  SEN_INV_S_0P5 U843 ( .A(n1316), .X(n445) );
  SEN_INV_2 U844 ( .A(n867), .X(n921) );
  SEN_ND2B_V1_1 U845 ( .A(n356), .B(n384), .X(n922) );
  SEN_MUXI2_DG_1 U846 ( .D0(n1214), .D1(n1213), .S(n396), .X(n1215) );
  SEN_ND2_G_1 U847 ( .A1(n1252), .A2(n240), .X(n1253) );
  SEN_NR2_G_1 U848 ( .A1(n1025), .A2(n949), .X(n892) );
  SEN_AN2_S_4 U849 ( .A1(n826), .A2(n827), .X(n312) );
  SEN_ND2B_S_0P5 U850 ( .A(B[14]), .B(n385), .X(n919) );
  SEN_NR2_S_0P5 U851 ( .A1(n1239), .A2(n317), .X(n294) );
  SEN_NR2_T_2 U852 ( .A1(n318), .A2(n295), .X(n319) );
  SEN_INV_S_0P5 U853 ( .A(n294), .X(n295) );
  SEN_NR2_S_0P8 U854 ( .A1(n380), .A2(n353), .X(n320) );
  SEN_ND2_S_0P5 U855 ( .A1(n1379), .A2(n370), .X(n298) );
  SEN_INV_S_0P5 U856 ( .A(n370), .X(n296) );
  SEN_INV_S_0P5 U857 ( .A(n1024), .X(n993) );
  SEN_ND2_S_1 U858 ( .A1(n1076), .A2(n1075), .X(n302) );
  SEN_ND2_S_0P5 U859 ( .A1(n1077), .A2(n1078), .X(n322) );
  SEN_ND2_S_0P5 U860 ( .A1(n825), .A2(n828), .X(n718) );
  SEN_OR3B_0P5 U861 ( .B1(n382), .B2(n383), .A(n846), .X(n300) );
  SEN_OR3B_2 U862 ( .B1(n382), .B2(n383), .A(n846), .X(n856) );
  SEN_INV_2 U863 ( .A(n753), .X(n321) );
  SEN_AN3B_0P5 U864 ( .B1(n1072), .B2(n1071), .A(n1070), .X(n1075) );
  SEN_INV_S_0P5 U865 ( .A(n1093), .X(n1092) );
  SEN_OAI211_0P5 U866 ( .A1(n1224), .A2(n242), .B1(n1223), .B2(n407), .X(n1227) );
  SEN_NR2_S_0P5 U867 ( .A1(n1056), .A2(n1001), .X(n512) );
  SEN_ND2_S_0P5 U868 ( .A1(n826), .A2(n827), .X(n821) );
  SEN_ND2_S_0P5 U869 ( .A1(n1379), .A2(n367), .X(n310) );
  SEN_ND2_S_0P5 U870 ( .A1(n359), .A2(n388), .X(n1072) );
  SEN_OR3B_4 U871 ( .B1(n396), .B2(n397), .A(n1243), .X(n1244) );
  SEN_OR2_DG_1 U872 ( .A1(n1320), .A2(n410), .X(n305) );
  SEN_OR2_DG_1 U873 ( .A1(n376), .A2(n349), .X(n308) );
  SEN_INV_1 U874 ( .A(n486), .X(n638) );
  SEN_INV_2 U875 ( .A(n537), .X(n540) );
  SEN_NR2B_V1DG_1 U876 ( .A(n1109), .B(n508), .X(n509) );
  SEN_ND2_S_0P5 U877 ( .A1(n415), .A2(n1287), .X(n1265) );
  SEN_INV_S_4 U878 ( .A(n1208), .X(n1243) );
  SEN_INV_S_0P5 U879 ( .A(n1310), .X(n1279) );
  SEN_ND2_S_1P5 U880 ( .A1(n1044), .A2(n1043), .X(Z[19]) );
  SEN_INV_S_0P5 U881 ( .A(n1346), .X(n317) );
  SEN_MUXI2_DG_1 U882 ( .D0(n1037), .D1(n266), .S(n361), .X(n1039) );
  SEN_ND2_S_0P5 U883 ( .A1(n379), .A2(n352), .X(n751) );
  SEN_ND2_S_0P5 U884 ( .A1(n366), .A2(n396), .X(n1281) );
  SEN_ND2_S_0P5 U885 ( .A1(n381), .A2(B[10]), .X(n827) );
  SEN_ND2B_S_0P5 U886 ( .A(n412), .B(n1119), .X(n1117) );
  SEN_ND2_S_0P5 U887 ( .A1(n1053), .A2(n1052), .X(n1055) );
  SEN_INV_S_0P5 U888 ( .A(n1066), .X(n1069) );
  SEN_INV_S_0P5 U889 ( .A(n1188), .X(n1189) );
  SEN_INV_S_0P5 U890 ( .A(n1361), .X(n1358) );
  SEN_AOA211_DG_1 U891 ( .A1(n1110), .A2(n1109), .B(n1137), .C(n1108), .X(n326) );
  SEN_INV_S_0P5 U892 ( .A(n1319), .X(n451) );
  SEN_INV_S_0P5 U893 ( .A(n1349), .X(n1343) );
  SEN_ND2_G_1 U894 ( .A1(n1035), .A2(n1034), .X(n1041) );
  SEN_ND2B_S_0P5 U895 ( .A(n346), .B(n373), .X(n631) );
  SEN_ND2B_S_0P5 U896 ( .A(n376), .B(n349), .X(n495) );
  SEN_ND2_S_0P5 U897 ( .A1(n397), .A2(B[26]), .X(n1346) );
  SEN_OR2_DG_1 U898 ( .A1(n1291), .A2(n410), .X(n316) );
  SEN_INV_S_0P5 U899 ( .A(n419), .X(n417) );
  SEN_INV_S_0P5 U900 ( .A(n419), .X(n418) );
  SEN_ND2_S_0P5 U901 ( .A1(n415), .A2(n1222), .X(n1201) );
  SEN_AO2BB2_0P5 U902 ( .A1(n761), .A2(n411), .B1(n405), .B2(n760), .X(n764)
         );
  SEN_INV_S_0P5 U903 ( .A(n508), .X(n1082) );
  SEN_INV_S_0P5 U904 ( .A(n489), .X(n720) );
  SEN_AOAI211_1 U905 ( .A1(n459), .A2(n458), .B(n457), .C(n456), .X(n473) );
  SEN_ND2_S_0P5 U906 ( .A1(n756), .A2(n757), .X(n489) );
  SEN_ND2_S_0P5 U907 ( .A1(n421), .A2(n1202), .X(n1158) );
  SEN_OAI21_S_0P5 U908 ( .A1(n1142), .A2(n417), .B(n264), .X(n1123) );
  SEN_NR2_S_0P5 U909 ( .A1(n1171), .A2(n506), .X(n515) );
  SEN_BUF_AS_0P5 U910 ( .A(n422), .X(n421) );
  SEN_ND2B_S_0P5 U911 ( .A(n961), .B(n420), .X(n1006) );
  SEN_OAI21_S_0P5 U912 ( .A1(n1280), .A2(n1279), .B(n1306), .X(n1282) );
  SEN_NR2_G_1 U913 ( .A1(n973), .A2(n971), .X(n947) );
  SEN_INV_S_0P5 U914 ( .A(n460), .X(n1120) );
  SEN_ND2_S_0P5 U915 ( .A1(n1319), .A2(n1318), .X(n1356) );
  SEN_ND2_S_0P5 U916 ( .A1(n245), .A2(n441), .X(n443) );
  SEN_OA21_1 U917 ( .A1(n1202), .A2(n417), .B(n1294), .X(n327) );
  SEN_ND2_S_0P5 U918 ( .A1(n576), .A2(n575), .X(n577) );
  SEN_INV_S_0P5 U919 ( .A(n1367), .X(n1364) );
  SEN_MUXI2_S_0P5 U920 ( .D0(n571), .D1(n574), .S(n345), .X(n572) );
  SEN_NR2_S_0P5 U921 ( .A1(n382), .A2(n354), .X(n822) );
  SEN_ND2_S_0P5 U922 ( .A1(n260), .A2(n263), .X(n1054) );
  SEN_OAI21_G_1 U923 ( .A1(n566), .A2(n565), .B(n564), .X(Z[0]) );
  SEN_OR2_DG_1 U924 ( .A1(n356), .A2(n384), .X(n912) );
  SEN_ND2_S_0P5 U925 ( .A1(n1379), .A2(n369), .X(n332) );
  SEN_INV_S_0P5 U926 ( .A(n351), .X(n717) );
  SEN_ND2_S_0P5 U927 ( .A1(n1131), .A2(n1130), .X(n1135) );
  SEN_OA21_4 U928 ( .A1(n1222), .A2(n1221), .B(n1220), .X(n325) );
  SEN_INV_S_4 U929 ( .A(n1203), .X(n1222) );
  SEN_INV_S_0P5 U930 ( .A(n413), .X(n412) );
  SEN_INV_1 U931 ( .A(n1080), .X(n1089) );
  SEN_INV_S_0P5 U932 ( .A(n1381), .X(n1332) );
  SEN_OAI21_S_0P5 U933 ( .A1(n733), .A2(n417), .B(n1294), .X(n723) );
  SEN_OAI21_S_0P5 U934 ( .A1(n865), .A2(n887), .B(n261), .X(n870) );
  SEN_OAI21_S_0P5 U935 ( .A1(n955), .A2(n417), .B(n1294), .X(n932) );
  SEN_OAI21_S_0P5 U936 ( .A1(n923), .A2(n950), .B(n1023), .X(n926) );
  SEN_NR3_T_0P5 U937 ( .A1(n1025), .A2(n1054), .A3(n949), .X(n923) );
  SEN_AOAI211_0P5 U938 ( .A1(n868), .A2(n1053), .B(n890), .C(n263), .X(n871)
         );
  SEN_NR2B_V1DG_1 U939 ( .A(n756), .B(n474), .X(n429) );
  SEN_AN3B_0P5 U940 ( .B1(n1020), .B2(n1019), .A(n1018), .X(n1022) );
  SEN_AOI21_S_0P5 U941 ( .A1(n1308), .A2(n1307), .B(n1347), .X(n1314) );
  SEN_INV_S_0P5 U942 ( .A(n1304), .X(n1308) );
  SEN_AOI221_2 U943 ( .A1(n517), .A2(n516), .B1(n515), .B2(n514), .C(n513), 
        .X(n520) );
  SEN_OAI21_S_0P5 U944 ( .A1(n1088), .A2(n417), .B(n1294), .X(n1045) );
  SEN_OAI21_S_0P5 U945 ( .A1(n787), .A2(n786), .B(n785), .X(n793) );
  SEN_INV_S_3 U946 ( .A(n961), .X(n1013) );
  SEN_INV_S_0P5 U947 ( .A(n522), .X(n1225) );
  SEN_ND2_S_0P5 U948 ( .A1(n1120), .A2(n1191), .X(n466) );
  SEN_ND2_S_0P5 U949 ( .A1(n992), .A2(n989), .X(n507) );
  SEN_OAI21_S_0P5 U950 ( .A1(n1222), .A2(n1221), .B(n1220), .X(n1236) );
  SEN_ND2_S_0P5 U951 ( .A1(n1024), .A2(n1023), .X(n1057) );
  SEN_ND2_S_0P5 U952 ( .A1(n1109), .A2(n255), .X(n464) );
  SEN_INV_S_2 U953 ( .A(n856), .X(n894) );
  SEN_BUF_AS_0P5 U954 ( .A(n416), .X(n413) );
  SEN_INV_S_0P5 U955 ( .A(n699), .X(n485) );
  SEN_ND3_S_1 U956 ( .A1(n493), .A2(n492), .A3(n491), .X(n501) );
  SEN_AOI21B_1 U957 ( .A1(n1190), .A2(n1187), .B(n1186), .X(n1200) );
  SEN_ND3_S_0P5 U958 ( .A1(n1193), .A2(n1192), .A3(n1191), .X(n1197) );
  SEN_OR3B_0P5 U959 ( .B1(n559), .B2(n343), .A(n335), .X(n1329) );
  SEN_OAI21_S_0P5 U960 ( .A1(n1141), .A2(n1140), .B(n330), .X(n1145) );
  SEN_ND2_S_0P5 U961 ( .A1(n1319), .A2(n1318), .X(n530) );
  SEN_ND2B_V1_1 U962 ( .A(n369), .B(n400), .X(n1361) );
  SEN_AOI21B_1 U963 ( .A1(n481), .A2(n480), .B(n479), .X(n482) );
  SEN_ND2_S_0P5 U964 ( .A1(n1361), .A2(n1360), .X(n1363) );
  SEN_ND2_S_0P5 U965 ( .A1(n387), .A2(n358), .X(n1015) );
  SEN_ND2B_S_0P5 U966 ( .A(n378), .B(n351), .X(n806) );
  SEN_NR2_S_0P5 U967 ( .A1(n388), .A2(n359), .X(n977) );
  SEN_AOAI211_1 U968 ( .A1(n338), .A2(n1216), .B(n1218), .C(n1215), .X(Z[25])
         );
  SEN_ND2B_S_0P5 U969 ( .A(n382), .B(n354), .X(n809) );
  SEN_ND2B_S_0P5 U970 ( .A(n388), .B(n359), .X(n992) );
  SEN_ND2_S_0P5 U971 ( .A1(n377), .A2(n350), .X(n825) );
  SEN_ND3_S_0P5 U972 ( .A1(n807), .A2(n806), .A3(n805), .X(n811) );
  SEN_INV_S_0P5 U973 ( .A(n339), .X(n1294) );
  SEN_ND2_S_0P5 U974 ( .A1(n365), .A2(n267), .X(n1182) );
  SEN_ND2B_S_0P5 U975 ( .A(n363), .B(n392), .X(n1108) );
  SEN_ND2B_S_0P5 U976 ( .A(n359), .B(n388), .X(n995) );
  SEN_INV_S_0P5 U977 ( .A(n338), .X(n1385) );
  SEN_ND2B_S_0P5 U978 ( .A(n386), .B(n357), .X(n988) );
  SEN_ND2_S_0P5 U979 ( .A1(n349), .A2(n376), .X(n676) );
  SEN_INV_S_0P5 U980 ( .A(n386), .X(n909) );
  SEN_INV_S_0P5 U981 ( .A(n357), .X(n910) );
  SEN_AOAI211_0P5 U982 ( .A1(n392), .A2(n1105), .B(n1385), .C(n363), .X(n1106)
         );
  SEN_ND2_S_0P5 U983 ( .A1(n353), .A2(n380), .X(n781) );
  SEN_ND2B_S_0P5 U984 ( .A(n372), .B(n345), .X(n494) );
  SEN_INV_S_0P5 U985 ( .A(n345), .X(n588) );
  SEN_OA21_2 U986 ( .A1(n326), .A2(n1139), .B(n1138), .X(n330) );
  SEN_INV_S_2 U987 ( .A(n895), .X(n955) );
  SEN_INV_S_3 U988 ( .A(n1143), .X(n1202) );
  SEN_OR3B_4 U989 ( .B1(n376), .B2(n377), .A(n700), .X(n701) );
  SEN_OAI22_S_0P5 U990 ( .A1(n242), .A2(n831), .B1(n830), .B2(n409), .X(n834)
         );
  SEN_INV_S_0P5 U991 ( .A(n847), .X(n831) );
  SEN_OAI211_0P5 U992 ( .A1(n760), .A2(n403), .B1(n759), .B2(n406), .X(n765)
         );
  SEN_ND2B_S_0P5 U993 ( .A(n412), .B(n761), .X(n759) );
  SEN_OAI221_0P5 U994 ( .A1(n587), .A2(n243), .B1(n411), .B2(n570), .C(n406), 
        .X(n574) );
  SEN_INV_S_0P5 U995 ( .A(n604), .X(n605) );
  SEN_INV_S_0P5 U996 ( .A(n1060), .X(n949) );
  SEN_OAI221_0P5 U997 ( .A1(n848), .A2(n411), .B1(n847), .B2(n402), .C(n406), 
        .X(n835) );
  SEN_OAI221_0P5 U998 ( .A1(n736), .A2(n411), .B1(n734), .B2(n243), .C(n406), 
        .X(n722) );
  SEN_ND2_S_0P5 U999 ( .A1(n415), .A2(n1203), .X(n1204) );
  SEN_INV_S_0P5 U1000 ( .A(n852), .X(n849) );
  SEN_OAI22_S_0P5 U1001 ( .A1(n603), .A2(n402), .B1(n604), .B2(n409), .X(n614)
         );
  SEN_INV_S_0P5 U1002 ( .A(n606), .X(n603) );
  SEN_INV_S_0P5 U1003 ( .A(n957), .X(n954) );
  SEN_OAI211_0P5 U1004 ( .A1(n1000), .A2(n402), .B1(n999), .B2(n407), .X(n1002) );
  SEN_ND2B_S_0P5 U1005 ( .A(n412), .B(n998), .X(n999) );
  SEN_OAI211_0P5 U1006 ( .A1(n870), .A2(n242), .B1(n869), .B2(n406), .X(n875)
         );
  SEN_ND2B_S_0P5 U1007 ( .A(n411), .B(n871), .X(n869) );
  SEN_OAI211_0P5 U1008 ( .A1(n636), .A2(n402), .B1(n407), .B2(n635), .X(n640)
         );
  SEN_ND2_S_0P5 U1009 ( .A1(n415), .A2(n637), .X(n635) );
  SEN_ND3_S_0P5 U1010 ( .A1(n243), .A2(n410), .A3(n406), .X(n555) );
  SEN_OAI22_S_0P5 U1011 ( .A1(n243), .A2(n872), .B1(n871), .B2(n409), .X(n874)
         );
  SEN_INV_S_0P5 U1012 ( .A(n870), .X(n872) );
  SEN_OAI22_S_0P5 U1013 ( .A1(n600), .A2(n236), .B1(n601), .B2(n409), .X(n594)
         );
  SEN_OAI21_S_0P5 U1014 ( .A1(n1137), .A2(n1140), .B(n326), .X(n1119) );
  SEN_OAI22_S_0P5 U1015 ( .A1(n682), .A2(n242), .B1(n698), .B2(n409), .X(n685)
         );
  SEN_AO2BB2_0P5 U1016 ( .A1(n637), .A2(n411), .B1(n405), .B2(n636), .X(n639)
         );
  SEN_AO2BB2_0P5 U1017 ( .A1(n1119), .A2(n411), .B1(n405), .B2(n1118), .X(
        n1121) );
  SEN_AO2BB2_0P5 U1018 ( .A1(n1081), .A2(n411), .B1(n404), .B2(n1080), .X(
        n1083) );
  SEN_AO2BB2_0P5 U1019 ( .A1(n719), .A2(n411), .B1(n405), .B2(n734), .X(n721)
         );
  SEN_ND2_S_0P5 U1020 ( .A1(n244), .A2(n793), .X(n788) );
  SEN_ND2_S_0P5 U1021 ( .A1(n942), .A2(n1074), .X(n847) );
  SEN_ND2_S_0P5 U1022 ( .A1(n275), .A2(n1060), .X(n830) );
  SEN_INV_S_0P5 U1023 ( .A(n718), .X(n702) );
  SEN_INV_S_0P5 U1024 ( .A(n651), .X(n627) );
  SEN_ND2B_S_0P5 U1025 ( .A(n948), .B(n275), .X(n985) );
  SEN_ND3_S_0P5 U1026 ( .A1(n407), .A2(n681), .A3(n680), .X(n686) );
  SEN_ND2_S_0P5 U1027 ( .A1(n405), .A2(n682), .X(n681) );
  SEN_ND2_S_0P5 U1028 ( .A1(n415), .A2(n698), .X(n680) );
  SEN_ND2B_S_0P5 U1029 ( .A(n1118), .B(n404), .X(n1116) );
  SEN_OAI211_0P5 U1030 ( .A1(n1091), .A2(n411), .B1(n407), .B2(n1079), .X(
        n1084) );
  SEN_ND2_S_0P5 U1031 ( .A1(n405), .A2(n1089), .X(n1079) );
  SEN_INV_S_0P5 U1032 ( .A(n832), .X(n833) );
  SEN_INV_S_0P5 U1033 ( .A(n1348), .X(n1340) );
  SEN_INV_S_0P5 U1034 ( .A(n683), .X(n684) );
  SEN_INV_S_0P5 U1035 ( .A(n928), .X(n929) );
  SEN_OAI211_0P5 U1036 ( .A1(n704), .A2(n411), .B1(n407), .B2(n703), .X(n708)
         );
  SEN_INV_S_0P5 U1037 ( .A(n715), .X(n704) );
  SEN_ND2_S_0P5 U1038 ( .A1(n244), .A2(n702), .X(n703) );
  SEN_INV_S_0P5 U1039 ( .A(n1347), .X(n1353) );
  SEN_INV_S_0P5 U1040 ( .A(n581), .X(n573) );
  SEN_INV_S_0P5 U1041 ( .A(n1123), .X(n1098) );
  SEN_INV_S_0P5 U1042 ( .A(n1045), .X(n1035) );
  SEN_INV_S_0P5 U1043 ( .A(n1070), .X(n1017) );
  SEN_INV_S_0P5 U1044 ( .A(n782), .X(n754) );
  SEN_ND2_S_0P5 U1045 ( .A1(n415), .A2(n1175), .X(n1174) );
  SEN_NR2B_V1_1 U1046 ( .A(n1165), .B(n518), .X(n519) );
  SEN_INV_S_0P5 U1047 ( .A(n896), .X(n897) );
  SEN_OAI21_S_0P5 U1048 ( .A1(n1132), .A2(n322), .B(n1115), .X(n1118) );
  SEN_INV_S_0P5 U1049 ( .A(n1136), .X(n1115) );
  SEN_OAI221_0P5 U1050 ( .A1(n301), .A2(n236), .B1(n679), .B2(n410), .C(n406), 
        .X(n665) );
  SEN_AO21B_1 U1051 ( .A1(n1306), .A2(n1304), .B(n1312), .X(n1284) );
  SEN_NR3B_1 U1052 ( .A(n255), .B1(n1057), .B2(n1056), .X(n1061) );
  SEN_ND2_S_0P5 U1053 ( .A1(n414), .A2(n1264), .X(n1262) );
  SEN_AO21B_1 U1054 ( .A1(n945), .A2(n1016), .B(n975), .X(n946) );
  SEN_NR2_S_0P5 U1055 ( .A1(n866), .A2(n949), .X(n868) );
  SEN_INV_S_0P5 U1056 ( .A(n589), .X(n600) );
  SEN_ND2B_S_0P5 U1057 ( .A(n627), .B(n626), .X(n589) );
  SEN_OAI22_S_0P5 U1058 ( .A1(n662), .A2(n402), .B1(n663), .B2(n409), .X(n672)
         );
  SEN_INV_S_0P5 U1059 ( .A(n301), .X(n662) );
  SEN_ND3_S_0P5 U1060 ( .A1(n495), .A2(n324), .A3(n633), .X(n497) );
  SEN_INV_S_0P5 U1061 ( .A(n256), .X(n499) );
  SEN_AN2_S_0P5 U1062 ( .A1(n565), .A2(n559), .X(n336) );
  SEN_INV_S_0P5 U1063 ( .A(n977), .X(n978) );
  SEN_INV_S_0P5 U1064 ( .A(n1015), .X(n979) );
  SEN_AOAI211_0P5 U1065 ( .A1(n953), .A2(n952), .B(n951), .C(n1024), .X(n956)
         );
  SEN_INV_S_0P5 U1066 ( .A(n983), .X(n952) );
  SEN_AO21B_1 U1067 ( .A1(n950), .A2(n1023), .B(n989), .X(n951) );
  SEN_INV_S_0P5 U1068 ( .A(n1318), .X(n1286) );
  SEN_ND2_S_0P5 U1069 ( .A1(n1191), .A2(n1193), .X(n1137) );
  SEN_INV_S_0P5 U1070 ( .A(n757), .X(n735) );
  SEN_OR3B_0P5 U1071 ( .B1(n1056), .B2(n1057), .A(n1060), .X(n1026) );
  SEN_INV_S_0P5 U1072 ( .A(n898), .X(n893) );
  SEN_AOAI211_0P5 U1073 ( .A1(n777), .A2(n337), .B(n775), .C(n776), .X(n761)
         );
  SEN_AOAI211_0P5 U1074 ( .A1(n660), .A2(n634), .B(n657), .C(n656), .X(n637)
         );
  SEN_INV_S_0P5 U1075 ( .A(n654), .X(n634) );
  SEN_NR3_0P5 U1076 ( .A1(n985), .A2(n984), .A3(n983), .X(n996) );
  SEN_ND2_S_0P5 U1077 ( .A1(n1024), .A2(n1060), .X(n984) );
  SEN_OAI22_S_0P5 U1078 ( .A1(n569), .A2(n403), .B1(n410), .B2(n568), .X(n571)
         );
  SEN_OAI21_S_0P5 U1079 ( .A1(n498), .A2(n602), .B(n631), .X(n604) );
  SEN_INV_S_0P5 U1080 ( .A(n324), .X(n602) );
  SEN_OAI21_S_0P5 U1081 ( .A1(n916), .A2(n945), .B(n1016), .X(n925) );
  SEN_NR3_0P5 U1082 ( .A1(n1018), .A2(n1068), .A3(n238), .X(n916) );
  SEN_AOAI211_0P5 U1083 ( .A1(n432), .A2(n431), .B(n430), .C(n429), .X(n436)
         );
  SEN_AN2_S_0P5 U1084 ( .A1(n755), .A2(n812), .X(n431) );
  SEN_ND2_S_0P5 U1085 ( .A1(n720), .A2(n806), .X(n430) );
  SEN_ND2_S_0P5 U1086 ( .A1(n677), .A2(n658), .X(n426) );
  SEN_INV_S_0P5 U1087 ( .A(n948), .X(n438) );
  SEN_ND2_S_0P5 U1088 ( .A1(n873), .A2(n917), .X(n437) );
  SEN_AN2_S_0P5 U1089 ( .A1(n521), .A2(n1190), .X(n526) );
  SEN_ND2_S_0P5 U1090 ( .A1(n1225), .A2(n1220), .X(n525) );
  SEN_OAI21B_0P5 U1091 ( .A1(n778), .A2(n777), .B(n808), .X(n791) );
  SEN_ND2_S_0P5 U1092 ( .A1(n1311), .A2(n1338), .X(n1304) );
  SEN_ND2_S_0P5 U1093 ( .A1(n1024), .A2(n989), .X(n928) );
  SEN_NR3_0P5 U1094 ( .A1(n973), .A2(n972), .A3(n971), .X(n982) );
  SEN_ND2_S_0P5 U1095 ( .A1(n293), .A2(n1015), .X(n972) );
  SEN_NR2B_V1_1 U1096 ( .A(n1315), .B(n528), .X(n531) );
  SEN_INV_S_0P5 U1097 ( .A(n821), .X(n785) );
  SEN_INV_S_0P5 U1098 ( .A(n1068), .X(n1020) );
  SEN_OAI21B_0P5 U1099 ( .A1(n418), .A2(n598), .B(n581), .X(n586) );
  SEN_INV_S_0P5 U1100 ( .A(n1167), .X(n1166) );
  SEN_OAI21_S_0P5 U1101 ( .A1(n629), .A2(n648), .B(n647), .X(n636) );
  SEN_NR2_S_0P5 U1102 ( .A1(n646), .A2(n627), .X(n629) );
  SEN_OAI21_S_0P5 U1103 ( .A1(n644), .A2(n418), .B(n1294), .X(n617) );
  SEN_OAI21_S_0P5 U1104 ( .A1(n700), .A2(n418), .B(n1294), .X(n687) );
  SEN_OAI21_S_0P5 U1105 ( .A1(n789), .A2(n417), .B(n1294), .X(n766) );
  SEN_OAI21_S_0P5 U1106 ( .A1(n894), .A2(n417), .B(n1294), .X(n876) );
  SEN_ND2_S_0P5 U1107 ( .A1(n1310), .A2(n1311), .X(n1341) );
  SEN_OAI21_S_0P5 U1108 ( .A1(n274), .A2(n600), .B(n625), .X(n606) );
  SEN_ND2_S_0P5 U1109 ( .A1(n263), .A2(n1053), .X(n948) );
  SEN_INV_S_0P5 U1110 ( .A(n1111), .X(n1090) );
  SEN_ND2B_S_0P5 U1111 ( .A(n1001), .B(n992), .X(n454) );
  SEN_INV_S_0P5 U1112 ( .A(n440), .X(n455) );
  SEN_NR2_S_0P5 U1113 ( .A1(n461), .A2(n466), .X(n440) );
  SEN_OAI21_S_0P5 U1114 ( .A1(n1243), .A2(n417), .B(n1294), .X(n1228) );
  SEN_OAI21_S_0P5 U1115 ( .A1(n846), .A2(n417), .B(n1294), .X(n836) );
  SEN_OAI21_S_0P5 U1116 ( .A1(n1013), .A2(n417), .B(n1294), .X(n1004) );
  SEN_ND4B_1 U1117 ( .A(n465), .B1(n464), .B2(n463), .B3(n462), .X(n472) );
  SEN_INV_S_0P5 U1118 ( .A(n1239), .X(n1345) );
  SEN_ND2_S_0P5 U1119 ( .A1(n1280), .A2(n1281), .X(n1239) );
  SEN_NR3B_1 U1120 ( .A(n776), .B1(n762), .B2(n832), .X(n492) );
  SEN_ND2_S_0P5 U1121 ( .A1(n1192), .A2(n1028), .X(n510) );
  SEN_ND2_S_0P5 U1122 ( .A1(n415), .A2(n1176), .X(n1177) );
  SEN_INV_S_0P5 U1123 ( .A(n1317), .X(n1360) );
  SEN_ND2_S_0P5 U1124 ( .A1(n1316), .A2(n1315), .X(n1317) );
  SEN_ND2_S_0P5 U1125 ( .A1(n988), .A2(n987), .X(n950) );
  SEN_INV_S_0P5 U1126 ( .A(n697), .X(n682) );
  SEN_OAI21_S_0P5 U1127 ( .A1(n418), .A2(n582), .B(n1294), .X(n581) );
  SEN_NR2_S_0P5 U1128 ( .A1(n1358), .A2(n1324), .X(n529) );
  SEN_ND2_S_0P5 U1129 ( .A1(n976), .A2(n974), .X(n945) );
  SEN_ND2_S_0P5 U1130 ( .A1(n917), .A2(n867), .X(n890) );
  SEN_INV_S_0P5 U1131 ( .A(n1191), .X(n506) );
  SEN_ND2_S_0P5 U1132 ( .A1(n911), .A2(n912), .X(n887) );
  SEN_ND2_S_0P5 U1133 ( .A1(n1110), .A2(n1193), .X(n508) );
  SEN_ND2_S_0P5 U1134 ( .A1(n1306), .A2(n1305), .X(n1347) );
  SEN_ND2B_S_0P5 U1135 ( .A(n418), .B(n644), .X(n620) );
  SEN_OR4B_1 U1136 ( .B1(n446), .B2(n445), .B3(n1358), .A(n444), .X(n448) );
  SEN_ND2_S_0P5 U1137 ( .A1(n1220), .A2(n1186), .X(n446) );
  SEN_ND2_S_0P5 U1138 ( .A1(n995), .A2(n1024), .X(n457) );
  SEN_INV_S_0P5 U1139 ( .A(n490), .X(n873) );
  SEN_ND2_S_0P5 U1140 ( .A1(n1052), .A2(n1059), .X(n866) );
  SEN_INV_S_0P5 U1141 ( .A(n568), .X(n570) );
  SEN_ND2B_S_0P5 U1142 ( .A(n743), .B(n420), .X(n769) );
  SEN_ND2B_S_0P5 U1143 ( .A(n300), .B(n420), .X(n879) );
  SEN_ND2B_S_0P5 U1144 ( .A(n667), .B(n421), .X(n690) );
  SEN_ND2_S_0P5 U1145 ( .A1(n1082), .A2(n1192), .X(n461) );
  SEN_ND2_S_0P5 U1146 ( .A1(n1337), .A2(n1352), .X(n1348) );
  SEN_ND2_S_0P5 U1147 ( .A1(n421), .A2(n1088), .X(n1048) );
  SEN_ND2_S_0P5 U1148 ( .A1(n1186), .A2(n1190), .X(n518) );
  SEN_INV_S_0P5 U1149 ( .A(n806), .X(n484) );
  SEN_OR4B_1 U1150 ( .B1(n452), .B2(n1324), .B3(n451), .A(n450), .X(n453) );
  SEN_ND2_S_0P5 U1151 ( .A1(n1179), .A2(n1167), .X(n452) );
  SEN_ND2B_S_0P5 U1152 ( .A(n272), .B(n413), .X(n1242) );
  SEN_NR2B_V1_1 U1153 ( .A(n263), .B(n490), .X(n479) );
  SEN_ND2_S_0P5 U1154 ( .A1(n421), .A2(n955), .X(n936) );
  SEN_ND2_S_0P5 U1155 ( .A1(n421), .A2(n733), .X(n727) );
  SEN_ND2_S_0P5 U1156 ( .A1(n421), .A2(n846), .X(n840) );
  SEN_ND2_S_0P5 U1157 ( .A1(n1349), .A2(n1348), .X(n1351) );
  SEN_INV_S_0P5 U1158 ( .A(n1324), .X(n1325) );
  SEN_INV_S_0P5 U1159 ( .A(n762), .X(n763) );
  SEN_NR2_S_0P5 U1160 ( .A1(n461), .A2(n460), .X(n462) );
  SEN_ND2_S_0P5 U1161 ( .A1(n1120), .A2(n1108), .X(n513) );
  SEN_ND2_S_0P5 U1162 ( .A1(n1190), .A2(n1189), .X(n1198) );
  SEN_INV_S_0P5 U1163 ( .A(n1338), .X(n1339) );
  SEN_BUF_AS_0P5 U1164 ( .A(n416), .X(n415) );
  SEN_ND2_S_0P5 U1165 ( .A1(n591), .A2(n590), .X(n593) );
  SEN_ND2_S_0P5 U1166 ( .A1(n414), .A2(n601), .X(n590) );
  SEN_AOI21_S_0P5 U1167 ( .A1(n405), .A2(n600), .B(n408), .X(n591) );
  SEN_MUXI2_S_0P5 U1168 ( .D0(n1160), .D1(n1159), .S(n395), .X(n1184) );
  SEN_MUXI2_S_0P5 U1169 ( .D0(n1181), .D1(n1180), .S(n1179), .X(n1183) );
  SEN_ND4_S_0P5 U1170 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .X(n216)
         );
  SEN_OAI221_0P5 U1171 ( .A1(n1329), .A2(n691), .B1(n690), .B2(n376), .C(n1381), .X(n692) );
  SEN_INV_S_0P5 U1172 ( .A(n350), .X(n691) );
  SEN_OAI221_0P5 U1173 ( .A1(n1329), .A2(n780), .B1(n769), .B2(n380), .C(n1381), .X(n770) );
  SEN_OAI221_0P5 U1174 ( .A1(n1329), .A2(n886), .B1(n879), .B2(n384), .C(n1381), .X(n880) );
  SEN_OAI221_0P5 U1175 ( .A1(n1329), .A2(n1007), .B1(n1006), .B2(n388), .C(
        n1381), .X(n1008) );
  SEN_INV_S_0P5 U1176 ( .A(n360), .X(n1007) );
  SEN_OAI21_S_0P5 U1177 ( .A1(n392), .A2(n363), .B(n1111), .X(n1132) );
  SEN_AO21B_1 U1178 ( .A1(n887), .A2(n261), .B(n913), .X(n888) );
  SEN_INV_S_0P5 U1179 ( .A(n261), .X(n885) );
  SEN_ND2_S_0P5 U1180 ( .A1(n375), .A2(n348), .X(n649) );
  SEN_AO21B_1 U1181 ( .A1(n890), .A2(n263), .B(n918), .X(n891) );
  SEN_ND2B_S_0P5 U1182 ( .A(n360), .B(n389), .X(n1058) );
  SEN_ND2_S_0P5 U1183 ( .A1(n364), .A2(n394), .X(n1161) );
  SEN_INV_S_0P5 U1184 ( .A(n394), .X(n1163) );
  SEN_MUXI2_S_0P5 U1185 ( .D0(n614), .D1(n608), .S(n347), .X(n607) );
  SEN_MUXI2_S_0P5 U1186 ( .D0(n672), .D1(n665), .S(n349), .X(n664) );
  SEN_MUXI2_S_0P5 U1187 ( .D0(n861), .D1(n854), .S(n356), .X(n853) );
  SEN_OAI21_S_0P5 U1188 ( .A1(n1359), .A2(n1358), .B(n1357), .X(n1367) );
  SEN_INV_S_0P5 U1189 ( .A(n1356), .X(n1359) );
  SEN_MUXI2_S_0P5 U1190 ( .D0(n1127), .D1(n1126), .S(n393), .X(n1128) );
  SEN_OAI21_S_0P5 U1191 ( .A1(n1124), .A2(n417), .B(n1098), .X(n1127) );
  SEN_OAI221_0P5 U1192 ( .A1(n266), .A2(n1130), .B1(n1125), .B2(n392), .C(
        n1381), .X(n1126) );
  SEN_INV_S_0P5 U1193 ( .A(n392), .X(n1124) );
  SEN_ND2_S_0P5 U1194 ( .A1(n367), .A2(n398), .X(n1306) );
  SEN_ND2_S_0P5 U1195 ( .A1(n1281), .A2(n1346), .X(n1307) );
  SEN_OAI211_0P5 U1196 ( .A1(n1048), .A2(n390), .B1(n269), .B2(n1047), .X(
        n1049) );
  SEN_ND2B_S_0P5 U1197 ( .A(n1329), .B(n362), .X(n1047) );
  SEN_ND2_S_0P5 U1198 ( .A1(n368), .A2(n1379), .X(n1272) );
  SEN_OAI211_0P5 U1199 ( .A1(n936), .A2(n386), .B1(n269), .B2(n935), .X(n937)
         );
  SEN_ND2_S_0P5 U1200 ( .A1(n358), .A2(n1379), .X(n935) );
  SEN_OAI211_0P5 U1201 ( .A1(n727), .A2(n378), .B1(n269), .B2(n726), .X(n728)
         );
  SEN_ND2_S_0P5 U1202 ( .A1(n352), .A2(n1379), .X(n726) );
  SEN_OAI211_0P5 U1203 ( .A1(n840), .A2(n382), .B1(n269), .B2(n839), .X(n841)
         );
  SEN_ND2_S_0P5 U1204 ( .A1(n355), .A2(n1379), .X(n839) );
  SEN_OAI211_0P5 U1205 ( .A1(n1158), .A2(n394), .B1(n269), .B2(n1157), .X(
        n1159) );
  SEN_ND2B_S_0P5 U1206 ( .A(n1329), .B(n365), .X(n1157) );
  SEN_ND2_S_0P5 U1207 ( .A1(n1218), .A2(n1217), .X(n1310) );
  SEN_INV_S_0P5 U1208 ( .A(n396), .X(n1217) );
  SEN_INV_S_0P5 U1209 ( .A(n1099), .X(n1096) );
  SEN_INV_S_0P5 U1210 ( .A(n371), .X(n582) );
  SEN_MUXI2_S_0P5 U1211 ( .D0(n748), .D1(n741), .S(n353), .X(n740) );
  SEN_ND2_S_0P5 U1212 ( .A1(n341), .A2(n540), .X(n539) );
  SEN_ND2_S_0P5 U1213 ( .A1(n363), .A2(n392), .X(n1112) );
  SEN_ND2B_S_0P5 U1214 ( .A(n395), .B(n365), .X(n1190) );
  SEN_AO21B_1 U1215 ( .A1(n415), .A2(n1145), .B(n1144), .X(n1149) );
  SEN_MUXI2_S_0P5 U1216 ( .D0(n640), .D1(n639), .S(n638), .X(n642) );
  SEN_MUXI2_S_0P5 U1217 ( .D0(n624), .D1(n623), .S(n375), .X(n643) );
  SEN_MUXI2_S_0P5 U1218 ( .D0(n1294), .D1(n556), .S(n371), .X(n562) );
  SEN_AOI21_S_0P5 U1219 ( .A1(n560), .A2(n555), .B(n554), .X(n556) );
  SEN_ND2_S_0P5 U1220 ( .A1(n418), .A2(n1381), .X(n554) );
  SEN_ND2_S_0P5 U1221 ( .A1(n369), .A2(n400), .X(n1352) );
  SEN_AOAI211_0P5 U1222 ( .A1(n338), .A2(n1155), .B(n1164), .C(n1154), .X(
        Z[23]) );
  SEN_ND2_S_0P5 U1223 ( .A1(n394), .A2(n1146), .X(n1155) );
  SEN_AOAI211_0P5 U1224 ( .A1(n338), .A2(n804), .B(n803), .C(n802), .X(Z[11])
         );
  SEN_INV_S_0P5 U1225 ( .A(n354), .X(n803) );
  SEN_ND2_S_0P5 U1226 ( .A1(n382), .A2(n794), .X(n804) );
  SEN_MUXI2_S_0P5 U1227 ( .D0(n801), .D1(n800), .S(n382), .X(n802) );
  SEN_ND2B_S_0P5 U1228 ( .A(n394), .B(n364), .X(n1167) );
  SEN_AOAI211_0P5 U1229 ( .A1(n630), .A2(n424), .B(n256), .C(n423), .X(n428)
         );
  SEN_ND3B_0P5 U1230 ( .A(n344), .B1(n371), .B2(n494), .X(n424) );
  SEN_NR2B_V1_1 U1231 ( .A(n631), .B(n653), .X(n423) );
  SEN_INV_S_0P5 U1232 ( .A(n533), .X(n535) );
  SEN_ND2_S_0P5 U1233 ( .A1(n259), .A2(n1016), .X(n971) );
  SEN_ND2_S_0P5 U1234 ( .A1(n814), .A2(n1052), .X(n434) );
  SEN_ND2_S_0P5 U1235 ( .A1(n1023), .A2(n260), .X(n983) );
  SEN_AOI21B_0P5 U1236 ( .A1(n1364), .A2(n1363), .B(n1362), .X(n1365) );
  SEN_ND2B_S_0P5 U1237 ( .A(n367), .B(n398), .X(n1315) );
  SEN_OAI21_S_0P5 U1238 ( .A1(n400), .A2(n369), .B(n1312), .X(n1337) );
  SEN_AN2_S_0P5 U1239 ( .A1(n216), .A2(n567), .X(n338) );
  SEN_ND3_S_0P5 U1240 ( .A1(n553), .A2(n565), .A3(n341), .X(n1381) );
  SEN_EN2_0P5 U1241 ( .A1(n340), .A2(n552), .X(n553) );
  SEN_ND2B_S_0P5 U1242 ( .A(n397), .B(n1240), .X(n1311) );
  SEN_ND2B_S_0P5 U1243 ( .A(n389), .B(n360), .X(n1028) );
  SEN_AOAI211_0P5 U1244 ( .A1(n478), .A2(n477), .B(n476), .C(n475), .X(n481)
         );
  SEN_ND2_S_0P5 U1245 ( .A1(n758), .A2(n757), .X(n477) );
  SEN_ND2_S_0P5 U1246 ( .A1(n809), .A2(n805), .X(n476) );
  SEN_ND2_S_0P5 U1247 ( .A1(n395), .A2(n365), .X(n1280) );
  SEN_ND2B_S_0P5 U1248 ( .A(n366), .B(n396), .X(n1220) );
  SEN_ND2B_S_0P5 U1249 ( .A(n364), .B(n394), .X(n1165) );
  SEN_ND2B_S_0P5 U1250 ( .A(n418), .B(n401), .X(n1377) );
  SEN_INV_S_0P5 U1251 ( .A(n344), .X(n560) );
  SEN_ND2_S_0P5 U1252 ( .A1(n1138), .A2(n1168), .X(n460) );
  SEN_INV_S_0P5 U1253 ( .A(n523), .X(n1238) );
  SEN_ND3_S_0P5 U1254 ( .A1(n1138), .A2(n1165), .A3(n329), .X(n470) );
  SEN_ND3_S_0P5 U1255 ( .A1(n269), .A2(n584), .A3(n583), .X(n585) );
  SEN_ND2_S_0P5 U1256 ( .A1(n346), .A2(n1379), .X(n583) );
  SEN_ND3B_0P5 U1257 ( .A(n418), .B1(n582), .B2(n598), .X(n584) );
  SEN_ND2_S_0P5 U1258 ( .A1(n1258), .A2(n1257), .X(n1338) );
  SEN_INV_S_0P5 U1259 ( .A(n398), .X(n1257) );
  SEN_INV_S_0P5 U1260 ( .A(n364), .X(n1164) );
  SEN_ND2B_S_0P5 U1261 ( .A(n400), .B(n369), .X(n1319) );
  SEN_ND2B_S_0P5 U1262 ( .A(n365), .B(n395), .X(n1186) );
  SEN_INV_S_0P5 U1263 ( .A(n507), .X(n483) );
  SEN_AN2_S_0P5 U1264 ( .A1(n917), .A2(n867), .X(n480) );
  SEN_ND2_S_0P5 U1265 ( .A1(n391), .A2(n362), .X(n1113) );
  SEN_ND2B_S_0P5 U1266 ( .A(n401), .B(n1342), .X(n1349) );
  SEN_INV_S_0P5 U1267 ( .A(n369), .X(n1302) );
  SEN_ND2_S_0P5 U1268 ( .A1(n396), .A2(n1205), .X(n1216) );
  SEN_ND2_S_0P5 U1269 ( .A1(n398), .A2(n1247), .X(n1256) );
  SEN_AOAI211_0P5 U1270 ( .A1(n338), .A2(n714), .B(n717), .C(n713), .X(Z[7])
         );
  SEN_ND2_S_0P5 U1271 ( .A1(n378), .A2(n705), .X(n714) );
  SEN_MUXI2_S_0P5 U1272 ( .D0(n712), .D1(n711), .S(n378), .X(n713) );
  SEN_ND2_S_0P5 U1273 ( .A1(n724), .A2(n706), .X(n712) );
  SEN_AOAI211_0P5 U1274 ( .A1(n338), .A2(n580), .B(n588), .C(n579), .X(Z[1])
         );
  SEN_ND2_S_0P5 U1275 ( .A1(n372), .A2(n571), .X(n580) );
  SEN_MUXI2_S_0P5 U1276 ( .D0(n578), .D1(n577), .S(n372), .X(n579) );
  SEN_ND2_S_0P5 U1277 ( .A1(n573), .A2(n572), .X(n578) );
  SEN_INV_S_0P5 U1278 ( .A(n359), .X(n969) );
  SEN_ND2_S_0P5 U1279 ( .A1(n388), .A2(n958), .X(n970) );
  SEN_ND3B_0P5 U1280 ( .A(n622), .B1(n621), .B2(n269), .X(n623) );
  SEN_ND2B_S_0P5 U1281 ( .A(n266), .B(n348), .X(n621) );
  SEN_NR2_S_0P5 U1282 ( .A1(n620), .A2(n374), .X(n622) );
  SEN_OR3B_0P5 U1283 ( .B1(n547), .B2(n340), .A(n336), .X(n1370) );
  SEN_ND2B_S_0P5 U1284 ( .A(n1137), .B(n1168), .X(n1141) );
  SEN_ND2_S_0P5 U1285 ( .A1(n1173), .A2(n1172), .X(n1175) );
  SEN_INV_S_0P5 U1286 ( .A(n1187), .X(n1173) );
  SEN_OR4B_1 U1287 ( .B1(n1171), .B2(n1170), .B3(n1169), .A(n1195), .X(n1172)
         );
  SEN_ND3_S_0P5 U1288 ( .A1(n1168), .A2(n1191), .A3(n1167), .X(n1169) );
  SEN_OR3B_2 U1289 ( .B1(n386), .B2(n387), .A(n955), .X(n961) );
  SEN_AN2_S_0P5 U1290 ( .A1(n690), .A2(n269), .X(n668) );
  SEN_MUXI2_S_0P5 U1291 ( .D0(n666), .D1(n266), .S(n349), .X(n669) );
  SEN_INV_S_0P5 U1292 ( .A(n665), .X(n666) );
  SEN_AN2_S_0P5 U1293 ( .A1(n269), .A2(n1048), .X(n1038) );
  SEN_AN3_0P5 U1294 ( .A1(n342), .A2(n340), .A3(n336), .X(n339) );
  SEN_OR2_DG_1 U1295 ( .A1(n399), .A2(n368), .X(n1312) );
  SEN_NR2_S_0P5 U1296 ( .A1(n451), .A2(n1324), .X(n447) );
  SEN_ND2_S_0P5 U1297 ( .A1(n399), .A2(n368), .X(n1305) );
  SEN_INV_S_0P5 U1298 ( .A(n378), .X(n716) );
  SEN_OR3B_1 U1299 ( .B1(n384), .B2(n385), .A(n894), .X(n895) );
  SEN_ND2_S_0P5 U1300 ( .A1(n1191), .A2(n534), .X(n465) );
  SEN_ND2B_S_0P5 U1301 ( .A(n418), .B(n400), .X(n1328) );
  SEN_NR2_S_0P5 U1302 ( .A1(n361), .A2(n390), .X(n1064) );
  SEN_ND2B_S_0P5 U1303 ( .A(n396), .B(n366), .X(n521) );
  SEN_ND2_S_0P5 U1304 ( .A1(n361), .A2(n390), .X(n1114) );
  SEN_OR2_DG_1 U1305 ( .A1(n391), .A2(n362), .X(n1111) );
  SEN_OR2_1 U1306 ( .A1(n373), .A2(n346), .X(n628) );
  SEN_INV_S_0P5 U1307 ( .A(n342), .X(n547) );
  SEN_ND2_S_0P5 U1308 ( .A1(n368), .A2(n1385), .X(n1277) );
  SEN_ND3_S_0P5 U1309 ( .A1(n845), .A2(n844), .A3(n843), .X(Z[12]) );
  SEN_ND2_S_0P5 U1310 ( .A1(n355), .A2(n267), .X(n844) );
  SEN_MUXI2_S_0P5 U1311 ( .D0(n842), .D1(n841), .S(n383), .X(n843) );
  SEN_MUXI2_S_0P5 U1312 ( .D0(n835), .D1(n834), .S(n833), .X(n845) );
  SEN_ND3_S_0P5 U1313 ( .A1(n941), .A2(n940), .A3(n939), .X(Z[16]) );
  SEN_ND2_S_0P5 U1314 ( .A1(n358), .A2(n267), .X(n940) );
  SEN_MUXI2_S_0P5 U1315 ( .D0(n938), .D1(n937), .S(n387), .X(n939) );
  SEN_MUXI2_S_0P5 U1316 ( .D0(n931), .D1(n930), .S(n929), .X(n941) );
  SEN_ND3_S_0P5 U1317 ( .A1(n732), .A2(n731), .A3(n730), .X(Z[8]) );
  SEN_ND2_S_0P5 U1318 ( .A1(n352), .A2(n1385), .X(n731) );
  SEN_MUXI2_S_0P5 U1319 ( .D0(n729), .D1(n728), .S(n379), .X(n730) );
  SEN_MUXI2_S_0P5 U1320 ( .D0(n722), .D1(n721), .S(n720), .X(n732) );
  SEN_ND3_S_0P5 U1321 ( .A1(n696), .A2(n695), .A3(n694), .X(Z[6]) );
  SEN_ND2_S_0P5 U1322 ( .A1(n350), .A2(n1385), .X(n695) );
  SEN_MUXI2_S_0P5 U1323 ( .D0(n686), .D1(n685), .S(n684), .X(n696) );
  SEN_MUXI2_S_0P5 U1324 ( .D0(n693), .D1(n692), .S(n377), .X(n694) );
  SEN_ND3_S_0P5 U1325 ( .A1(n1012), .A2(n1011), .A3(n1010), .X(Z[18]) );
  SEN_ND2_S_0P5 U1326 ( .A1(n360), .A2(n1385), .X(n1011) );
  SEN_MUXI2_S_0P5 U1327 ( .D0(n1009), .D1(n1008), .S(n389), .X(n1010) );
  SEN_INV_S_0P5 U1328 ( .A(n366), .X(n1218) );
  SEN_INV_S_0P5 U1329 ( .A(n367), .X(n1258) );
  SEN_NR2_S_0P5 U1330 ( .A1(n1329), .A2(n1342), .X(n1331) );
  SEN_INV_0P65 U1331 ( .A(n1372), .X(n416) );
  SEN_OR3B_0P5 U1332 ( .B1(n565), .B2(n341), .A(n335), .X(n1372) );
  SEN_INV_S_0P5 U1333 ( .A(n1374), .X(n422) );
  SEN_OR3B_0P5 U1334 ( .B1(n551), .B2(n342), .A(n336), .X(n1374) );
  SEN_ND2B_S_0P5 U1335 ( .A(n340), .B(n341), .X(n544) );
  SEN_NR2_S_0P5 U1336 ( .A1(n901), .A2(n1332), .X(n904) );
  SEN_INV_0P5 U1337 ( .A(n936), .X(n901) );
  SEN_NR2_S_0P5 U1338 ( .A1(n1209), .A2(n1332), .X(n1212) );
  SEN_NR2_S_0P5 U1339 ( .A1(n1250), .A2(n1332), .X(n1252) );
  SEN_ND2_S_0P5 U1340 ( .A1(n710), .A2(n709), .X(n711) );
  SEN_NR2_S_0P5 U1341 ( .A1(n707), .A2(n1332), .X(n710) );
  SEN_MUXI2_S_0P5 U1342 ( .D0(n708), .D1(n1379), .S(n351), .X(n709) );
  SEN_INV_S_0P5 U1343 ( .A(n727), .X(n707) );
  SEN_AOI21_S_0P5 U1344 ( .A1(n582), .A2(n419), .B(n1332), .X(n576) );
  SEN_MUXI2_S_0P5 U1345 ( .D0(n574), .D1(n1379), .S(n345), .X(n575) );
  SEN_NR2_S_0P5 U1346 ( .A1(n962), .A2(n1332), .X(n965) );
  SEN_INV_0P5 U1347 ( .A(n1006), .X(n962) );
  SEN_ND2_S_0P5 U1348 ( .A1(n799), .A2(n798), .X(n800) );
  SEN_NR2_S_0P5 U1349 ( .A1(n796), .A2(n1332), .X(n799) );
  SEN_MUXI2_S_0P5 U1350 ( .D0(n797), .D1(n1379), .S(n354), .X(n798) );
  SEN_INV_0P5 U1351 ( .A(n840), .X(n796) );
  SEN_NR3_0P5 U1352 ( .A1(n563), .A2(n562), .A3(n561), .X(n564) );
  SEN_NR2_S_0P5 U1353 ( .A1(n567), .A2(n560), .X(n561) );
  SEN_INV_S_0P5 U1354 ( .A(n1004), .X(n960) );
  SEN_ND2_S_0P5 U1355 ( .A1(n837), .A2(n795), .X(n801) );
  SEN_MUXI2_S_0P5 U1356 ( .D0(n794), .D1(n797), .S(n354), .X(n795) );
  SEN_ND3_S_0P5 U1357 ( .A1(n1087), .A2(n1086), .A3(n1085), .X(Z[20]) );
  SEN_ND2_S_0P5 U1358 ( .A1(n362), .A2(n1385), .X(n1085) );
  SEN_MUXI2_S_0P5 U1359 ( .D0(n1050), .D1(n1049), .S(n391), .X(n1087) );
  SEN_MUXI2_S_0P5 U1360 ( .D0(n1084), .D1(n1083), .S(n1082), .X(n1086) );
  SEN_ND3_S_0P5 U1361 ( .A1(n597), .A2(n596), .A3(n595), .X(Z[2]) );
  SEN_ND2_S_0P5 U1362 ( .A1(n346), .A2(n1385), .X(n595) );
  SEN_MUXI2_S_0P5 U1363 ( .D0(n594), .D1(n593), .S(n256), .X(n596) );
  SEN_MUXI2_S_0P5 U1364 ( .D0(n586), .D1(n585), .S(n373), .X(n597) );
  SEN_AN2_S_0P5 U1365 ( .A1(n879), .A2(n269), .X(n857) );
  SEN_AN2_S_0P5 U1366 ( .A1(n1125), .A2(n269), .X(n1101) );
  SEN_ND2B_S_0P5 U1367 ( .A(n611), .B(n610), .X(n612) );
  SEN_AN2_S_0P5 U1368 ( .A1(n269), .A2(n620), .X(n610) );
  SEN_MUXI2_S_0P5 U1369 ( .D0(n609), .D1(n266), .S(n347), .X(n611) );
  SEN_INV_S_0P5 U1370 ( .A(n608), .X(n609) );
  SEN_AN2_S_0P5 U1371 ( .A1(n769), .A2(n1381), .X(n744) );
  SEN_ND2_S_0P5 U1372 ( .A1(n327), .A2(n1156), .X(n1160) );
  SEN_ND2B_S_0P5 U1373 ( .A(n418), .B(n394), .X(n1156) );
  SEN_ND2_S_0P5 U1374 ( .A1(n1035), .A2(n1046), .X(n1050) );
  SEN_ND2B_S_0P5 U1375 ( .A(n418), .B(n390), .X(n1046) );
  SEN_ND2_S_0P5 U1376 ( .A1(n619), .A2(n618), .X(n624) );
  SEN_ND2_S_0P5 U1377 ( .A1(n374), .A2(n420), .X(n619) );
  SEN_INV_S_0P5 U1378 ( .A(n617), .X(n618) );
  SEN_ND2_S_0P5 U1379 ( .A1(n689), .A2(n688), .X(n693) );
  SEN_ND2_S_0P5 U1380 ( .A1(n376), .A2(n420), .X(n689) );
  SEN_INV_S_0P5 U1381 ( .A(n687), .X(n688) );
  SEN_ND2_S_0P5 U1382 ( .A1(n768), .A2(n767), .X(n771) );
  SEN_ND2_S_0P5 U1383 ( .A1(n380), .A2(n420), .X(n768) );
  SEN_INV_S_0P5 U1384 ( .A(n766), .X(n767) );
  SEN_ND2_S_0P5 U1385 ( .A1(n878), .A2(n877), .X(n881) );
  SEN_ND2_S_0P5 U1386 ( .A1(n384), .A2(n420), .X(n878) );
  SEN_INV_S_0P5 U1387 ( .A(n876), .X(n877) );
  SEN_ND2_S_0P5 U1388 ( .A1(n1229), .A2(n1207), .X(n1232) );
  SEN_ND2_S_0P5 U1389 ( .A1(n396), .A2(n420), .X(n1229) );
  SEN_ND2_S_0P5 U1390 ( .A1(n398), .A2(n419), .X(n1271) );
  SEN_ND2_S_0P5 U1391 ( .A1(n725), .A2(n724), .X(n729) );
  SEN_ND2_S_0P5 U1392 ( .A1(n378), .A2(n420), .X(n725) );
  SEN_INV_S_0P5 U1393 ( .A(n723), .X(n724) );
  SEN_ND2_S_0P5 U1394 ( .A1(n838), .A2(n837), .X(n842) );
  SEN_ND2_S_0P5 U1395 ( .A1(n382), .A2(n420), .X(n838) );
  SEN_INV_S_0P5 U1396 ( .A(n836), .X(n837) );
  SEN_ND2_S_0P5 U1397 ( .A1(n934), .A2(n933), .X(n938) );
  SEN_ND2_S_0P5 U1398 ( .A1(n386), .A2(n420), .X(n934) );
  SEN_INV_S_0P5 U1399 ( .A(n932), .X(n933) );
  SEN_ND2_S_0P5 U1400 ( .A1(n1005), .A2(n960), .X(n1009) );
  SEN_ND2_S_0P5 U1401 ( .A1(n388), .A2(n420), .X(n1005) );
  SEN_AOAI211_0P5 U1402 ( .A1(n384), .A2(n861), .B(n1385), .C(n356), .X(n862)
         );
  SEN_MUXI2_S_0P5 U1403 ( .D0(n860), .D1(n859), .S(n384), .X(n863) );
  SEN_AOAI211_0P5 U1404 ( .A1(n376), .A2(n672), .B(n1385), .C(n349), .X(n673)
         );
  SEN_MUXI2_S_0P5 U1405 ( .D0(n671), .D1(n670), .S(n376), .X(n674) );
  SEN_ND2_S_0P5 U1406 ( .A1(n688), .A2(n664), .X(n671) );
  SEN_ND2_S_0P5 U1407 ( .A1(n616), .A2(n615), .X(Z[3]) );
  SEN_AOAI211_0P5 U1408 ( .A1(n374), .A2(n614), .B(n1385), .C(n347), .X(n615)
         );
  SEN_MUXI2_S_0P5 U1409 ( .D0(n613), .D1(n612), .S(n374), .X(n616) );
  SEN_ND2_S_0P5 U1410 ( .A1(n618), .A2(n607), .X(n613) );
  SEN_ND2_S_0P5 U1411 ( .A1(n750), .A2(n749), .X(Z[9]) );
  SEN_MUXI2_S_0P5 U1412 ( .D0(n747), .D1(n746), .S(n380), .X(n750) );
  SEN_ND2_S_0P5 U1413 ( .A1(n767), .A2(n740), .X(n747) );
  SEN_INV_S_0P5 U1414 ( .A(n393), .X(n1131) );
  SEN_INV_S_0P5 U1415 ( .A(B[30]), .X(n1342) );
  SEN_INV_S_0P5 U1416 ( .A(B[26]), .X(n1240) );
  SEN_INV_S_0P5 U1417 ( .A(B[22]), .X(n1130) );
  SEN_ND2B_S_0P5 U1418 ( .A(n370), .B(A[31]), .X(n534) );
  SEN_ND2B_S_0P5 U1419 ( .A(n397), .B(B[26]), .X(n523) );
  SEN_OAI211_0P5 U1420 ( .A1(n550), .A2(n216), .B1(n549), .B2(n548), .X(n563)
         );
  SEN_EN2_0P5 U1421 ( .A1(n344), .A2(SEL), .X(n550) );
  SEN_ND2B_S_0P5 U1422 ( .A(n1329), .B(n587), .X(n548) );
  SEN_ND2_S_0P5 U1423 ( .A1(n570), .A2(n555), .X(n549) );
  SEN_ND2_S_0P5 U1424 ( .A1(n401), .A2(B[30]), .X(n1350) );
  SEN_OAI211_0P5 U1425 ( .A1(n338), .A2(n1130), .B1(n1129), .B2(n1128), .X(
        Z[22]) );
  SEN_MUXI2_S_0P5 U1426 ( .D0(n1122), .D1(n1121), .S(n1120), .X(n1129) );
  SEN_OR3B_0P5 U1427 ( .B1(n559), .B2(n343), .A(n558), .X(n567) );
  SEN_EN2_0P5 U1428 ( .A1(n340), .A2(n557), .X(n558) );
  SEN_ND2_S_0P5 U1429 ( .A1(n342), .A2(SEL), .X(n557) );
  SEN_ND2B_S_0P5 U1430 ( .A(A[31]), .B(n370), .X(n533) );
  SEN_ND2B_S_0P5 U1431 ( .A(SEL), .B(n342), .X(n552) );
  SEN_ND2_S_0P5 U1432 ( .A1(B[30]), .A2(n267), .X(n1334) );
  SEN_ND3_S_0P5 U1433 ( .A1(n884), .A2(n883), .A3(n882), .X(Z[14]) );
  SEN_ND2_S_0P5 U1434 ( .A1(B[14]), .A2(n1385), .X(n883) );
  SEN_MUXI2_S_0P5 U1435 ( .D0(n881), .D1(n880), .S(n385), .X(n882) );
  SEN_MUXI2_S_0P5 U1436 ( .D0(n875), .D1(n874), .S(n873), .X(n884) );
  SEN_ND2_S_0P5 U1437 ( .A1(B[26]), .A2(n1385), .X(n1234) );
  SEN_ND3_S_0P5 U1438 ( .A1(n774), .A2(n773), .A3(n772), .X(Z[10]) );
  SEN_ND2_S_0P5 U1439 ( .A1(B[10]), .A2(n1385), .X(n773) );
  SEN_MUXI2_S_0P5 U1440 ( .D0(n771), .D1(n770), .S(n381), .X(n772) );
  SEN_MUXI2_S_0P5 U1441 ( .D0(n765), .D1(n764), .S(n763), .X(n774) );
  SEN_BUF_AS_0P5 U1442 ( .A(B[31]), .X(n370) );
  SEN_AOAI211_0P5 U1443 ( .A1(n786), .A2(n754), .B(n779), .C(n258), .X(n760)
         );
  SEN_INV_S_0P5 U1444 ( .A(n282), .X(n1178) );
  SEN_ND2_S_0P5 U1445 ( .A1(n1114), .A2(n322), .X(n1080) );
  SEN_OAI211_0P5 U1446 ( .A1(n282), .A2(n403), .B1(n407), .B2(n1174), .X(n1181) );
  SEN_OAI22_S_0P5 U1447 ( .A1(n237), .A2(n403), .B1(n1145), .B2(n409), .X(
        n1146) );
  SEN_AOI21B_0P5 U1448 ( .A1(n244), .A2(n237), .B(n407), .X(n1144) );
  SEN_AOI221_4 U1449 ( .A1(B[22]), .A2(n393), .B1(n1136), .B2(n1135), .C(n1134), .X(n1162) );
endmodule

