
module ShiftLR ( Z, X, S, LEFT, LOG, clock );
  output [31:0] Z;
  input [31:0] X;
  input [4:0] S;
  input LEFT, LOG, clock;
  wire   left_cg, log_cg, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n74, n78, n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90,
         n92, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n247, n248, n249, n250, n251,
         n252, n253, n254, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416;
  wire   [31:0] input_cg;
  wire   [4:0] shift_cg;

  SEN_FDPQ_4 \shift_cg_reg[0]  ( .D(S[0]), .CK(clock), .Q(shift_cg[0]) );
  SEN_FDPQ_4 left_cg_reg ( .D(LEFT), .CK(clock), .Q(left_cg) );
  SEN_FDPQ_D_1 log_cg_reg ( .D(LOG), .CK(clock), .Q(log_cg) );
  SEN_FDPQ_D_1 \input_cg_reg[7]  ( .D(X[7]), .CK(clock), .Q(input_cg[7]) );
  SEN_FDPQ_D_1 \input_cg_reg[6]  ( .D(X[6]), .CK(clock), .Q(input_cg[6]) );
  SEN_FDPQ_D_1 \input_cg_reg[5]  ( .D(X[5]), .CK(clock), .Q(input_cg[5]) );
  SEN_FDPQ_D_1 \input_cg_reg[4]  ( .D(X[4]), .CK(clock), .Q(input_cg[4]) );
  SEN_FDPQ_D_1 \input_cg_reg[22]  ( .D(X[22]), .CK(clock), .Q(input_cg[22]) );
  SEN_FDPQ_D_1 \input_cg_reg[21]  ( .D(X[21]), .CK(clock), .Q(input_cg[21]) );
  SEN_FDPQ_D_1 \input_cg_reg[20]  ( .D(X[20]), .CK(clock), .Q(input_cg[20]) );
  SEN_FDPQ_D_1 \input_cg_reg[15]  ( .D(X[15]), .CK(clock), .Q(input_cg[15]) );
  SEN_FDPQ_D_1 \input_cg_reg[13]  ( .D(X[13]), .CK(clock), .Q(input_cg[13]) );
  SEN_FDPQ_D_1 \input_cg_reg[29]  ( .D(X[29]), .CK(clock), .Q(input_cg[29]) );
  SEN_FDPQ_D_1 \input_cg_reg[14]  ( .D(X[14]), .CK(clock), .Q(input_cg[14]) );
  SEN_FDPQ_D_1 \input_cg_reg[12]  ( .D(X[12]), .CK(clock), .Q(input_cg[12]) );
  SEN_FDPQ_D_1 \input_cg_reg[10]  ( .D(X[10]), .CK(clock), .Q(input_cg[10]) );
  SEN_FDPQ_D_1 \input_cg_reg[9]  ( .D(X[9]), .CK(clock), .Q(input_cg[9]) );
  SEN_FDPQ_D_1 \input_cg_reg[8]  ( .D(X[8]), .CK(clock), .Q(input_cg[8]) );
  SEN_FDPQ_D_1 \input_cg_reg[23]  ( .D(X[23]), .CK(clock), .Q(input_cg[23]) );
  SEN_FDPQ_D_1 \input_cg_reg[30]  ( .D(X[30]), .CK(clock), .Q(input_cg[30]) );
  SEN_FDPQ_D_1 \input_cg_reg[28]  ( .D(X[28]), .CK(clock), .Q(input_cg[28]) );
  SEN_FDPQ_D_1 \input_cg_reg[0]  ( .D(X[0]), .CK(clock), .Q(input_cg[0]) );
  SEN_FDPQ_D_1 \input_cg_reg[17]  ( .D(X[17]), .CK(clock), .Q(input_cg[17]) );
  SEN_FDPQ_D_1 \input_cg_reg[3]  ( .D(X[3]), .CK(clock), .Q(input_cg[3]) );
  SEN_FDPQ_D_1 \input_cg_reg[2]  ( .D(X[2]), .CK(clock), .Q(input_cg[2]) );
  SEN_FDPQ_D_1 \input_cg_reg[1]  ( .D(X[1]), .CK(clock), .Q(input_cg[1]) );
  SEN_FDPQ_D_1 \input_cg_reg[11]  ( .D(X[11]), .CK(clock), .Q(input_cg[11]) );
  SEN_FDPQ_D_1 \input_cg_reg[27]  ( .D(X[27]), .CK(clock), .Q(input_cg[27]) );
  SEN_FDPQ_D_1 \input_cg_reg[18]  ( .D(X[18]), .CK(clock), .Q(input_cg[18]) );
  SEN_FDPQ_D_1 \input_cg_reg[19]  ( .D(X[19]), .CK(clock), .Q(input_cg[19]) );
  SEN_FDPQ_D_1 \input_cg_reg[26]  ( .D(X[26]), .CK(clock), .Q(input_cg[26]) );
  SEN_FDPQ_D_1 \input_cg_reg[16]  ( .D(X[16]), .CK(clock), .Q(input_cg[16]) );
  SEN_FDPQ_D_1 \input_cg_reg[24]  ( .D(X[24]), .CK(clock), .Q(input_cg[24]) );
  SEN_FDPQ_D_1 \input_cg_reg[25]  ( .D(X[25]), .CK(clock), .Q(input_cg[25]) );
  SEN_FDPQ_D_1 \input_cg_reg[31]  ( .D(X[31]), .CK(clock), .Q(input_cg[31]) );
  SEN_FDPQ_D_1 \shift_cg_reg[2]  ( .D(S[2]), .CK(clock), .Q(shift_cg[2]) );
  SEN_FDPQ_D_1 \shift_cg_reg[4]  ( .D(S[4]), .CK(clock), .Q(shift_cg[4]) );
  SEN_FDPQ_1 \shift_cg_reg[3]  ( .D(S[3]), .CK(clock), .Q(shift_cg[3]) );
  SEN_NR2_T_1P5 U290 ( .A1(log_cg), .A2(n296), .X(n152) );
  SEN_OA2BB2_1 U291 ( .A1(n80), .A2(n170), .B1(n108), .B2(n188), .X(n211) );
  SEN_INV_1 U292 ( .A(n253), .X(n332) );
  SEN_OR2_5 U293 ( .A1(n357), .A2(left_cg), .X(n294) );
  SEN_ND2_G_3 U294 ( .A1(n357), .A2(left_cg), .X(n137) );
  SEN_BUF_S_6 U295 ( .A(n212), .X(n357) );
  SEN_OAI211_3 U296 ( .A1(n66), .A2(n309), .B1(n39), .B2(n172), .X(n151) );
  SEN_AN2_S_1 U297 ( .A1(n408), .A2(n33), .X(n400) );
  SEN_EN2_S_4 U298 ( .A1(shift_cg[4]), .A2(n254), .X(n387) );
  SEN_AOI221_2 U299 ( .A1(n24), .A2(n79), .B1(n290), .B2(n272), .C(n223), .X(
        n209) );
  SEN_ND2_T_4 U300 ( .A1(n333), .A2(left_cg), .X(n254) );
  SEN_INV_2 U301 ( .A(n294), .X(n359) );
  SEN_NR2_G_0P65 U302 ( .A1(n387), .A2(left_cg), .X(n298) );
  SEN_NR2_G_1 U303 ( .A1(n387), .A2(left_cg), .X(n220) );
  SEN_INV_0P65 U304 ( .A(n32), .X(n398) );
  SEN_INV_S_0P5 U305 ( .A(n30), .X(n257) );
  SEN_AOI22_S_2 U306 ( .A1(n83), .A2(n23), .B1(n80), .B2(n290), .X(n206) );
  SEN_OAI221_2 U307 ( .A1(n188), .A2(n378), .B1(n38), .B2(n270), .C(n189), .X(
        n179) );
  SEN_AOI222_3 U308 ( .A1(n416), .A2(n287), .B1(n409), .B2(n191), .C1(n407), 
        .C2(n274), .X(n192) );
  SEN_AOI222_2 U309 ( .A1(n415), .A2(n268), .B1(n408), .B2(n117), .C1(n406), 
        .C2(n99), .X(n119) );
  SEN_AOI222_2 U310 ( .A1(n415), .A2(n99), .B1(n408), .B2(n268), .C1(n406), 
        .C2(n97), .X(n111) );
  SEN_OAI221_1 U311 ( .A1(n118), .A2(n414), .B1(n70), .B2(n410), .C(n119), .X(
        Z[4]) );
  SEN_AO221_2 U312 ( .A1(n300), .A2(input_cg[16]), .B1(n402), .B2(input_cg[0]), 
        .C(n32), .X(n115) );
  SEN_INV_S_0P5 U313 ( .A(n34), .X(n258) );
  SEN_AOI221_2 U314 ( .A1(n115), .A2(n79), .B1(n170), .B2(n272), .C(n226), .X(
        n213) );
  SEN_AOI222_1 U315 ( .A1(n416), .A2(n221), .B1(n409), .B2(n224), .C1(n407), 
        .C2(n8), .X(n225) );
  SEN_AOI222_2 U316 ( .A1(n415), .A2(n97), .B1(n408), .B2(n99), .C1(n406), 
        .C2(n95), .X(n100) );
  SEN_NR2_2 U317 ( .A1(n35), .A2(n405), .X(n376) );
  SEN_INV_S_3 U318 ( .A(n176), .X(n35) );
  SEN_AO2BB2_1 U319 ( .A1(n315), .A2(n166), .B1(n327), .B2(n290), .X(n185) );
  SEN_INV_2 U320 ( .A(n103), .X(n259) );
  SEN_INV_S_3 U321 ( .A(n259), .X(n260) );
  SEN_ND2_0P5 U322 ( .A1(left_cg), .A2(n253), .X(n252) );
  SEN_AOI222_2 U323 ( .A1(n415), .A2(n117), .B1(n408), .B2(n11), .C1(n406), 
        .C2(n268), .X(n124) );
  SEN_AO222_2 U324 ( .A1(n415), .A2(n11), .B1(n408), .B2(n146), .C1(n406), 
        .C2(n117), .X(n334) );
  SEN_INV_3 U325 ( .A(n118), .X(n11) );
  SEN_BUF_S_4 U326 ( .A(n200), .X(n305) );
  SEN_OAI22_T_0P5 U327 ( .A1(n108), .A2(n113), .B1(n314), .B2(n188), .X(n226)
         );
  SEN_AN3_S_2 U328 ( .A1(n394), .A2(n395), .A3(n302), .X(n113) );
  SEN_AOI222_2 U329 ( .A1(n416), .A2(n179), .B1(n409), .B2(n274), .C1(n407), 
        .C2(n22), .X(n184) );
  SEN_OAI222_2 U330 ( .A1(n107), .A2(n270), .B1(n101), .B2(n108), .C1(n147), 
        .C2(n405), .X(n117) );
  SEN_INV_1P25 U331 ( .A(n317), .X(n270) );
  SEN_OA222_2 U332 ( .A1(n69), .A2(n247), .B1(n53), .B2(n310), .C1(n292), .C2(
        n173), .X(n147) );
  SEN_INV_4 U333 ( .A(n136), .X(n261) );
  SEN_INV_S_3 U334 ( .A(n261), .X(n262) );
  SEN_INV_S_6 U335 ( .A(n261), .X(n263) );
  SEN_INV_S_3 U336 ( .A(n261), .X(n264) );
  SEN_BUF_3 U337 ( .A(n229), .X(n306) );
  SEN_AOI22_0P75 U338 ( .A1(n299), .A2(input_cg[15]), .B1(n359), .B2(
        input_cg[31]), .X(n229) );
  SEN_INV_1 U339 ( .A(n116), .X(n265) );
  SEN_INV_S_3 U340 ( .A(n265), .X(n266) );
  SEN_INV_3 U341 ( .A(n138), .X(n30) );
  SEN_OAI211_2 U342 ( .A1(n67), .A2(n309), .B1(n39), .B2(n177), .X(n176) );
  SEN_AOI22_T_2 U343 ( .A1(n160), .A2(input_cg[23]), .B1(n173), .B2(n178), .X(
        n177) );
  SEN_AN3_2 U344 ( .A1(n384), .A2(n385), .A3(n386), .X(n188) );
  SEN_INV_S_2 U345 ( .A(n110), .X(n267) );
  SEN_INV_2 U346 ( .A(n267), .X(n268) );
  SEN_AO221_2 U347 ( .A1(n196), .A2(n197), .B1(n198), .B2(n409), .C(n199), .X(
        Z[1]) );
  SEN_ND2_4 U348 ( .A1(n197), .A2(n85), .X(n238) );
  SEN_AN2_DG_1 U349 ( .A1(n197), .A2(n130), .X(n404) );
  SEN_NR2_G_3 U350 ( .A1(n413), .A2(n371), .X(n197) );
  SEN_INV_S_3 U351 ( .A(n291), .X(n292) );
  SEN_INV_S_0P5 U352 ( .A(n317), .X(n269) );
  SEN_INV_S_6 U353 ( .A(n81), .X(n271) );
  SEN_INV_S_0P5 U354 ( .A(n104), .X(n272) );
  SEN_INV_S_1 U355 ( .A(n269), .X(n273) );
  SEN_ND2_0P8 U356 ( .A1(n405), .A2(n82), .X(n104) );
  SEN_INV_S_2 U357 ( .A(n104), .X(n317) );
  SEN_INV_2 U358 ( .A(n318), .X(n81) );
  SEN_ND3_S_4 U359 ( .A1(n364), .A2(n365), .A3(n233), .X(n224) );
  SEN_ND3_S_4 U360 ( .A1(n335), .A2(n336), .A3(n302), .X(n178) );
  SEN_OAI221_1 U361 ( .A1(n153), .A2(n414), .B1(n45), .B2(n410), .C(n154), .X(
        Z[28]) );
  SEN_AN3_S_2 U362 ( .A1(n319), .A2(n320), .A3(n321), .X(n222) );
  SEN_ND2_0P5 U363 ( .A1(n407), .A2(n20), .X(n321) );
  SEN_BUF_S_3 U364 ( .A(n181), .X(n303) );
  SEN_AOI221_2 U365 ( .A1(input_cg[30]), .A2(n299), .B1(input_cg[14]), .B2(
        n402), .C(n32), .X(n181) );
  SEN_OAI222_2 U366 ( .A1(n70), .A2(n247), .B1(n54), .B2(n310), .C1(n266), 
        .C2(n173), .X(n200) );
  SEN_OA2BB2_4 U367 ( .A1(n140), .A2(n130), .B1(n141), .B2(n130), .X(n128) );
  SEN_AOI222_2 U368 ( .A1(n84), .A2(n142), .B1(n272), .B2(n143), .C1(n83), 
        .C2(n283), .X(n141) );
  SEN_BUF_S_3 U369 ( .A(n183), .X(n274) );
  SEN_INV_2 U370 ( .A(n238), .X(n415) );
  SEN_AOI22_S_1P5 U371 ( .A1(n300), .A2(input_cg[13]), .B1(n359), .B2(
        input_cg[29]), .X(n109) );
  SEN_INV_4 U372 ( .A(n190), .X(n37) );
  SEN_AOI221_4 U373 ( .A1(input_cg[0]), .A2(n78), .B1(n74), .B2(input_cg[16]), 
        .C(n152), .X(n190) );
  SEN_AN2_S_1 U374 ( .A1(n415), .A2(n92), .X(n324) );
  SEN_OAI221_2 U375 ( .A1(n126), .A2(n307), .B1(n288), .B2(n270), .C(n239), 
        .X(n92) );
  SEN_AOI222_3 U376 ( .A1(n415), .A2(n30), .B1(n408), .B2(n34), .C1(n406), 
        .C2(n140), .X(n154) );
  SEN_AOI222_3 U377 ( .A1(n415), .A2(n282), .B1(n408), .B2(n276), .C1(n406), 
        .C2(n285), .X(n234) );
  SEN_INV_0P8 U378 ( .A(n412), .X(n411) );
  SEN_INV_0P65 U379 ( .A(n88), .X(n412) );
  SEN_NR3_T_1 U380 ( .A1(n379), .A2(n380), .A3(n32), .X(n219) );
  SEN_OA2BB2_1 U381 ( .A1(n80), .A2(n178), .B1(n108), .B2(n175), .X(n194) );
  SEN_OA2BB2_DG_2 U382 ( .A1(n80), .A2(n115), .B1(n108), .B2(n266), .X(n114)
         );
  SEN_ND2_2 U383 ( .A1(n173), .A2(n123), .X(n108) );
  SEN_INV_S_2 U384 ( .A(n90), .X(n275) );
  SEN_INV_2 U385 ( .A(n275), .X(n276) );
  SEN_OR2_2P5 U386 ( .A1(n41), .A2(n130), .X(n353) );
  SEN_INV_S_2 U387 ( .A(n208), .X(n277) );
  SEN_INV_2 U388 ( .A(n277), .X(n278) );
  SEN_INV_1 U389 ( .A(n404), .X(n279) );
  SEN_INV_0P5 U390 ( .A(n404), .X(n280) );
  SEN_INV_1 U391 ( .A(n404), .X(n360) );
  SEN_INV_1 U392 ( .A(n404), .X(n414) );
  SEN_OAI221_2 U393 ( .A1(n240), .A2(n279), .B1(n43), .B2(n238), .C(n241), .X(
        Z[0]) );
  SEN_AOI22_T_1P5 U394 ( .A1(n371), .A2(n196), .B1(n412), .B2(input_cg[0]), 
        .X(n241) );
  SEN_AOI221_2 U395 ( .A1(n17), .A2(n79), .B1(n178), .B2(n272), .C(n215), .X(
        n201) );
  SEN_INV_S_2 U396 ( .A(n94), .X(n281) );
  SEN_INV_2 U397 ( .A(n281), .X(n282) );
  SEN_OAI221_1 U398 ( .A1(n193), .A2(n307), .B1(n155), .B2(n271), .C(n194), 
        .X(n183) );
  SEN_INV_1P5 U399 ( .A(n152), .X(n39) );
  SEN_OAI221_1 U400 ( .A1(n168), .A2(n360), .B1(n48), .B2(n410), .C(n169), .X(
        Z[25]) );
  SEN_INV_5 U401 ( .A(n137), .X(n78) );
  SEN_INV_2 U402 ( .A(n262), .X(n74) );
  SEN_OAI211_3 U403 ( .A1(n65), .A2(n309), .B1(n39), .B2(n165), .X(n142) );
  SEN_AN2_DG_2 U404 ( .A1(n415), .A2(n276), .X(n391) );
  SEN_AN2_2 U405 ( .A1(n415), .A2(n34), .X(n399) );
  SEN_AN3_S_2 U406 ( .A1(n388), .A2(n389), .A3(n390), .X(n193) );
  SEN_INV_2 U407 ( .A(n221), .X(n14) );
  SEN_ND2_S_0P5 U408 ( .A1(n409), .A2(n221), .X(n320) );
  SEN_OAI221_2 U409 ( .A1(n306), .A2(n308), .B1(n175), .B2(n271), .C(n230), 
        .X(n221) );
  SEN_AOI222_2 U410 ( .A1(n416), .A2(n274), .B1(n409), .B2(n287), .C1(n407), 
        .C2(n179), .X(n187) );
  SEN_INV_S_1P5 U411 ( .A(n238), .X(n416) );
  SEN_BUF_S_1 U412 ( .A(n144), .X(n283) );
  SEN_ND2B_2 U413 ( .A(shift_cg[2]), .B(n358), .X(n253) );
  SEN_INV_S_2 U414 ( .A(n227), .X(n284) );
  SEN_INV_2 U415 ( .A(n284), .X(n285) );
  SEN_OR2_2P5 U416 ( .A1(n361), .A2(n362), .X(n297) );
  SEN_AN2_S_1 U417 ( .A1(n409), .A2(n311), .X(n362) );
  SEN_INV_S_2 U418 ( .A(n186), .X(n286) );
  SEN_INV_2 U419 ( .A(n286), .X(n287) );
  SEN_AN2_1 U420 ( .A1(n407), .A2(n278), .X(n347) );
  SEN_INV_S_4 U421 ( .A(n312), .X(n316) );
  SEN_INV_1P5 U422 ( .A(n209), .X(n20) );
  SEN_ND2_T_2 U423 ( .A1(n353), .A2(n354), .X(n196) );
  SEN_INV_S_2 U424 ( .A(n146), .X(n41) );
  SEN_OAI222_2 U425 ( .A1(n120), .A2(n271), .B1(n121), .B2(n328), .C1(n122), 
        .C2(n405), .X(n99) );
  SEN_INV_3 U426 ( .A(n148), .X(n34) );
  SEN_OAI221_1 U427 ( .A1(n258), .A2(n414), .B1(n44), .B2(n410), .C(n149), .X(
        Z[29]) );
  SEN_AOI222_3 U428 ( .A1(n290), .A2(n79), .B1(n283), .B2(n80), .C1(n142), 
        .C2(n405), .X(n148) );
  SEN_AOI221_4 U429 ( .A1(input_cg[2]), .A2(n78), .B1(input_cg[18]), .B2(n74), 
        .C(n152), .X(n161) );
  SEN_INV_2 U430 ( .A(n168), .X(n22) );
  SEN_AOI221_2 U431 ( .A1(n23), .A2(n79), .B1(n283), .B2(n273), .C(n185), .X(
        n168) );
  SEN_NR2_S_1 U432 ( .A1(n264), .A2(n173), .X(n160) );
  SEN_INV_2 U433 ( .A(n207), .X(n23) );
  SEN_AOI221_2 U434 ( .A1(n300), .A2(input_cg[25]), .B1(n402), .B2(input_cg[9]), .C(n32), .X(n207) );
  SEN_NR3_T_2 U435 ( .A1(n368), .A2(n369), .A3(n370), .X(n210) );
  SEN_AOI22_S_1 U436 ( .A1(n83), .A2(n28), .B1(n80), .B2(n31), .X(n204) );
  SEN_INV_2 U437 ( .A(n107), .X(n24) );
  SEN_AOI221_2 U438 ( .A1(n300), .A2(input_cg[17]), .B1(n402), .B2(input_cg[1]), .C(n32), .X(n107) );
  SEN_BUF_S_2 U439 ( .A(n203), .X(n288) );
  SEN_INV_2 U440 ( .A(n120), .X(n17) );
  SEN_AOI221_2 U441 ( .A1(n299), .A2(input_cg[19]), .B1(n402), .B2(input_cg[3]), .C(n32), .X(n120) );
  SEN_EO2_2 U442 ( .A1(shift_cg[4]), .A2(n254), .X(n212) );
  SEN_INV_S_2 U443 ( .A(n164), .X(n289) );
  SEN_INV_2 U444 ( .A(n289), .X(n290) );
  SEN_OAI22_T_0P5 U445 ( .A1(n108), .A2(n193), .B1(n316), .B2(n175), .X(n215)
         );
  SEN_OA222_1 U446 ( .A1(n68), .A2(n247), .B1(n52), .B2(n310), .C1(n232), .C2(
        n173), .X(n127) );
  SEN_INV_1 U447 ( .A(n109), .X(n291) );
  SEN_AOI222_3 U448 ( .A1(n115), .A2(n273), .B1(n50), .B2(n83), .C1(n305), 
        .C2(n84), .X(n118) );
  SEN_AN2_1 U449 ( .A1(n299), .A2(input_cg[26]), .X(n379) );
  SEN_ND2_G_1 U450 ( .A1(n300), .A2(n173), .X(n247) );
  SEN_INV_2 U451 ( .A(n153), .X(n33) );
  SEN_AOI221_1 U452 ( .A1(input_cg[3]), .A2(n78), .B1(n402), .B2(input_cg[19]), 
        .C(n152), .X(n155) );
  SEN_OAI221_1 U453 ( .A1(n125), .A2(n102), .B1(n303), .B2(n271), .C(n218), 
        .X(n208) );
  SEN_AN2_1 U454 ( .A1(n408), .A2(n167), .X(n341) );
  SEN_NR2_1 U455 ( .A1(shift_cg[1]), .A2(shift_cg[0]), .X(n358) );
  SEN_INV_2 U456 ( .A(n106), .X(n312) );
  SEN_ND2_G_1 U457 ( .A1(n84), .A2(n82), .X(n106) );
  SEN_AN3_1 U458 ( .A1(n355), .A2(n356), .A3(n295), .X(n242) );
  SEN_OAI222_1 U459 ( .A1(n125), .A2(n271), .B1(n126), .B2(n328), .C1(n127), 
        .C2(n405), .X(n110) );
  SEN_OAI221_1 U460 ( .A1(n288), .A2(n102), .B1(n161), .B2(n271), .C(n204), 
        .X(n186) );
  SEN_AN2_S_1 U461 ( .A1(n407), .A2(n167), .X(n352) );
  SEN_AN2_S_1 U462 ( .A1(n406), .A2(n30), .X(n401) );
  SEN_INV_S_1 U463 ( .A(input_cg[31]), .X(n40) );
  SEN_ND2_2 U464 ( .A1(n387), .A2(left_cg), .X(n136) );
  SEN_INV_4 U465 ( .A(n405), .X(n84) );
  SEN_INV_S_1 U466 ( .A(n108), .X(n83) );
  SEN_INV_S_1 U467 ( .A(n224), .X(n3) );
  SEN_ND3_S_0P5 U468 ( .A1(n343), .A2(n344), .A3(n217), .X(Z[15]) );
  SEN_AOI222_1 U469 ( .A1(n416), .A2(n278), .B1(n409), .B2(n20), .C1(n407), 
        .C2(n15), .X(n214) );
  SEN_NR3_T_2 U470 ( .A1(n340), .A2(n341), .A3(n342), .X(n169) );
  SEN_OA2BB2_1 U471 ( .A1(n416), .A2(n131), .B1(n86), .B2(n128), .X(n139) );
  SEN_OR3_2 U472 ( .A1(n374), .A2(n375), .A3(n376), .X(n140) );
  SEN_AN2_S_1 U473 ( .A1(n416), .A2(n191), .X(n361) );
  SEN_OAI221_0P5 U474 ( .A1(n209), .A2(n414), .B1(n57), .B2(n411), .C(n210), 
        .X(Z[17]) );
  SEN_INV_S_1 U475 ( .A(n220), .X(n377) );
  SEN_BUF_3 U476 ( .A(n220), .X(n300) );
  SEN_INV_S_1 U477 ( .A(n412), .X(n410) );
  SEN_INV_S_1 U478 ( .A(n117), .X(n304) );
  SEN_OR2_1 U479 ( .A1(n86), .A2(n130), .X(n293) );
  SEN_INV_2 U480 ( .A(n301), .X(n302) );
  SEN_INV_S_1 U481 ( .A(n293), .X(n407) );
  SEN_INV_S_1 U482 ( .A(n403), .X(n408) );
  SEN_OA22_1 U483 ( .A1(n147), .A2(n84), .B1(n101), .B2(n315), .X(n295) );
  SEN_OR2_1 U484 ( .A1(n40), .A2(left_cg), .X(n296) );
  SEN_BUF_3 U485 ( .A(n298), .X(n299) );
  SEN_ND4_1 U486 ( .A1(n357), .A2(n79), .A3(n130), .A4(n86), .X(n88) );
  SEN_INV_4 U487 ( .A(n102), .X(n79) );
  SEN_ND2_S_3 U488 ( .A1(n331), .A2(n332), .X(n333) );
  SEN_AOI22_1 U489 ( .A1(n83), .A2(n170), .B1(n80), .B2(n37), .X(n189) );
  SEN_NR3_T_2 U490 ( .A1(n381), .A2(n382), .A3(n383), .X(n163) );
  SEN_AN2_S_1 U491 ( .A1(n408), .A2(n162), .X(n382) );
  SEN_OAI221_1 U492 ( .A1(n257), .A2(n360), .B1(n42), .B2(n410), .C(n139), .X(
        Z[30]) );
  SEN_OA222_3 U493 ( .A1(n67), .A2(n247), .B1(n51), .B2(n310), .C1(n306), .C2(
        n173), .X(n122) );
  SEN_INV_2 U494 ( .A(n216), .X(n301) );
  SEN_AN2_1 U495 ( .A1(n408), .A2(n278), .X(n369) );
  SEN_AOI22_S_4 U496 ( .A1(n160), .A2(input_cg[24]), .B1(n173), .B2(n37), .X(
        n172) );
  SEN_ND2_2 U497 ( .A1(n84), .A2(n173), .X(n102) );
  SEN_INV_1 U498 ( .A(n173), .X(n82) );
  SEN_ND2_T_1 U499 ( .A1(n359), .A2(n173), .X(n248) );
  SEN_EO2_G_4 U500 ( .A1(n252), .A2(shift_cg[3]), .X(n173) );
  SEN_OA2BB2_DG_1 U501 ( .A1(n83), .A2(n24), .B1(n314), .B2(n260), .X(n235) );
  SEN_OAI22_T_0P5 U502 ( .A1(n108), .A2(n260), .B1(n316), .B2(n207), .X(n223)
         );
  SEN_AOI221_2 U503 ( .A1(n299), .A2(input_cg[21]), .B1(n402), .B2(input_cg[5]), .C(n32), .X(n103) );
  SEN_AOI22_S_1 U504 ( .A1(n300), .A2(input_cg[12]), .B1(n359), .B2(
        input_cg[28]), .X(n116) );
  SEN_OA2BB2_2 U505 ( .A1(n160), .A2(input_cg[26]), .B1(n82), .B2(n161), .X(
        n159) );
  SEN_OA2BB2_2 U506 ( .A1(n160), .A2(input_cg[25]), .B1(n82), .B2(n166), .X(
        n165) );
  SEN_ND2_G_1 U507 ( .A1(n152), .A2(n387), .X(n216) );
  SEN_AOI222_2 U508 ( .A1(n415), .A2(n140), .B1(n408), .B2(n30), .C1(n406), 
        .C2(n131), .X(n149) );
  SEN_OAI221_1 U509 ( .A1(n377), .A2(n45), .B1(n264), .B2(n62), .C(n302), .X(
        n170) );
  SEN_ND2_S_0P5 U510 ( .A1(n84), .A2(n173), .X(n307) );
  SEN_ND2_S_0P5 U511 ( .A1(n84), .A2(n173), .X(n308) );
  SEN_ND2_S_0P5 U512 ( .A1(n84), .A2(n173), .X(n378) );
  SEN_NR3_T_2 U513 ( .A1(n399), .A2(n400), .A3(n401), .X(n157) );
  SEN_OAI211_3 U514 ( .A1(n64), .A2(n309), .B1(n39), .B2(n159), .X(n135) );
  SEN_OA2BB2_1 U515 ( .A1(n130), .A2(n131), .B1(n130), .B2(n132), .X(n129) );
  SEN_AOI222_1 U516 ( .A1(n133), .A2(n83), .B1(n134), .B2(n273), .C1(n135), 
        .C2(n84), .X(n132) );
  SEN_OAI221_1 U517 ( .A1(n113), .A2(n308), .B1(n190), .B2(n271), .C(n211), 
        .X(n195) );
  SEN_OAI221_1 U518 ( .A1(n377), .A2(n44), .B1(n264), .B2(n61), .C(n302), .X(
        n164) );
  SEN_BUF_3 U519 ( .A(n158), .X(n309) );
  SEN_EO2_1 U520 ( .A1(shift_cg[2]), .A2(n256), .X(n123) );
  SEN_INV_4 U521 ( .A(n302), .X(n32) );
  SEN_BUF_S_3 U522 ( .A(n248), .X(n310) );
  SEN_ND2_S_0P65 U523 ( .A1(n299), .A2(input_cg[23]), .X(n388) );
  SEN_AOI222_3 U524 ( .A1(n31), .A2(n79), .B1(n133), .B2(n80), .C1(n135), .C2(
        n405), .X(n138) );
  SEN_AN2_2 U525 ( .A1(n407), .A2(n282), .X(n393) );
  SEN_OAI221_1 U526 ( .A1(n266), .A2(n308), .B1(n188), .B2(n271), .C(n237), 
        .X(n94) );
  SEN_AOI222_3 U527 ( .A1(n170), .A2(n79), .B1(n171), .B2(n80), .C1(n151), 
        .C2(n405), .X(n153) );
  SEN_EO2_DG_2 U528 ( .A1(n251), .A2(shift_cg[1]), .X(n130) );
  SEN_BUF_S_3 U529 ( .A(n195), .X(n311) );
  SEN_INV_S_3 U530 ( .A(n312), .X(n313) );
  SEN_INV_0P8 U531 ( .A(n312), .X(n314) );
  SEN_INV_0P65 U532 ( .A(n312), .X(n315) );
  SEN_INV_4 U533 ( .A(n313), .X(n80) );
  SEN_OA2BB2_DG_1 U534 ( .A1(n83), .A2(n115), .B1(n315), .B2(n113), .X(n237)
         );
  SEN_INV_S_1 U535 ( .A(n317), .X(n318) );
  SEN_OAI221_1 U536 ( .A1(n121), .A2(n102), .B1(n193), .B2(n270), .C(n236), 
        .X(n90) );
  SEN_OAI222_2 U537 ( .A1(n38), .A2(n328), .B1(n150), .B2(n270), .C1(n36), 
        .C2(n405), .X(n131) );
  SEN_ND2_S_0P5 U538 ( .A1(n416), .A2(n8), .X(n319) );
  SEN_OR2_DG_1 U539 ( .A1(n12), .A2(n360), .X(n322) );
  SEN_OR2_DG_1 U540 ( .A1(n66), .A2(n410), .X(n323) );
  SEN_ND3_S_1 U541 ( .A1(n322), .A2(n323), .A3(n96), .X(Z[8]) );
  SEN_AN2_S_0P5 U542 ( .A1(n408), .A2(n95), .X(n325) );
  SEN_AN2_DG_1 U543 ( .A1(n406), .A2(n276), .X(n326) );
  SEN_NR3_T_2 U544 ( .A1(n324), .A2(n325), .A3(n326), .X(n96) );
  SEN_OAI221_1 U545 ( .A1(n101), .A2(n378), .B1(n260), .B2(n270), .C(n105), 
        .X(n95) );
  SEN_INV_1 U546 ( .A(n293), .X(n406) );
  SEN_INV_1 U547 ( .A(n108), .X(n327) );
  SEN_INV_0P8 U548 ( .A(n327), .X(n328) );
  SEN_OR2_DG_1 U549 ( .A1(n201), .A2(n414), .X(n329) );
  SEN_OR2_DG_1 U550 ( .A1(n55), .A2(n411), .X(n330) );
  SEN_ND3_T_0P8 U551 ( .A1(n329), .A2(n330), .A3(n202), .X(Z[19]) );
  SEN_NR2_S_3 U552 ( .A1(n363), .A2(n297), .X(n202) );
  SEN_AN2_S_0P5 U553 ( .A1(n407), .A2(n287), .X(n363) );
  SEN_INV_S_1 U554 ( .A(shift_cg[3]), .X(n331) );
  SEN_AO221_1 U555 ( .A1(n198), .A2(n404), .B1(input_cg[2]), .B2(n412), .C(
        n334), .X(Z[2]) );
  SEN_INV_S_1 U556 ( .A(n198), .X(n43) );
  SEN_OR2_DG_1 U557 ( .A1(n377), .A2(n40), .X(n335) );
  SEN_OR2_DG_1 U558 ( .A1(n263), .A2(n59), .X(n336) );
  SEN_OR2_DG_1 U559 ( .A1(n175), .A2(n102), .X(n337) );
  SEN_OR2_DG_1 U560 ( .A1(n155), .A2(n316), .X(n338) );
  SEN_OR2_2P5 U561 ( .A1(n35), .A2(n84), .X(n339) );
  SEN_ND3_T_4 U562 ( .A1(n337), .A2(n338), .A3(n339), .X(n162) );
  SEN_AN3_S_2 U563 ( .A1(n396), .A2(n397), .A3(n398), .X(n175) );
  SEN_INV_1 U564 ( .A(n162), .X(n29) );
  SEN_AN2_1 U565 ( .A1(n415), .A2(n162), .X(n340) );
  SEN_AN2_DG_1 U566 ( .A1(n406), .A2(n33), .X(n342) );
  SEN_OAI221_1 U567 ( .A1(n303), .A2(n328), .B1(n161), .B2(n315), .C(n182), 
        .X(n167) );
  SEN_OR2_DG_1 U568 ( .A1(n14), .A2(n279), .X(n343) );
  SEN_OR2_DG_1 U569 ( .A1(n59), .A2(n411), .X(n344) );
  SEN_AN2_S_0P5 U570 ( .A1(n416), .A2(n20), .X(n345) );
  SEN_AN2_DG_1 U571 ( .A1(n409), .A2(n8), .X(n346) );
  SEN_NR3_T_2 U572 ( .A1(n345), .A2(n346), .A3(n347), .X(n217) );
  SEN_OR2_DG_1 U573 ( .A1(n16), .A2(n280), .X(n348) );
  SEN_OR2_DG_1 U574 ( .A1(n51), .A2(n411), .X(n349) );
  SEN_ND3_S_1 U575 ( .A1(n348), .A2(n349), .A3(n180), .X(Z[23]) );
  SEN_AN2_S_0P5 U576 ( .A1(n416), .A2(n22), .X(n350) );
  SEN_AN2_S_0P5 U577 ( .A1(n409), .A2(n179), .X(n351) );
  SEN_NR3_T_2 U578 ( .A1(n350), .A2(n351), .A3(n352), .X(n180) );
  SEN_OA22_DG_1 U579 ( .A1(n314), .A2(n288), .B1(n108), .B2(n125), .X(n233) );
  SEN_OA22_DG_1 U580 ( .A1(n315), .A2(n107), .B1(n108), .B2(n292), .X(n105) );
  SEN_OA22_DG_1 U581 ( .A1(n314), .A2(n120), .B1(n108), .B2(n306), .X(n236) );
  SEN_OA2BB2_DG_1 U582 ( .A1(n80), .A2(n28), .B1(n108), .B2(n288), .X(n218) );
  SEN_OR2_1 U583 ( .A1(n242), .A2(n85), .X(n354) );
  SEN_ND2_S_0P5 U584 ( .A1(n243), .A2(input_cg[1]), .X(n355) );
  SEN_ND2_S_0P5 U585 ( .A1(n244), .A2(input_cg[17]), .X(n356) );
  SEN_INV_S_0P5 U586 ( .A(n130), .X(n85) );
  SEN_NR2_0P5 U587 ( .A1(n378), .A2(n377), .X(n243) );
  SEN_NR2B_V1DG_1 U588 ( .A(n359), .B(n308), .X(n244) );
  SEN_OR2_DG_1 U589 ( .A1(n232), .A2(n102), .X(n364) );
  SEN_OR2_DG_1 U590 ( .A1(n219), .A2(n270), .X(n365) );
  SEN_AOI22_S_1 U591 ( .A1(n299), .A2(input_cg[14]), .B1(n359), .B2(
        input_cg[30]), .X(n232) );
  SEN_AOI221_1 U592 ( .A1(input_cg[28]), .A2(n74), .B1(n78), .B2(input_cg[12]), 
        .C(n152), .X(n150) );
  SEN_AOI221_1 U593 ( .A1(input_cg[27]), .A2(n402), .B1(n78), .B2(input_cg[11]), .C(n152), .X(n156) );
  SEN_ND2_S_0P5 U594 ( .A1(n78), .A2(n82), .X(n158) );
  SEN_INV_2 U595 ( .A(n201), .X(n15) );
  SEN_AN3_S_1 U596 ( .A1(n372), .A2(n373), .A3(n398), .X(n125) );
  SEN_AN2_S_0P5 U597 ( .A1(n416), .A2(n15), .X(n368) );
  SEN_AN2_1 U598 ( .A1(n407), .A2(n311), .X(n370) );
  SEN_ND2_0P8 U599 ( .A1(input_cg[1]), .A2(n78), .X(n366) );
  SEN_ND2_T_0P5 U600 ( .A1(n402), .A2(input_cg[17]), .X(n367) );
  SEN_AN3_S_2 U601 ( .A1(n366), .A2(n367), .A3(n39), .X(n166) );
  SEN_INV_3 U602 ( .A(n263), .X(n402) );
  SEN_BUF_1 U603 ( .A(shift_cg[0]), .X(n371) );
  SEN_ND2_S_0P5 U604 ( .A1(n299), .A2(input_cg[18]), .X(n372) );
  SEN_ND2_S_0P5 U605 ( .A1(n402), .A2(input_cg[2]), .X(n373) );
  SEN_NR2_S_0P5 U606 ( .A1(n155), .A2(n328), .X(n374) );
  SEN_NR2_S_0P5 U607 ( .A1(n156), .A2(n270), .X(n375) );
  SEN_BUF_6 U608 ( .A(n123), .X(n405) );
  SEN_INV_1 U609 ( .A(n219), .X(n28) );
  SEN_ND2_S_0P5 U610 ( .A1(n402), .A2(input_cg[7]), .X(n389) );
  SEN_AN2_1 U611 ( .A1(n406), .A2(n34), .X(n383) );
  SEN_OAI221_1 U612 ( .A1(n27), .A2(n279), .B1(n47), .B2(n410), .C(n163), .X(
        Z[26]) );
  SEN_AN2_S_0P5 U613 ( .A1(n74), .A2(input_cg[10]), .X(n380) );
  SEN_OAI221_1 U614 ( .A1(n26), .A2(n414), .B1(n65), .B2(n411), .C(n89), .X(
        Z[9]) );
  SEN_AN2_S_0P5 U615 ( .A1(n409), .A2(n92), .X(n392) );
  SEN_AN2_S_0P5 U616 ( .A1(n415), .A2(n33), .X(n381) );
  SEN_ND2_S_0P5 U617 ( .A1(n299), .A2(input_cg[24]), .X(n384) );
  SEN_ND2_G_0P65 U618 ( .A1(n402), .A2(input_cg[8]), .X(n385) );
  SEN_INV_0P5 U619 ( .A(n32), .X(n386) );
  SEN_INV_S_0P5 U620 ( .A(n32), .X(n390) );
  SEN_OA22_DG_1 U621 ( .A1(n108), .A2(n120), .B1(n314), .B2(n193), .X(n230) );
  SEN_OA22_DG_1 U622 ( .A1(n316), .A2(n125), .B1(n108), .B2(n232), .X(n239) );
  SEN_AOI221_1 U623 ( .A1(n300), .A2(input_cg[22]), .B1(n402), .B2(input_cg[6]), .C(n32), .X(n203) );
  SEN_AOI222_1 U624 ( .A1(n416), .A2(n167), .B1(n409), .B2(n22), .C1(n407), 
        .C2(n162), .X(n174) );
  SEN_NR3_T_2 U625 ( .A1(n391), .A2(n392), .A3(n393), .X(n89) );
  SEN_ND2_S_0P5 U626 ( .A1(n300), .A2(input_cg[20]), .X(n394) );
  SEN_ND2_S_0P5 U627 ( .A1(n74), .A2(input_cg[4]), .X(n395) );
  SEN_ND2_S_0P5 U628 ( .A1(n300), .A2(input_cg[27]), .X(n396) );
  SEN_ND2_S_0P5 U629 ( .A1(n402), .A2(input_cg[11]), .X(n397) );
  SEN_INV_1 U630 ( .A(n112), .X(n50) );
  SEN_INV_1 U631 ( .A(n303), .X(n31) );
  SEN_AOI22_0P5 U632 ( .A1(n300), .A2(input_cg[9]), .B1(n359), .B2(
        input_cg[25]), .X(n101) );
  SEN_AOI22_0P5 U633 ( .A1(n299), .A2(input_cg[11]), .B1(n359), .B2(
        input_cg[27]), .X(n121) );
  SEN_OAI221_1 U634 ( .A1(n121), .A2(n316), .B1(n122), .B2(n84), .C(n249), .X(
        n146) );
  SEN_AOI22_0P5 U635 ( .A1(n300), .A2(input_cg[10]), .B1(n359), .B2(
        input_cg[26]), .X(n126) );
  SEN_INV_S_0P5 U636 ( .A(n167), .X(n27) );
  SEN_OAI221_0P5 U637 ( .A1(n263), .A2(n42), .B1(n137), .B2(n60), .C(n39), .X(
        n134) );
  SEN_OAI221_0P5 U638 ( .A1(n69), .A2(n137), .B1(n263), .B2(n53), .C(n39), .X(
        n144) );
  SEN_OAI221_0P5 U639 ( .A1(n68), .A2(n137), .B1(n264), .B2(n52), .C(n39), .X(
        n133) );
  SEN_INV_2 U640 ( .A(n213), .X(n8) );
  SEN_OAI221_0P5 U641 ( .A1(n70), .A2(n137), .B1(n263), .B2(n54), .C(n39), .X(
        n171) );
  SEN_INV_S_0P5 U642 ( .A(n99), .X(n18) );
  SEN_OAI221_1 U643 ( .A1(n112), .A2(n378), .B1(n113), .B2(n271), .C(n114), 
        .X(n97) );
  SEN_OAI221_0P5 U644 ( .A1(n61), .A2(n137), .B1(n264), .B2(n44), .C(n39), .X(
        n143) );
  SEN_INV_S_0P5 U645 ( .A(n268), .X(n6) );
  SEN_INV_S_0P5 U646 ( .A(n191), .X(n21) );
  SEN_INV_S_0P5 U647 ( .A(n274), .X(n16) );
  SEN_INV_S_0P5 U648 ( .A(n287), .X(n5) );
  SEN_INV_S_0P5 U649 ( .A(n285), .X(n19) );
  SEN_INV_S_0P5 U650 ( .A(n92), .X(n2) );
  SEN_INV_S_0P5 U651 ( .A(n282), .X(n7) );
  SEN_INV_S_0P5 U652 ( .A(n95), .X(n26) );
  SEN_INV_S_0P5 U653 ( .A(n97), .X(n12) );
  SEN_OR2_1 U654 ( .A1(n85), .A2(n86), .X(n403) );
  SEN_INV_S_0P5 U655 ( .A(n151), .X(n36) );
  SEN_OAI221_0P5 U656 ( .A1(n126), .A2(n314), .B1(n127), .B2(n84), .C(n250), 
        .X(n198) );
  SEN_AOI22_0P5 U657 ( .A1(n300), .A2(input_cg[8]), .B1(n359), .B2(
        input_cg[24]), .X(n112) );
  SEN_AOI222_0P5 U658 ( .A1(n405), .A2(n305), .B1(n244), .B2(input_cg[16]), 
        .C1(n80), .C2(n50), .X(n240) );
  SEN_INV_S_0P5 U659 ( .A(n179), .X(n10) );
  SEN_INV_S_0P5 U660 ( .A(n276), .X(n13) );
  SEN_INV_S_0P5 U661 ( .A(n278), .X(n4) );
  SEN_NR2B_V1_1 U662 ( .A(left_cg), .B(n358), .X(n256) );
  SEN_INV_S_1 U663 ( .A(n171), .X(n38) );
  SEN_INV_S_1 U664 ( .A(n403), .X(n409) );
  SEN_INV_S_1 U665 ( .A(n88), .X(n413) );
  SEN_OAI221_1 U666 ( .A1(n292), .A2(n307), .B1(n207), .B2(n270), .C(n235), 
        .X(n227) );
  SEN_OAI221_1 U667 ( .A1(n260), .A2(n307), .B1(n166), .B2(n270), .C(n206), 
        .X(n191) );
  SEN_OAI221_1 U668 ( .A1(n304), .A2(n360), .B1(n69), .B2(n410), .C(n111), .X(
        Z[5]) );
  SEN_OAI221_1 U669 ( .A1(n2), .A2(n360), .B1(n64), .B2(n410), .C(n234), .X(
        Z[10]) );
  SEN_OAI221_1 U670 ( .A1(n19), .A2(n280), .B1(n61), .B2(n411), .C(n225), .X(
        Z[13]) );
  SEN_OAI221_1 U671 ( .A1(n18), .A2(n280), .B1(n67), .B2(n410), .C(n98), .X(
        Z[7]) );
  SEN_AOI222_1 U672 ( .A1(n415), .A2(n95), .B1(n408), .B2(n97), .C1(n406), 
        .C2(n92), .X(n98) );
  SEN_OAI221_1 U673 ( .A1(n5), .A2(n280), .B1(n52), .B2(n411), .C(n184), .X(
        Z[22]) );
  SEN_OAI221_1 U674 ( .A1(n3), .A2(n414), .B1(n60), .B2(n411), .C(n222), .X(
        Z[14]) );
  SEN_OAI221_1 U675 ( .A1(n9), .A2(n360), .B1(n54), .B2(n411), .C(n192), .X(
        Z[20]) );
  SEN_OAI221_1 U676 ( .A1(n6), .A2(n279), .B1(n68), .B2(n410), .C(n100), .X(
        Z[6]) );
  SEN_OAI221_1 U677 ( .A1(n7), .A2(n279), .B1(n62), .B2(n411), .C(n228), .X(
        Z[12]) );
  SEN_AOI222_1 U678 ( .A1(n416), .A2(n224), .B1(n409), .B2(n285), .C1(n407), 
        .C2(n221), .X(n228) );
  SEN_OAI221_1 U679 ( .A1(n21), .A2(n280), .B1(n53), .B2(n411), .C(n187), .X(
        Z[21]) );
  SEN_AOI22_S_1 U680 ( .A1(n79), .A2(n28), .B1(n273), .B2(n133), .X(n182) );
  SEN_AOI22_1 U681 ( .A1(n243), .A2(input_cg[3]), .B1(n244), .B2(input_cg[19]), 
        .X(n249) );
  SEN_AOI22_1 U682 ( .A1(n243), .A2(input_cg[2]), .B1(n244), .B2(input_cg[18]), 
        .X(n250) );
  SEN_INV_S_1 U683 ( .A(input_cg[25]), .X(n48) );
  SEN_OAI221_1 U684 ( .A1(n41), .A2(n414), .B1(n71), .B2(n410), .C(n124), .X(
        Z[3]) );
  SEN_INV_S_1 U685 ( .A(input_cg[3]), .X(n71) );
  SEN_OAI221_1 U686 ( .A1(n10), .A2(n360), .B1(n49), .B2(n411), .C(n174), .X(
        Z[24]) );
  SEN_INV_S_1 U687 ( .A(input_cg[24]), .X(n49) );
  SEN_OAI221_1 U688 ( .A1(n13), .A2(n414), .B1(n63), .B2(n410), .C(n231), .X(
        Z[11]) );
  SEN_INV_S_1 U689 ( .A(input_cg[11]), .X(n63) );
  SEN_AOI222_1 U690 ( .A1(n415), .A2(n285), .B1(n409), .B2(n282), .C1(n407), 
        .C2(n224), .X(n231) );
  SEN_INV_S_1 U691 ( .A(input_cg[26]), .X(n47) );
  SEN_OAI221_1 U692 ( .A1(n213), .A2(n360), .B1(n58), .B2(n411), .C(n214), .X(
        Z[16]) );
  SEN_INV_S_1 U693 ( .A(input_cg[16]), .X(n58) );
  SEN_INV_S_1 U694 ( .A(input_cg[17]), .X(n57) );
  SEN_INV_S_1 U695 ( .A(input_cg[19]), .X(n55) );
  SEN_OAI221_1 U696 ( .A1(n29), .A2(n280), .B1(n46), .B2(n410), .C(n157), .X(
        Z[27]) );
  SEN_INV_S_1 U697 ( .A(input_cg[27]), .X(n46) );
  SEN_OAI221_1 U698 ( .A1(n4), .A2(n279), .B1(n56), .B2(n411), .C(n205), .X(
        Z[18]) );
  SEN_INV_S_1 U699 ( .A(input_cg[18]), .X(n56) );
  SEN_AOI222_1 U700 ( .A1(n416), .A2(n311), .B1(n408), .B2(n15), .C1(n407), 
        .C2(n191), .X(n205) );
  SEN_INV_S_1 U701 ( .A(input_cg[29]), .X(n44) );
  SEN_INV_S_1 U702 ( .A(input_cg[13]), .X(n61) );
  SEN_INV_S_1 U703 ( .A(input_cg[9]), .X(n65) );
  SEN_INV_S_1 U704 ( .A(input_cg[10]), .X(n64) );
  SEN_INV_S_1 U705 ( .A(input_cg[20]), .X(n54) );
  SEN_INV_S_1 U706 ( .A(input_cg[4]), .X(n70) );
  SEN_INV_S_1 U707 ( .A(input_cg[21]), .X(n53) );
  SEN_INV_S_1 U708 ( .A(input_cg[22]), .X(n52) );
  SEN_INV_S_1 U709 ( .A(input_cg[7]), .X(n67) );
  SEN_INV_S_1 U710 ( .A(input_cg[5]), .X(n69) );
  SEN_INV_S_1 U711 ( .A(input_cg[6]), .X(n68) );
  SEN_INV_S_1 U712 ( .A(input_cg[12]), .X(n62) );
  SEN_INV_S_1 U713 ( .A(input_cg[14]), .X(n60) );
  SEN_INV_S_1 U714 ( .A(input_cg[8]), .X(n66) );
  SEN_INV_S_1 U715 ( .A(input_cg[15]), .X(n59) );
  SEN_INV_S_1 U716 ( .A(input_cg[23]), .X(n51) );
  SEN_AO22_1 U717 ( .A1(n406), .A2(n11), .B1(n413), .B2(input_cg[1]), .X(n199)
         );
  SEN_INV_S_1 U718 ( .A(input_cg[28]), .X(n45) );
  SEN_INV_S_1 U719 ( .A(input_cg[30]), .X(n42) );
  SEN_ND2_S_0P5 U720 ( .A1(n371), .A2(left_cg), .X(n251) );
  SEN_INV_S_1 U721 ( .A(n371), .X(n86) );
  SEN_INV_S_1 U722 ( .A(n311), .X(n9) );
  SEN_OAI222_1 U723 ( .A1(n371), .A2(n128), .B1(n129), .B2(n86), .C1(n40), 
        .C2(n411), .X(Z[31]) );
  SEN_FDPQ_2 \shift_cg_reg[1]  ( .D(S[1]), .CK(clock), .Q(shift_cg[1]) );
endmodule

