
module ShiftLR ( Z, X, S, LEFT, LOG, clock );
  output [31:0] Z;
  input [31:0] X;
  input [4:0] S;
  input LEFT, LOG, clock;
  wire   left_cg, log_cg, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n89, n90, n92, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294;
  wire   [31:0] input_cg;
  wire   [4:0] shift_cg;

  SEN_FDPQ_D_1 log_cg_reg ( .D(LOG), .CK(clock), .Q(log_cg) );
  SEN_FDPQ_D_1 \input_cg_reg[7]  ( .D(X[7]), .CK(clock), .Q(input_cg[7]) );
  SEN_FDPQ_D_1 \input_cg_reg[6]  ( .D(X[6]), .CK(clock), .Q(input_cg[6]) );
  SEN_FDPQ_D_1 \input_cg_reg[5]  ( .D(X[5]), .CK(clock), .Q(input_cg[5]) );
  SEN_FDPQ_D_1 \input_cg_reg[4]  ( .D(X[4]), .CK(clock), .Q(input_cg[4]) );
  SEN_FDPQ_D_1 \input_cg_reg[22]  ( .D(X[22]), .CK(clock), .Q(input_cg[22]) );
  SEN_FDPQ_D_1 \input_cg_reg[21]  ( .D(X[21]), .CK(clock), .Q(input_cg[21]) );
  SEN_FDPQ_D_1 \input_cg_reg[20]  ( .D(X[20]), .CK(clock), .Q(input_cg[20]) );
  SEN_FDPQ_D_1 \input_cg_reg[15]  ( .D(X[15]), .CK(clock), .Q(input_cg[15]) );
  SEN_FDPQ_D_1 \input_cg_reg[13]  ( .D(X[13]), .CK(clock), .Q(input_cg[13]) );
  SEN_FDPQ_D_1 \input_cg_reg[31]  ( .D(X[31]), .CK(clock), .Q(input_cg[31]) );
  SEN_FDPQ_D_1 \input_cg_reg[29]  ( .D(X[29]), .CK(clock), .Q(input_cg[29]) );
  SEN_FDPQ_D_1 \input_cg_reg[14]  ( .D(X[14]), .CK(clock), .Q(input_cg[14]) );
  SEN_FDPQ_D_1 \input_cg_reg[12]  ( .D(X[12]), .CK(clock), .Q(input_cg[12]) );
  SEN_FDPQ_D_1 \input_cg_reg[10]  ( .D(X[10]), .CK(clock), .Q(input_cg[10]) );
  SEN_FDPQ_D_1 \input_cg_reg[9]  ( .D(X[9]), .CK(clock), .Q(input_cg[9]) );
  SEN_FDPQ_D_1 \input_cg_reg[8]  ( .D(X[8]), .CK(clock), .Q(input_cg[8]) );
  SEN_FDPQ_D_1 \input_cg_reg[23]  ( .D(X[23]), .CK(clock), .Q(input_cg[23]) );
  SEN_FDPQ_D_1 \input_cg_reg[30]  ( .D(X[30]), .CK(clock), .Q(input_cg[30]) );
  SEN_FDPQ_D_1 \input_cg_reg[28]  ( .D(X[28]), .CK(clock), .Q(input_cg[28]) );
  SEN_FDPQ_D_1 \input_cg_reg[0]  ( .D(X[0]), .CK(clock), .Q(input_cg[0]) );
  SEN_FDPQ_D_1 \input_cg_reg[17]  ( .D(X[17]), .CK(clock), .Q(input_cg[17]) );
  SEN_FDPQ_D_1 \input_cg_reg[3]  ( .D(X[3]), .CK(clock), .Q(input_cg[3]) );
  SEN_FDPQ_D_1 \input_cg_reg[2]  ( .D(X[2]), .CK(clock), .Q(input_cg[2]) );
  SEN_FDPQ_D_1 \input_cg_reg[1]  ( .D(X[1]), .CK(clock), .Q(input_cg[1]) );
  SEN_FDPQ_D_1 \input_cg_reg[11]  ( .D(X[11]), .CK(clock), .Q(input_cg[11]) );
  SEN_FDPQ_D_1 \input_cg_reg[27]  ( .D(X[27]), .CK(clock), .Q(input_cg[27]) );
  SEN_FDPQ_D_1 \input_cg_reg[18]  ( .D(X[18]), .CK(clock), .Q(input_cg[18]) );
  SEN_FDPQ_D_1 \input_cg_reg[19]  ( .D(X[19]), .CK(clock), .Q(input_cg[19]) );
  SEN_FDPQ_D_1 \input_cg_reg[26]  ( .D(X[26]), .CK(clock), .Q(input_cg[26]) );
  SEN_FDPQ_D_1 \input_cg_reg[25]  ( .D(X[25]), .CK(clock), .Q(input_cg[25]) );
  SEN_FDPQ_D_1 \input_cg_reg[16]  ( .D(X[16]), .CK(clock), .Q(input_cg[16]) );
  SEN_FDPQ_D_1 \input_cg_reg[24]  ( .D(X[24]), .CK(clock), .Q(input_cg[24]) );
  SEN_FDPQ_D_1 \shift_cg_reg[4]  ( .D(S[4]), .CK(clock), .Q(shift_cg[4]) );
  SEN_FDPQ_D_1 \shift_cg_reg[2]  ( .D(S[2]), .CK(clock), .Q(shift_cg[2]) );
  SEN_FDPQ_D_1 \shift_cg_reg[3]  ( .D(S[3]), .CK(clock), .Q(shift_cg[3]) );
  SEN_FDPQ_1 \shift_cg_reg[0]  ( .D(S[0]), .CK(clock), .Q(shift_cg[0]) );
  SEN_FDPQ_1 left_cg_reg ( .D(LEFT), .CK(clock), .Q(left_cg) );
  SEN_INV_S_1 U290 ( .A(n281), .X(n291) );
  SEN_OAI221_0P5 U291 ( .A1(n16), .A2(n292), .B1(n51), .B2(n289), .C(n180), 
        .X(Z[23]) );
  SEN_NR2_S_0P5 U292 ( .A1(n75), .A2(left_cg), .X(n269) );
  SEN_INV_2 U293 ( .A(n212), .X(n75) );
  SEN_ND2_G_0P65 U294 ( .A1(n269), .A2(n173), .X(n247) );
  SEN_AN2_2 U295 ( .A1(n197), .A2(n130), .X(n281) );
  SEN_OAI211_2 U296 ( .A1(n66), .A2(n158), .B1(n39), .B2(n172), .X(n151) );
  SEN_INV_1P5 U297 ( .A(n153), .X(n33) );
  SEN_ND2B_V1_2 U298 ( .A(shift_cg[2]), .B(n255), .X(n253) );
  SEN_AOI221_1 U299 ( .A1(n220), .A2(input_cg[24]), .B1(n74), .B2(input_cg[8]), 
        .C(n32), .X(n188) );
  SEN_OAI222_0P5 U300 ( .A1(n175), .A2(n102), .B1(n155), .B2(n258), .C1(n35), 
        .C2(n84), .X(n162) );
  SEN_AN4_0P5 U301 ( .A1(n212), .A2(n79), .A3(n130), .A4(n86), .X(n257) );
  SEN_ND2_G_1 U302 ( .A1(n212), .A2(left_cg), .X(n137) );
  SEN_NR2_1 U303 ( .A1(n75), .A2(left_cg), .X(n220) );
  SEN_ND2_S_0P5 U304 ( .A1(n84), .A2(n82), .X(n258) );
  SEN_OAI221_0P5 U305 ( .A1(n121), .A2(n258), .B1(n122), .B2(n84), .C(n249), 
        .X(n146) );
  SEN_OAI22_S_0P5 U306 ( .A1(n147), .A2(n84), .B1(n101), .B2(n258), .X(n245)
         );
  SEN_INV_2 U307 ( .A(n282), .X(n84) );
  SEN_ND2_S_0P5 U308 ( .A1(n84), .A2(n82), .X(n106) );
  SEN_INV_S_1 U309 ( .A(n79), .X(n259) );
  SEN_INV_S_1 U310 ( .A(n102), .X(n79) );
  SEN_INV_S_1 U311 ( .A(n136), .X(n260) );
  SEN_INV_S_1 U312 ( .A(n136), .X(n74) );
  SEN_INV_S_1 U313 ( .A(n81), .X(n261) );
  SEN_ND2_G_1 U314 ( .A1(n275), .A2(shift_cg[4]), .X(n278) );
  SEN_ND2_G_1 U315 ( .A1(n254), .A2(n276), .X(n277) );
  SEN_ND2_0P5 U316 ( .A1(n152), .A2(n75), .X(n216) );
  SEN_OAI222_0P75 U317 ( .A1(n107), .A2(n104), .B1(n101), .B2(n108), .C1(n147), 
        .C2(n282), .X(n117) );
  SEN_BUF_S_1 U318 ( .A(n123), .X(n282) );
  SEN_ND2_G_1 U319 ( .A1(n273), .A2(n274), .X(n173) );
  SEN_ND2_G_1 U320 ( .A1(n271), .A2(shift_cg[3]), .X(n274) );
  SEN_INV_S_1 U321 ( .A(n254), .X(n275) );
  SEN_AN2_S_1 U322 ( .A1(n293), .A2(n11), .X(n262) );
  SEN_AN2_S_0P5 U323 ( .A1(n285), .A2(n146), .X(n263) );
  SEN_AN2_S_1 U324 ( .A1(n283), .A2(n117), .X(n264) );
  SEN_NR3_G_1 U325 ( .A1(n262), .A2(n263), .A3(n264), .X(n145) );
  SEN_INV_S_1 U326 ( .A(n216), .X(n32) );
  SEN_INV_S_0P5 U327 ( .A(n120), .X(n17) );
  SEN_INV_1 U328 ( .A(n137), .X(n78) );
  SEN_AOI22_S_1 U329 ( .A1(n160), .A2(input_cg[24]), .B1(n173), .B2(n37), .X(
        n172) );
  SEN_INV_S_1 U330 ( .A(shift_cg[4]), .X(n276) );
  SEN_ND2_S_0P5 U331 ( .A1(n173), .A2(n282), .X(n265) );
  SEN_OAI221_0P5 U332 ( .A1(n113), .A2(n102), .B1(n190), .B2(n104), .C(n211), 
        .X(n195) );
  SEN_INV_S_0P5 U333 ( .A(n287), .X(n290) );
  SEN_AOI222_0P5 U334 ( .A1(n170), .A2(n79), .B1(n171), .B2(n80), .C1(n151), 
        .C2(n282), .X(n153) );
  SEN_NR2B_V1_1 U335 ( .A(n246), .B(n102), .X(n244) );
  SEN_AOI22_0P5 U336 ( .A1(n79), .A2(n28), .B1(n81), .B2(n133), .X(n182) );
  SEN_AN3_S_1 U337 ( .A1(n266), .A2(n267), .A3(n268), .X(n214) );
  SEN_ND2_G_1 U338 ( .A1(n294), .A2(n208), .X(n266) );
  SEN_ND2_S_0P5 U339 ( .A1(n284), .A2(n15), .X(n268) );
  SEN_AOI22_0P5 U340 ( .A1(n160), .A2(input_cg[23]), .B1(n173), .B2(n178), .X(
        n177) );
  SEN_INV_S_1 U341 ( .A(n106), .X(n80) );
  SEN_INV_1 U342 ( .A(n108), .X(n83) );
  SEN_INV_S_1 U343 ( .A(n104), .X(n81) );
  SEN_INV_1 U344 ( .A(n201), .X(n15) );
  SEN_INV_1 U345 ( .A(n209), .X(n20) );
  SEN_OAI221_0P5 U346 ( .A1(n153), .A2(n292), .B1(n45), .B2(n288), .C(n154), 
        .X(Z[28]) );
  SEN_ND2_G_1 U347 ( .A1(n84), .A2(n173), .X(n102) );
  SEN_OAI221_1 U348 ( .A1(n232), .A2(n259), .B1(n219), .B2(n261), .C(n233), 
        .X(n224) );
  SEN_OAI221_0P5 U349 ( .A1(n201), .A2(n291), .B1(n55), .B2(n289), .C(n202), 
        .X(Z[19]) );
  SEN_EO2_S_0P5 U350 ( .A1(n251), .A2(shift_cg[1]), .X(n130) );
  SEN_OAI21_S_3 U351 ( .A1(shift_cg[3]), .A2(n253), .B(left_cg), .X(n254) );
  SEN_ND2_S_0P5 U352 ( .A1(n286), .A2(n20), .X(n267) );
  SEN_OAI221_0P5 U353 ( .A1(n213), .A2(n291), .B1(n58), .B2(n289), .C(n214), 
        .X(Z[16]) );
  SEN_INV_1 U354 ( .A(n290), .X(n289) );
  SEN_INV_0P65 U355 ( .A(n290), .X(n288) );
  SEN_INV_S_0P5 U356 ( .A(n281), .X(n292) );
  SEN_OAI222_0P5 U357 ( .A1(n125), .A2(n104), .B1(n126), .B2(n108), .C1(n127), 
        .C2(n282), .X(n110) );
  SEN_OAI222_0P5 U358 ( .A1(n120), .A2(n104), .B1(n121), .B2(n108), .C1(n122), 
        .C2(n282), .X(n99) );
  SEN_OAI22_S_0P5 U359 ( .A1(n108), .A2(n113), .B1(n258), .B2(n188), .X(n226)
         );
  SEN_OAI22_S_0P5 U360 ( .A1(n265), .A2(n193), .B1(n106), .B2(n175), .X(n215)
         );
  SEN_ND2_S_0P5 U361 ( .A1(n270), .A2(n287), .X(n238) );
  SEN_OA222_0P5 U362 ( .A1(n67), .A2(n247), .B1(n51), .B2(n248), .C1(n229), 
        .C2(n173), .X(n122) );
  SEN_OA222_0P5 U363 ( .A1(n69), .A2(n247), .B1(n53), .B2(n248), .C1(n109), 
        .C2(n173), .X(n147) );
  SEN_INV_1 U364 ( .A(n146), .X(n41) );
  SEN_OAI222_0P5 U365 ( .A1(n70), .A2(n247), .B1(n54), .B2(n248), .C1(n116), 
        .C2(n173), .X(n200) );
  SEN_AOI22_0P5 U366 ( .A1(n269), .A2(input_cg[12]), .B1(n246), .B2(
        input_cg[28]), .X(n116) );
  SEN_OAI221_0P5 U367 ( .A1(n126), .A2(n258), .B1(n127), .B2(n84), .C(n250), 
        .X(n198) );
  SEN_AOI222_0P5 U368 ( .A1(n282), .A2(n200), .B1(n244), .B2(input_cg[16]), 
        .C1(n80), .C2(n50), .X(n240) );
  SEN_ND2_2 U369 ( .A1(n277), .A2(n278), .X(n212) );
  SEN_AN2_S_0P5 U370 ( .A1(n287), .A2(n86), .X(n197) );
  SEN_AN2_S_1 U371 ( .A1(n85), .A2(n86), .X(n270) );
  SEN_ND2_0P8 U372 ( .A1(n252), .A2(n272), .X(n273) );
  SEN_INV_1 U373 ( .A(n252), .X(n271) );
  SEN_INV_S_0P5 U374 ( .A(shift_cg[3]), .X(n272) );
  SEN_ND2_T_0P5 U375 ( .A1(left_cg), .A2(n253), .X(n252) );
  SEN_ND2_S_0P5 U376 ( .A1(n246), .A2(n173), .X(n248) );
  SEN_OA222_0P5 U377 ( .A1(n68), .A2(n247), .B1(n52), .B2(n248), .C1(n232), 
        .C2(n173), .X(n127) );
  SEN_ND2_S_0P5 U378 ( .A1(n173), .A2(n282), .X(n108) );
  SEN_ND2_S_0P5 U379 ( .A1(n78), .A2(n82), .X(n158) );
  SEN_INV_1 U380 ( .A(n138), .X(n30) );
  SEN_INV_1 U381 ( .A(n148), .X(n34) );
  SEN_INV_1 U382 ( .A(n118), .X(n11) );
  SEN_INV_1 U383 ( .A(n213), .X(n8) );
  SEN_INV_1 U384 ( .A(n168), .X(n22) );
  SEN_OAI221_0P5 U385 ( .A1(n103), .A2(n102), .B1(n166), .B2(n104), .C(n206), 
        .X(n191) );
  SEN_AOI22_S_1 U386 ( .A1(n83), .A2(n23), .B1(n80), .B2(n164), .X(n206) );
  SEN_OAI221_0P5 U387 ( .A1(n203), .A2(n102), .B1(n161), .B2(n104), .C(n204), 
        .X(n186) );
  SEN_AOI22_S_1 U388 ( .A1(n83), .A2(n28), .B1(n80), .B2(n31), .X(n204) );
  SEN_OAI221_0P5 U389 ( .A1(n73), .A2(n45), .B1(n136), .B2(n62), .C(n216), .X(
        n170) );
  SEN_OAI221_0P5 U390 ( .A1(n181), .A2(n265), .B1(n161), .B2(n258), .C(n182), 
        .X(n167) );
  SEN_OAI221_0P5 U391 ( .A1(n73), .A2(n44), .B1(n136), .B2(n61), .C(n216), .X(
        n164) );
  SEN_OAI221_0P5 U392 ( .A1(n69), .A2(n137), .B1(n136), .B2(n53), .C(n39), .X(
        n144) );
  SEN_OAI221_0P5 U393 ( .A1(n68), .A2(n137), .B1(n136), .B2(n52), .C(n39), .X(
        n133) );
  SEN_AO2BB2_0P5 U394 ( .A1(n258), .A2(n166), .B1(n83), .B2(n164), .X(n185) );
  SEN_OAI221_0P5 U395 ( .A1(n73), .A2(n40), .B1(n136), .B2(n59), .C(n216), .X(
        n178) );
  SEN_NR2_S_0P5 U396 ( .A1(n136), .A2(n173), .X(n160) );
  SEN_OAI221_0P5 U397 ( .A1(n70), .A2(n137), .B1(n136), .B2(n54), .C(n39), .X(
        n171) );
  SEN_ND2_G_1 U398 ( .A1(n282), .A2(n82), .X(n104) );
  SEN_AOI222_0P5 U399 ( .A1(n84), .A2(n142), .B1(n81), .B2(n143), .C1(n83), 
        .C2(n144), .X(n141) );
  SEN_OAI221_0P5 U400 ( .A1(n61), .A2(n137), .B1(n136), .B2(n44), .C(n39), .X(
        n143) );
  SEN_OAI221_0P5 U401 ( .A1(n138), .A2(n292), .B1(n42), .B2(n288), .C(n139), 
        .X(Z[30]) );
  SEN_INV_S_0P5 U402 ( .A(n227), .X(n19) );
  SEN_INV_S_0P5 U403 ( .A(n221), .X(n14) );
  SEN_INV_S_0P5 U404 ( .A(n224), .X(n3) );
  SEN_INV_S_0P5 U405 ( .A(n117), .X(n25) );
  SEN_INV_S_0P5 U406 ( .A(n110), .X(n6) );
  SEN_INV_S_0P5 U407 ( .A(n186), .X(n5) );
  SEN_INV_S_0P5 U408 ( .A(n191), .X(n21) );
  SEN_INV_S_0P5 U409 ( .A(n195), .X(n9) );
  SEN_INV_S_0P5 U410 ( .A(n92), .X(n2) );
  SEN_INV_S_0P5 U411 ( .A(n99), .X(n18) );
  SEN_INV_S_0P5 U412 ( .A(n183), .X(n16) );
  SEN_INV_S_0P5 U413 ( .A(n95), .X(n26) );
  SEN_INV_S_0P5 U414 ( .A(n97), .X(n12) );
  SEN_INV_1 U415 ( .A(n190), .X(n37) );
  SEN_NR3_0P5 U416 ( .A1(log_cg), .A2(left_cg), .A3(n40), .X(n152) );
  SEN_AOI221_0P5 U417 ( .A1(n220), .A2(input_cg[27]), .B1(n74), .B2(
        input_cg[11]), .C(n32), .X(n175) );
  SEN_AOI221_0P5 U418 ( .A1(n220), .A2(input_cg[23]), .B1(n74), .B2(
        input_cg[7]), .C(n32), .X(n193) );
  SEN_AOI221_0P5 U419 ( .A1(n220), .A2(input_cg[20]), .B1(n74), .B2(
        input_cg[4]), .C(n32), .X(n113) );
  SEN_AOI221_0P5 U420 ( .A1(n269), .A2(input_cg[21]), .B1(n260), .B2(
        input_cg[5]), .C(n32), .X(n103) );
  SEN_AOI221_0P5 U421 ( .A1(n220), .A2(input_cg[22]), .B1(n260), .B2(
        input_cg[6]), .C(n32), .X(n203) );
  SEN_AOI221_0P5 U422 ( .A1(n220), .A2(input_cg[18]), .B1(n74), .B2(
        input_cg[2]), .C(n32), .X(n125) );
  SEN_AOI221_0P5 U423 ( .A1(n269), .A2(input_cg[19]), .B1(n260), .B2(
        input_cg[3]), .C(n32), .X(n120) );
  SEN_AOI221_0P5 U424 ( .A1(input_cg[30]), .A2(n220), .B1(input_cg[14]), .B2(
        n74), .C(n32), .X(n181) );
  SEN_AOI221_0P5 U425 ( .A1(n269), .A2(input_cg[25]), .B1(n74), .B2(
        input_cg[9]), .C(n32), .X(n207) );
  SEN_AOI221_0P5 U426 ( .A1(input_cg[3]), .A2(n78), .B1(n260), .B2(
        input_cg[19]), .C(n152), .X(n155) );
  SEN_AOI221_0P5 U427 ( .A1(n269), .A2(input_cg[17]), .B1(n260), .B2(
        input_cg[1]), .C(n32), .X(n107) );
  SEN_AOI221_0P5 U428 ( .A1(input_cg[28]), .A2(n260), .B1(n78), .B2(
        input_cg[12]), .C(n152), .X(n150) );
  SEN_INV_S_0P5 U429 ( .A(n151), .X(n36) );
  SEN_AOI221_0P5 U430 ( .A1(input_cg[27]), .A2(n260), .B1(n78), .B2(
        input_cg[11]), .C(n152), .X(n156) );
  SEN_AOI221_0P5 U431 ( .A1(n269), .A2(input_cg[26]), .B1(n260), .B2(
        input_cg[10]), .C(n32), .X(n219) );
  SEN_AOI22_0P5 U432 ( .A1(n269), .A2(input_cg[15]), .B1(n246), .B2(
        input_cg[31]), .X(n229) );
  SEN_AOI22_0P5 U433 ( .A1(n269), .A2(input_cg[13]), .B1(n246), .B2(
        input_cg[29]), .X(n109) );
  SEN_AOI22_0P5 U434 ( .A1(n269), .A2(input_cg[11]), .B1(n246), .B2(
        input_cg[27]), .X(n121) );
  SEN_AOI22_0P5 U435 ( .A1(n269), .A2(input_cg[10]), .B1(n246), .B2(
        input_cg[26]), .X(n126) );
  SEN_AOI22_0P5 U436 ( .A1(n269), .A2(input_cg[9]), .B1(n246), .B2(
        input_cg[25]), .X(n101) );
  SEN_AOI22_0P5 U437 ( .A1(n269), .A2(input_cg[14]), .B1(n246), .B2(
        input_cg[30]), .X(n232) );
  SEN_AOI22_0P5 U438 ( .A1(n269), .A2(input_cg[8]), .B1(n246), .B2(
        input_cg[24]), .X(n112) );
  SEN_OAI222_0P5 U439 ( .A1(shift_cg[0]), .A2(n128), .B1(n129), .B2(n86), .C1(
        n40), .C2(n289), .X(Z[31]) );
  SEN_OA2BB2_0P5 U440 ( .A1(n130), .A2(n131), .B1(n130), .B2(n132), .X(n129)
         );
  SEN_AOI222_0P5 U441 ( .A1(n133), .A2(n83), .B1(n134), .B2(n81), .C1(n135), 
        .C2(n84), .X(n132) );
  SEN_OAI221_0P5 U442 ( .A1(n136), .A2(n42), .B1(n137), .B2(n60), .C(n39), .X(
        n134) );
  SEN_INV_S_0P5 U443 ( .A(n162), .X(n29) );
  SEN_INV_S_0P5 U444 ( .A(n167), .X(n27) );
  SEN_INV_S_0P5 U445 ( .A(n90), .X(n13) );
  SEN_INV_S_0P5 U446 ( .A(n208), .X(n4) );
  SEN_INV_S_0P5 U447 ( .A(n179), .X(n10) );
  SEN_AOI22_0P5 U448 ( .A1(shift_cg[0]), .A2(n196), .B1(n290), .B2(input_cg[0]), .X(n241) );
  SEN_INV_S_0P5 U449 ( .A(shift_cg[0]), .X(n86) );
  SEN_NR2B_V1_1 U450 ( .A(left_cg), .B(n255), .X(n256) );
  SEN_INV_1 U451 ( .A(n176), .X(n35) );
  SEN_AO221_0P5 U452 ( .A1(n269), .A2(input_cg[16]), .B1(n260), .B2(
        input_cg[0]), .C(n32), .X(n115) );
  SEN_AOI221_1 U453 ( .A1(input_cg[0]), .A2(n78), .B1(n74), .B2(input_cg[16]), 
        .C(n152), .X(n190) );
  SEN_NR2_S_4 U454 ( .A1(shift_cg[1]), .A2(shift_cg[0]), .X(n255) );
  SEN_NR2_S_0P5 U455 ( .A1(n212), .A2(left_cg), .X(n246) );
  SEN_INV_S_1 U456 ( .A(n238), .X(n294) );
  SEN_INV_S_1 U457 ( .A(n238), .X(n293) );
  SEN_NR2_1 U458 ( .A1(n102), .A2(n73), .X(n243) );
  SEN_INV_S_1 U459 ( .A(n171), .X(n38) );
  SEN_INV_S_1 U460 ( .A(n280), .X(n283) );
  SEN_INV_S_1 U461 ( .A(n279), .X(n286) );
  SEN_INV_S_1 U462 ( .A(n279), .X(n285) );
  SEN_INV_S_1 U463 ( .A(n280), .X(n284) );
  SEN_OAI221_1 U464 ( .A1(n188), .A2(n259), .B1(n38), .B2(n261), .C(n189), .X(
        n179) );
  SEN_AOI22_1 U465 ( .A1(n83), .A2(n170), .B1(n80), .B2(n37), .X(n189) );
  SEN_OAI221_1 U466 ( .A1(n193), .A2(n102), .B1(n155), .B2(n104), .C(n194), 
        .X(n183) );
  SEN_OA2BB2_1 U467 ( .A1(n80), .A2(n178), .B1(n265), .B2(n175), .X(n194) );
  SEN_OA2BB2_1 U468 ( .A1(n80), .A2(n170), .B1(n265), .B2(n188), .X(n211) );
  SEN_OAI221_1 U469 ( .A1(n125), .A2(n259), .B1(n181), .B2(n261), .C(n218), 
        .X(n208) );
  SEN_OA2BB2_1 U470 ( .A1(n80), .A2(n28), .B1(n265), .B2(n203), .X(n218) );
  SEN_OAI221_1 U471 ( .A1(n101), .A2(n102), .B1(n103), .B2(n104), .C(n105), 
        .X(n95) );
  SEN_OA22_1 U472 ( .A1(n258), .A2(n107), .B1(n265), .B2(n109), .X(n105) );
  SEN_OAI221_1 U473 ( .A1(n126), .A2(n102), .B1(n203), .B2(n104), .C(n239), 
        .X(n92) );
  SEN_OA22_1 U474 ( .A1(n258), .A2(n125), .B1(n265), .B2(n232), .X(n239) );
  SEN_OAI221_1 U475 ( .A1(n121), .A2(n102), .B1(n193), .B2(n104), .C(n236), 
        .X(n90) );
  SEN_OA22_1 U476 ( .A1(n258), .A2(n120), .B1(n265), .B2(n229), .X(n236) );
  SEN_OAI221_1 U477 ( .A1(n116), .A2(n102), .B1(n188), .B2(n104), .C(n237), 
        .X(n94) );
  SEN_OA2BB2_1 U478 ( .A1(n83), .A2(n115), .B1(n258), .B2(n113), .X(n237) );
  SEN_OAI221_1 U479 ( .A1(n109), .A2(n259), .B1(n207), .B2(n261), .C(n235), 
        .X(n227) );
  SEN_OA2BB2_1 U480 ( .A1(n83), .A2(n24), .B1(n258), .B2(n103), .X(n235) );
  SEN_OA22_1 U481 ( .A1(n258), .A2(n203), .B1(n265), .B2(n125), .X(n233) );
  SEN_OAI221_1 U482 ( .A1(n229), .A2(n259), .B1(n175), .B2(n104), .C(n230), 
        .X(n221) );
  SEN_OA22_1 U483 ( .A1(n265), .A2(n120), .B1(n258), .B2(n193), .X(n230) );
  SEN_OAI221_1 U484 ( .A1(n112), .A2(n102), .B1(n113), .B2(n104), .C(n114), 
        .X(n97) );
  SEN_OA2BB2_1 U485 ( .A1(n80), .A2(n115), .B1(n265), .B2(n116), .X(n114) );
  SEN_INV_S_0P5 U486 ( .A(n173), .X(n82) );
  SEN_AOI221_1 U487 ( .A1(n115), .A2(n79), .B1(n170), .B2(n81), .C(n226), .X(
        n213) );
  SEN_AOI221_1 U488 ( .A1(n24), .A2(n79), .B1(n164), .B2(n81), .C(n223), .X(
        n209) );
  SEN_OAI22_1 U489 ( .A1(n265), .A2(n103), .B1(n258), .B2(n207), .X(n223) );
  SEN_AOI221_1 U490 ( .A1(n17), .A2(n79), .B1(n178), .B2(n81), .C(n215), .X(
        n201) );
  SEN_AOI221_1 U491 ( .A1(n23), .A2(n79), .B1(n144), .B2(n81), .C(n185), .X(
        n168) );
  SEN_AOI222_1 U492 ( .A1(n115), .A2(n81), .B1(n50), .B2(n83), .C1(n200), .C2(
        n84), .X(n118) );
  SEN_AOI222_1 U493 ( .A1(n31), .A2(n79), .B1(n133), .B2(n80), .C1(n135), .C2(
        n282), .X(n138) );
  SEN_AOI222_1 U494 ( .A1(n164), .A2(n79), .B1(n144), .B2(n80), .C1(n142), 
        .C2(n282), .X(n148) );
  SEN_OAI221_1 U495 ( .A1(n118), .A2(n292), .B1(n70), .B2(n288), .C(n119), .X(
        Z[4]) );
  SEN_AOI222_1 U496 ( .A1(n293), .A2(n110), .B1(n285), .B2(n117), .C1(n283), 
        .C2(n99), .X(n119) );
  SEN_OAI221_1 U497 ( .A1(n25), .A2(n292), .B1(n69), .B2(n288), .C(n111), .X(
        Z[5]) );
  SEN_AOI222_1 U498 ( .A1(n293), .A2(n99), .B1(n285), .B2(n110), .C1(n283), 
        .C2(n97), .X(n111) );
  SEN_OA2BB2_1 U499 ( .A1(n140), .A2(n130), .B1(n141), .B2(n130), .X(n128) );
  SEN_OAI221_1 U500 ( .A1(n148), .A2(n292), .B1(n44), .B2(n288), .C(n149), .X(
        Z[29]) );
  SEN_AOI222_1 U501 ( .A1(n293), .A2(n140), .B1(n285), .B2(n30), .C1(n283), 
        .C2(n131), .X(n149) );
  SEN_AOI222_1 U502 ( .A1(n293), .A2(n30), .B1(n285), .B2(n34), .C1(n283), 
        .C2(n140), .X(n154) );
  SEN_INV_S_1 U503 ( .A(n130), .X(n85) );
  SEN_OAI221_1 U504 ( .A1(n6), .A2(n292), .B1(n68), .B2(n288), .C(n100), .X(
        Z[6]) );
  SEN_AOI222_1 U505 ( .A1(n293), .A2(n97), .B1(n285), .B2(n99), .C1(n283), 
        .C2(n95), .X(n100) );
  SEN_OAI221_1 U506 ( .A1(n18), .A2(n292), .B1(n67), .B2(n288), .C(n98), .X(
        Z[7]) );
  SEN_AOI222_1 U507 ( .A1(n293), .A2(n95), .B1(n285), .B2(n97), .C1(n283), 
        .C2(n92), .X(n98) );
  SEN_INV_1 U508 ( .A(n181), .X(n31) );
  SEN_OAI221_1 U509 ( .A1(n9), .A2(n291), .B1(n54), .B2(n289), .C(n192), .X(
        Z[20]) );
  SEN_AOI222_1 U510 ( .A1(n294), .A2(n186), .B1(n286), .B2(n191), .C1(n284), 
        .C2(n183), .X(n192) );
  SEN_OAI221_1 U511 ( .A1(n21), .A2(n291), .B1(n53), .B2(n289), .C(n187), .X(
        Z[21]) );
  SEN_AOI222_1 U512 ( .A1(n294), .A2(n183), .B1(n286), .B2(n186), .C1(n284), 
        .C2(n179), .X(n187) );
  SEN_AOI222_1 U513 ( .A1(n294), .A2(n22), .B1(n286), .B2(n179), .C1(n284), 
        .C2(n167), .X(n180) );
  SEN_OAI221_1 U514 ( .A1(n5), .A2(n291), .B1(n52), .B2(n289), .C(n184), .X(
        Z[22]) );
  SEN_AOI222_1 U515 ( .A1(n294), .A2(n179), .B1(n286), .B2(n183), .C1(n284), 
        .C2(n22), .X(n184) );
  SEN_OAI221_1 U516 ( .A1(n26), .A2(n291), .B1(n65), .B2(n289), .C(n89), .X(
        Z[9]) );
  SEN_AOI222_1 U517 ( .A1(n294), .A2(n90), .B1(n286), .B2(n92), .C1(n284), 
        .C2(n94), .X(n89) );
  SEN_OAI221_1 U518 ( .A1(n2), .A2(n291), .B1(n64), .B2(n288), .C(n234), .X(
        Z[10]) );
  SEN_AOI222_1 U519 ( .A1(n293), .A2(n94), .B1(n285), .B2(n90), .C1(n283), 
        .C2(n227), .X(n234) );
  SEN_OAI221_1 U520 ( .A1(n7), .A2(n291), .B1(n62), .B2(n289), .C(n228), .X(
        Z[12]) );
  SEN_INV_S_1 U521 ( .A(n94), .X(n7) );
  SEN_AOI222_1 U522 ( .A1(n294), .A2(n224), .B1(n285), .B2(n227), .C1(n284), 
        .C2(n221), .X(n228) );
  SEN_OAI221_1 U523 ( .A1(n19), .A2(n291), .B1(n61), .B2(n289), .C(n225), .X(
        Z[13]) );
  SEN_AOI222_1 U524 ( .A1(n294), .A2(n221), .B1(n286), .B2(n224), .C1(n284), 
        .C2(n8), .X(n225) );
  SEN_OAI221_1 U525 ( .A1(n3), .A2(n291), .B1(n60), .B2(n289), .C(n222), .X(
        Z[14]) );
  SEN_AOI222_1 U526 ( .A1(n294), .A2(n8), .B1(n286), .B2(n221), .C1(n283), 
        .C2(n20), .X(n222) );
  SEN_OAI221_1 U527 ( .A1(n14), .A2(n291), .B1(n59), .B2(n289), .C(n217), .X(
        Z[15]) );
  SEN_AOI222_1 U528 ( .A1(n294), .A2(n20), .B1(n286), .B2(n8), .C1(n284), .C2(
        n208), .X(n217) );
  SEN_OAI221_1 U529 ( .A1(n12), .A2(n292), .B1(n66), .B2(n288), .C(n96), .X(
        Z[8]) );
  SEN_AOI222_1 U530 ( .A1(n293), .A2(n92), .B1(n285), .B2(n95), .C1(n283), 
        .C2(n90), .X(n96) );
  SEN_INV_1 U531 ( .A(n219), .X(n28) );
  SEN_INV_S_1 U532 ( .A(n220), .X(n73) );
  SEN_INV_1 U533 ( .A(n207), .X(n23) );
  SEN_INV_S_1 U534 ( .A(n152), .X(n39) );
  SEN_INV_1 U535 ( .A(n107), .X(n24) );
  SEN_OA2BB2_1 U536 ( .A1(n293), .A2(n131), .B1(n86), .B2(n128), .X(n139) );
  SEN_OR2_1 U537 ( .A1(n85), .A2(n86), .X(n279) );
  SEN_OR2_1 U538 ( .A1(n86), .A2(n130), .X(n280) );
  SEN_INV_S_1 U539 ( .A(n198), .X(n43) );
  SEN_INV_S_1 U540 ( .A(n112), .X(n50) );
  SEN_INV_1 U541 ( .A(n257), .X(n287) );
  SEN_OAI222_1 U542 ( .A1(n155), .A2(n265), .B1(n156), .B2(n104), .C1(n35), 
        .C2(n282), .X(n140) );
  SEN_OAI222_1 U543 ( .A1(n38), .A2(n265), .B1(n150), .B2(n261), .C1(n36), 
        .C2(n282), .X(n131) );
  SEN_AOI221_1 U544 ( .A1(input_cg[1]), .A2(n78), .B1(n260), .B2(input_cg[17]), 
        .C(n152), .X(n166) );
  SEN_AOI221_1 U545 ( .A1(input_cg[2]), .A2(n78), .B1(input_cg[18]), .B2(n260), 
        .C(n152), .X(n161) );
  SEN_ND2_S_0P5 U546 ( .A1(shift_cg[0]), .A2(left_cg), .X(n251) );
  SEN_AOI22_1 U547 ( .A1(n243), .A2(input_cg[3]), .B1(n244), .B2(input_cg[19]), 
        .X(n249) );
  SEN_OAI211_1 U548 ( .A1(n64), .A2(n158), .B1(n39), .B2(n159), .X(n135) );
  SEN_OA2BB2_1 U549 ( .A1(n160), .A2(input_cg[26]), .B1(n82), .B2(n161), .X(
        n159) );
  SEN_OAI211_1 U550 ( .A1(n65), .A2(n158), .B1(n39), .B2(n165), .X(n142) );
  SEN_OA2BB2_1 U551 ( .A1(n160), .A2(input_cg[25]), .B1(n82), .B2(n166), .X(
        n165) );
  SEN_AOI22_1 U552 ( .A1(n243), .A2(input_cg[2]), .B1(n244), .B2(input_cg[18]), 
        .X(n250) );
  SEN_OAI221_1 U553 ( .A1(n41), .A2(n292), .B1(n71), .B2(n288), .C(n124), .X(
        Z[3]) );
  SEN_INV_S_1 U554 ( .A(input_cg[3]), .X(n71) );
  SEN_AOI222_1 U555 ( .A1(n293), .A2(n117), .B1(n285), .B2(n11), .C1(n283), 
        .C2(n110), .X(n124) );
  SEN_OAI211_1 U556 ( .A1(n67), .A2(n158), .B1(n39), .B2(n177), .X(n176) );
  SEN_ND2_G_1 U557 ( .A1(n75), .A2(left_cg), .X(n136) );
  SEN_OAI22_1 U558 ( .A1(n41), .A2(n130), .B1(n242), .B2(n85), .X(n196) );
  SEN_AOI221_1 U559 ( .A1(n243), .A2(input_cg[1]), .B1(n244), .B2(input_cg[17]), .C(n245), .X(n242) );
  SEN_INV_S_1 U560 ( .A(input_cg[16]), .X(n58) );
  SEN_OAI221_1 U561 ( .A1(n209), .A2(n291), .B1(n57), .B2(n289), .C(n210), .X(
        Z[17]) );
  SEN_INV_S_1 U562 ( .A(input_cg[17]), .X(n57) );
  SEN_AOI222_1 U563 ( .A1(n294), .A2(n15), .B1(n286), .B2(n208), .C1(n284), 
        .C2(n195), .X(n210) );
  SEN_OAI221_1 U564 ( .A1(n168), .A2(n292), .B1(n48), .B2(n288), .C(n169), .X(
        Z[25]) );
  SEN_INV_S_1 U565 ( .A(input_cg[25]), .X(n48) );
  SEN_AOI222_1 U566 ( .A1(n293), .A2(n162), .B1(n285), .B2(n167), .C1(n283), 
        .C2(n33), .X(n169) );
  SEN_INV_S_1 U567 ( .A(input_cg[19]), .X(n55) );
  SEN_AOI222_1 U568 ( .A1(n294), .A2(n191), .B1(n286), .B2(n195), .C1(n284), 
        .C2(n186), .X(n202) );
  SEN_OAI221_1 U569 ( .A1(n240), .A2(n291), .B1(n43), .B2(n238), .C(n241), .X(
        Z[0]) );
  SEN_OAI221_1 U570 ( .A1(n29), .A2(n292), .B1(n46), .B2(n288), .C(n157), .X(
        Z[27]) );
  SEN_INV_S_1 U571 ( .A(input_cg[27]), .X(n46) );
  SEN_AOI222_1 U572 ( .A1(n293), .A2(n34), .B1(n285), .B2(n33), .C1(n283), 
        .C2(n30), .X(n157) );
  SEN_OAI221_1 U573 ( .A1(n10), .A2(n292), .B1(n49), .B2(n289), .C(n174), .X(
        Z[24]) );
  SEN_INV_S_1 U574 ( .A(input_cg[24]), .X(n49) );
  SEN_AOI222_1 U575 ( .A1(n294), .A2(n167), .B1(n286), .B2(n22), .C1(n284), 
        .C2(n162), .X(n174) );
  SEN_OAI221_1 U576 ( .A1(n27), .A2(n292), .B1(n47), .B2(n288), .C(n163), .X(
        Z[26]) );
  SEN_INV_S_1 U577 ( .A(input_cg[26]), .X(n47) );
  SEN_AOI222_1 U578 ( .A1(n293), .A2(n33), .B1(n285), .B2(n162), .C1(n283), 
        .C2(n34), .X(n163) );
  SEN_OAI221_1 U579 ( .A1(n4), .A2(n291), .B1(n56), .B2(n289), .C(n205), .X(
        Z[18]) );
  SEN_INV_S_1 U580 ( .A(input_cg[18]), .X(n56) );
  SEN_AOI222_1 U581 ( .A1(n294), .A2(n195), .B1(n286), .B2(n15), .C1(n284), 
        .C2(n191), .X(n205) );
  SEN_OAI221_1 U582 ( .A1(n13), .A2(n291), .B1(n63), .B2(n288), .C(n231), .X(
        Z[11]) );
  SEN_INV_S_1 U583 ( .A(input_cg[11]), .X(n63) );
  SEN_AOI222_1 U584 ( .A1(n294), .A2(n227), .B1(n285), .B2(n94), .C1(n284), 
        .C2(n224), .X(n231) );
  SEN_OAI221_1 U585 ( .A1(n43), .A2(n292), .B1(n72), .B2(n288), .C(n145), .X(
        Z[2]) );
  SEN_INV_S_1 U586 ( .A(input_cg[2]), .X(n72) );
  SEN_EO2_S_0P5 U587 ( .A1(shift_cg[2]), .A2(n256), .X(n123) );
  SEN_INV_S_1 U588 ( .A(input_cg[31]), .X(n40) );
  SEN_INV_S_1 U589 ( .A(input_cg[29]), .X(n44) );
  SEN_INV_S_1 U590 ( .A(input_cg[13]), .X(n61) );
  SEN_INV_S_1 U591 ( .A(input_cg[20]), .X(n54) );
  SEN_INV_S_1 U592 ( .A(input_cg[4]), .X(n70) );
  SEN_INV_S_1 U593 ( .A(input_cg[21]), .X(n53) );
  SEN_INV_S_1 U594 ( .A(input_cg[22]), .X(n52) );
  SEN_INV_S_1 U595 ( .A(input_cg[7]), .X(n67) );
  SEN_INV_S_1 U596 ( .A(input_cg[5]), .X(n69) );
  SEN_INV_S_1 U597 ( .A(input_cg[6]), .X(n68) );
  SEN_INV_S_1 U598 ( .A(input_cg[12]), .X(n62) );
  SEN_INV_S_1 U599 ( .A(input_cg[28]), .X(n45) );
  SEN_INV_S_1 U600 ( .A(input_cg[30]), .X(n42) );
  SEN_INV_S_1 U601 ( .A(input_cg[14]), .X(n60) );
  SEN_INV_S_1 U602 ( .A(input_cg[9]), .X(n65) );
  SEN_INV_S_1 U603 ( .A(input_cg[8]), .X(n66) );
  SEN_INV_S_1 U604 ( .A(input_cg[10]), .X(n64) );
  SEN_INV_S_1 U605 ( .A(input_cg[15]), .X(n59) );
  SEN_INV_S_1 U606 ( .A(input_cg[23]), .X(n51) );
  SEN_AO221_1 U607 ( .A1(n196), .A2(n197), .B1(n198), .B2(n286), .C(n199), .X(
        Z[1]) );
  SEN_AO22_1 U608 ( .A1(n284), .A2(n11), .B1(n290), .B2(input_cg[1]), .X(n199)
         );
  SEN_FDPQ_D_1 \shift_cg_reg[1]  ( .D(S[1]), .CK(clock), .Q(shift_cg[1]) );
endmodule

