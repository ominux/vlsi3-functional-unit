
module Alu ( Z, A, B, INST, SEL );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  input SEL;
  wire   adder_cin, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n216,
         n217, \struct_adder/add_1_root_add_19_2/carry[31] ,
         \struct_adder/add_1_root_add_19_2/carry[30] ,
         \struct_adder/add_1_root_add_19_2/carry[29] ,
         \struct_adder/add_1_root_add_19_2/carry[28] ,
         \struct_adder/add_1_root_add_19_2/carry[27] ,
         \struct_adder/add_1_root_add_19_2/carry[26] ,
         \struct_adder/add_1_root_add_19_2/carry[25] ,
         \struct_adder/add_1_root_add_19_2/carry[24] ,
         \struct_adder/add_1_root_add_19_2/carry[23] ,
         \struct_adder/add_1_root_add_19_2/carry[22] ,
         \struct_adder/add_1_root_add_19_2/carry[21] ,
         \struct_adder/add_1_root_add_19_2/carry[20] ,
         \struct_adder/add_1_root_add_19_2/carry[19] ,
         \struct_adder/add_1_root_add_19_2/carry[18] ,
         \struct_adder/add_1_root_add_19_2/carry[17] ,
         \struct_adder/add_1_root_add_19_2/carry[16] ,
         \struct_adder/add_1_root_add_19_2/carry[15] ,
         \struct_adder/add_1_root_add_19_2/carry[14] ,
         \struct_adder/add_1_root_add_19_2/carry[13] ,
         \struct_adder/add_1_root_add_19_2/carry[12] ,
         \struct_adder/add_1_root_add_19_2/carry[11] ,
         \struct_adder/add_1_root_add_19_2/carry[10] ,
         \struct_adder/add_1_root_add_19_2/carry[9] ,
         \struct_adder/add_1_root_add_19_2/carry[8] ,
         \struct_adder/add_1_root_add_19_2/carry[7] ,
         \struct_adder/add_1_root_add_19_2/carry[6] ,
         \struct_adder/add_1_root_add_19_2/carry[5] ,
         \struct_adder/add_1_root_add_19_2/carry[4] ,
         \struct_adder/add_1_root_add_19_2/carry[3] ,
         \struct_adder/add_1_root_add_19_2/carry[2] ,
         \struct_adder/add_1_root_add_19_2/carry[1] , n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330;
  wire   [31:0] adder_a;
  wire   [31:0] adder_b;
  wire   [31:0] adder_out;

  SEN_LDPQ_D_1 adder_cin_reg ( .G(N188), .D(N189), .Q(adder_cin) );
  SEN_LDPQ_D_1 \adder_b_reg[30]  ( .G(n255), .D(N186), .Q(adder_b[30]) );
  SEN_LDPQ_D_1 \adder_b_reg[29]  ( .G(n255), .D(N185), .Q(adder_b[29]) );
  SEN_LDPQ_D_1 \adder_b_reg[28]  ( .G(n255), .D(N184), .Q(adder_b[28]) );
  SEN_LDPQ_D_1 \adder_b_reg[27]  ( .G(n255), .D(N183), .Q(adder_b[27]) );
  SEN_LDPQ_D_1 \adder_b_reg[26]  ( .G(n255), .D(N182), .Q(adder_b[26]) );
  SEN_LDPQ_D_1 \adder_b_reg[25]  ( .G(n255), .D(N181), .Q(adder_b[25]) );
  SEN_LDPQ_D_1 \adder_b_reg[24]  ( .G(n255), .D(N180), .Q(adder_b[24]) );
  SEN_LDPQ_D_1 \adder_b_reg[23]  ( .G(n255), .D(N179), .Q(adder_b[23]) );
  SEN_LDPQ_D_1 \adder_b_reg[22]  ( .G(n255), .D(N178), .Q(adder_b[22]) );
  SEN_LDPQ_D_1 \adder_b_reg[21]  ( .G(n255), .D(N177), .Q(adder_b[21]) );
  SEN_LDPQ_D_1 \adder_b_reg[20]  ( .G(n255), .D(N176), .Q(adder_b[20]) );
  SEN_LDPQ_D_1 \adder_b_reg[19]  ( .G(n255), .D(N175), .Q(adder_b[19]) );
  SEN_LDPQ_D_1 \adder_b_reg[18]  ( .G(n256), .D(N174), .Q(adder_b[18]) );
  SEN_LDPQ_D_1 \adder_b_reg[17]  ( .G(n256), .D(N173), .Q(adder_b[17]) );
  SEN_LDPQ_D_1 \adder_b_reg[16]  ( .G(n256), .D(N172), .Q(adder_b[16]) );
  SEN_LDPQ_D_1 \adder_b_reg[15]  ( .G(n256), .D(N171), .Q(adder_b[15]) );
  SEN_LDPQ_D_1 \adder_b_reg[14]  ( .G(n256), .D(N170), .Q(adder_b[14]) );
  SEN_LDPQ_D_1 \adder_b_reg[13]  ( .G(n256), .D(N169), .Q(adder_b[13]) );
  SEN_LDPQ_D_1 \adder_b_reg[12]  ( .G(n256), .D(N168), .Q(adder_b[12]) );
  SEN_LDPQ_D_1 \adder_b_reg[11]  ( .G(n256), .D(N167), .Q(adder_b[11]) );
  SEN_LDPQ_D_1 \adder_b_reg[10]  ( .G(n256), .D(N166), .Q(adder_b[10]) );
  SEN_LDPQ_D_1 \adder_b_reg[9]  ( .G(n256), .D(N165), .Q(adder_b[9]) );
  SEN_LDPQ_D_1 \adder_b_reg[8]  ( .G(n256), .D(N164), .Q(adder_b[8]) );
  SEN_LDPQ_D_1 \adder_b_reg[7]  ( .G(n256), .D(N163), .Q(adder_b[7]) );
  SEN_LDPQ_D_1 \adder_b_reg[6]  ( .G(n256), .D(N162), .Q(adder_b[6]) );
  SEN_LDPQ_D_1 \adder_b_reg[5]  ( .G(n256), .D(N161), .Q(adder_b[5]) );
  SEN_LDPQ_D_1 \adder_b_reg[4]  ( .G(n256), .D(N160), .Q(adder_b[4]) );
  SEN_LDPQ_D_1 \adder_b_reg[3]  ( .G(N188), .D(N159), .Q(adder_b[3]) );
  SEN_LDPQ_D_1 \adder_b_reg[2]  ( .G(N188), .D(N158), .Q(adder_b[2]) );
  SEN_LDPQ_D_1 \adder_b_reg[1]  ( .G(N188), .D(N157), .Q(adder_b[1]) );
  SEN_LDPQ_D_1 \adder_b_reg[0]  ( .G(N188), .D(N156), .Q(adder_b[0]) );
  SEN_LDPQ_D_1 \adder_a_reg[30]  ( .G(n253), .D(N154), .Q(adder_a[30]) );
  SEN_LDPQ_D_1 \adder_a_reg[29]  ( .G(n253), .D(N153), .Q(adder_a[29]) );
  SEN_LDPQ_D_1 \adder_a_reg[28]  ( .G(n253), .D(N152), .Q(adder_a[28]) );
  SEN_LDPQ_D_1 \adder_a_reg[27]  ( .G(n253), .D(N151), .Q(adder_a[27]) );
  SEN_LDPQ_D_1 \adder_a_reg[26]  ( .G(n253), .D(N150), .Q(adder_a[26]) );
  SEN_LDPQ_D_1 \adder_a_reg[25]  ( .G(n253), .D(N149), .Q(adder_a[25]) );
  SEN_LDPQ_D_1 \adder_a_reg[24]  ( .G(n253), .D(N148), .Q(adder_a[24]) );
  SEN_LDPQ_D_1 \adder_a_reg[23]  ( .G(n253), .D(N147), .Q(adder_a[23]) );
  SEN_LDPQ_D_1 \adder_a_reg[22]  ( .G(n253), .D(N146), .Q(adder_a[22]) );
  SEN_LDPQ_D_1 \adder_a_reg[21]  ( .G(n253), .D(N145), .Q(adder_a[21]) );
  SEN_LDPQ_D_1 \adder_a_reg[20]  ( .G(n253), .D(N144), .Q(adder_a[20]) );
  SEN_LDPQ_D_1 \adder_a_reg[19]  ( .G(n253), .D(N143), .Q(adder_a[19]) );
  SEN_LDPQ_D_1 \adder_a_reg[18]  ( .G(n253), .D(N142), .Q(adder_a[18]) );
  SEN_LDPQ_D_1 \adder_a_reg[17]  ( .G(n253), .D(N141), .Q(adder_a[17]) );
  SEN_LDPQ_D_1 \adder_a_reg[16]  ( .G(n254), .D(N140), .Q(adder_a[16]) );
  SEN_LDPQ_D_1 \adder_a_reg[15]  ( .G(n254), .D(N139), .Q(adder_a[15]) );
  SEN_LDPQ_D_1 \adder_a_reg[14]  ( .G(n254), .D(N138), .Q(adder_a[14]) );
  SEN_LDPQ_D_1 \adder_a_reg[13]  ( .G(n254), .D(N137), .Q(adder_a[13]) );
  SEN_LDPQ_D_1 \adder_a_reg[12]  ( .G(n254), .D(N136), .Q(adder_a[12]) );
  SEN_LDPQ_D_1 \adder_a_reg[11]  ( .G(n254), .D(N135), .Q(adder_a[11]) );
  SEN_LDPQ_D_1 \adder_a_reg[10]  ( .G(n254), .D(N134), .Q(adder_a[10]) );
  SEN_LDPQ_D_1 \adder_a_reg[9]  ( .G(n254), .D(N133), .Q(adder_a[9]) );
  SEN_LDPQ_D_1 \adder_a_reg[8]  ( .G(n254), .D(N132), .Q(adder_a[8]) );
  SEN_LDPQ_D_1 \adder_a_reg[7]  ( .G(n254), .D(N131), .Q(adder_a[7]) );
  SEN_LDPQ_D_1 \adder_a_reg[6]  ( .G(n254), .D(N130), .Q(adder_a[6]) );
  SEN_LDPQ_D_1 \adder_a_reg[5]  ( .G(n254), .D(N129), .Q(adder_a[5]) );
  SEN_LDPQ_D_1 \adder_a_reg[4]  ( .G(n254), .D(N128), .Q(adder_a[4]) );
  SEN_LDPQ_D_1 \adder_a_reg[3]  ( .G(n254), .D(N127), .Q(adder_a[3]) );
  SEN_LDPQ_D_1 \adder_a_reg[2]  ( .G(n254), .D(N126), .Q(adder_a[2]) );
  SEN_LDPQ_D_1 \adder_a_reg[1]  ( .G(n255), .D(N125), .Q(adder_a[1]) );
  SEN_LDPQ_D_1 \adder_a_reg[0]  ( .G(n255), .D(N124), .Q(adder_a[0]) );
  SEN_LDPQ_D_1 \adder_b_reg[31]  ( .G(n255), .D(N187), .Q(adder_b[31]) );
  SEN_LDPQ_D_1 \adder_a_reg[31]  ( .G(n253), .D(N155), .Q(adder_a[31]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_30  ( .A(adder_a[30]), .B(
        adder_b[30]), .CI(\struct_adder/add_1_root_add_19_2/carry[30] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[31] ), .S(adder_out[30]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_29  ( .A(adder_a[29]), .B(
        adder_b[29]), .CI(\struct_adder/add_1_root_add_19_2/carry[29] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[30] ), .S(adder_out[29]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_28  ( .A(adder_a[28]), .B(
        adder_b[28]), .CI(\struct_adder/add_1_root_add_19_2/carry[28] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[29] ), .S(adder_out[28]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_27  ( .A(adder_a[27]), .B(
        adder_b[27]), .CI(\struct_adder/add_1_root_add_19_2/carry[27] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[28] ), .S(adder_out[27]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_26  ( .A(adder_a[26]), .B(
        adder_b[26]), .CI(\struct_adder/add_1_root_add_19_2/carry[26] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[27] ), .S(adder_out[26]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_25  ( .A(adder_a[25]), .B(
        adder_b[25]), .CI(\struct_adder/add_1_root_add_19_2/carry[25] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[26] ), .S(adder_out[25]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_24  ( .A(adder_a[24]), .B(
        adder_b[24]), .CI(\struct_adder/add_1_root_add_19_2/carry[24] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[25] ), .S(adder_out[24]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_23  ( .A(adder_a[23]), .B(
        adder_b[23]), .CI(\struct_adder/add_1_root_add_19_2/carry[23] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[24] ), .S(adder_out[23]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_22  ( .A(adder_a[22]), .B(
        adder_b[22]), .CI(\struct_adder/add_1_root_add_19_2/carry[22] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[23] ), .S(adder_out[22]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_21  ( .A(adder_a[21]), .B(
        adder_b[21]), .CI(\struct_adder/add_1_root_add_19_2/carry[21] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[22] ), .S(adder_out[21]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_20  ( .A(adder_a[20]), .B(
        adder_b[20]), .CI(\struct_adder/add_1_root_add_19_2/carry[20] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[21] ), .S(adder_out[20]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_19  ( .A(adder_a[19]), .B(
        adder_b[19]), .CI(\struct_adder/add_1_root_add_19_2/carry[19] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[20] ), .S(adder_out[19]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_18  ( .A(adder_a[18]), .B(
        adder_b[18]), .CI(\struct_adder/add_1_root_add_19_2/carry[18] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[19] ), .S(adder_out[18]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_17  ( .A(adder_a[17]), .B(
        adder_b[17]), .CI(\struct_adder/add_1_root_add_19_2/carry[17] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[18] ), .S(adder_out[17]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_16  ( .A(adder_a[16]), .B(
        adder_b[16]), .CI(\struct_adder/add_1_root_add_19_2/carry[16] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[17] ), .S(adder_out[16]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_15  ( .A(adder_a[15]), .B(
        adder_b[15]), .CI(\struct_adder/add_1_root_add_19_2/carry[15] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[16] ), .S(adder_out[15]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_14  ( .A(adder_a[14]), .B(
        adder_b[14]), .CI(\struct_adder/add_1_root_add_19_2/carry[14] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[15] ), .S(adder_out[14]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_13  ( .A(adder_a[13]), .B(
        adder_b[13]), .CI(\struct_adder/add_1_root_add_19_2/carry[13] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[14] ), .S(adder_out[13]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_12  ( .A(adder_a[12]), .B(
        adder_b[12]), .CI(\struct_adder/add_1_root_add_19_2/carry[12] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[13] ), .S(adder_out[12]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_11  ( .A(adder_a[11]), .B(
        adder_b[11]), .CI(\struct_adder/add_1_root_add_19_2/carry[11] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[12] ), .S(adder_out[11]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_10  ( .A(adder_a[10]), .B(
        adder_b[10]), .CI(\struct_adder/add_1_root_add_19_2/carry[10] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[11] ), .S(adder_out[10]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_9  ( .A(adder_a[9]), .B(
        adder_b[9]), .CI(\struct_adder/add_1_root_add_19_2/carry[9] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[10] ), .S(adder_out[9]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_8  ( .A(adder_a[8]), .B(
        adder_b[8]), .CI(\struct_adder/add_1_root_add_19_2/carry[8] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[9] ), .S(adder_out[8]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_7  ( .A(adder_a[7]), .B(
        adder_b[7]), .CI(\struct_adder/add_1_root_add_19_2/carry[7] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[8] ), .S(adder_out[7]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_6  ( .A(adder_a[6]), .B(
        adder_b[6]), .CI(\struct_adder/add_1_root_add_19_2/carry[6] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[7] ), .S(adder_out[6]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_5  ( .A(adder_a[5]), .B(
        adder_b[5]), .CI(\struct_adder/add_1_root_add_19_2/carry[5] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[6] ), .S(adder_out[5]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_4  ( .A(adder_a[4]), .B(
        adder_b[4]), .CI(\struct_adder/add_1_root_add_19_2/carry[4] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[5] ), .S(adder_out[4]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_3  ( .A(adder_a[3]), .B(
        adder_b[3]), .CI(\struct_adder/add_1_root_add_19_2/carry[3] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[4] ), .S(adder_out[3]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_2  ( .A(adder_a[2]), .B(
        adder_b[2]), .CI(\struct_adder/add_1_root_add_19_2/carry[2] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[3] ), .S(adder_out[2]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_1  ( .A(adder_a[1]), .B(
        adder_b[1]), .CI(\struct_adder/add_1_root_add_19_2/carry[1] ), .CO(
        \struct_adder/add_1_root_add_19_2/carry[2] ), .S(adder_out[1]) );
  SEN_ADDF_0P5 \struct_adder/add_1_root_add_19_2/U1_0  ( .A(adder_a[0]), .B(
        adder_b[0]), .CI(adder_cin), .CO(
        \struct_adder/add_1_root_add_19_2/carry[1] ), .S(adder_out[0]) );
  SEN_AOI22_0P5 U316 ( .A1(n251), .A2(adder_out[27]), .B1(n247), .B2(n262), 
        .X(n123) );
  SEN_EN3_0P5 U317 ( .A1(adder_a[31]), .A2(adder_b[31]), .A3(
        \struct_adder/add_1_root_add_19_2/carry[31] ), .X(n218) );
  SEN_INV_S_0P5 U318 ( .A(n218), .X(adder_out[31]) );
  SEN_AOI22_0P5 U319 ( .A1(n251), .A2(adder_out[28]), .B1(n247), .B2(n261), 
        .X(n120) );
  SEN_MAJ3_0P5 U320 ( .A1(adder_out[31]), .A2(adder_a[31]), .A3(adder_b[31]), 
        .X(n185) );
  SEN_AOI22_0P5 U321 ( .A1(n251), .A2(adder_out[29]), .B1(n247), .B2(n260), 
        .X(n117) );
  SEN_AOI31_0P5 U322 ( .A1(INST[2]), .A2(INST[1]), .A3(INST[0]), .B(n323), .X(
        n217) );
  SEN_AOI22_0P5 U323 ( .A1(n251), .A2(adder_out[30]), .B1(n84), .B2(n259), .X(
        n111) );
  SEN_NR4_0P5 U324 ( .A1(adder_out[23]), .A2(adder_out[22]), .A3(adder_out[21]), .A4(adder_out[20]), .X(n219) );
  SEN_INV_S_0P5 U325 ( .A(n219), .X(n209) );
  SEN_AOI22_0P5 U326 ( .A1(n251), .A2(adder_out[31]), .B1(n84), .B2(n258), .X(
        n108) );
  SEN_MUXI2_S_0P5 U327 ( .D0(n223), .D1(n216), .S(B[0]), .X(N156) );
  SEN_INV_S_0P5 U328 ( .A(N188), .X(n257) );
  SEN_ND2_S_0P5 U329 ( .A1(n216), .A2(n223), .X(n220) );
  SEN_INV_S_0P5 U330 ( .A(n85), .X(n246) );
  SEN_INV_S_0P5 U331 ( .A(n241), .X(n239) );
  SEN_INV_S_0P5 U332 ( .A(n241), .X(n240) );
  SEN_INV_S_0P5 U333 ( .A(n87), .X(n238) );
  SEN_INV_S_0P5 U334 ( .A(n83), .X(n252) );
  SEN_INV_S_0P5 U335 ( .A(n84), .X(n249) );
  SEN_INV_S_0P5 U336 ( .A(n216), .X(n229) );
  SEN_INV_S_0P5 U337 ( .A(n214), .X(n235) );
  SEN_INV_S_0P5 U338 ( .A(n86), .X(n241) );
  SEN_INV_S_0P5 U339 ( .A(n257), .X(n256) );
  SEN_INV_S_0P5 U340 ( .A(n257), .X(n255) );
  SEN_INV_S_0P5 U341 ( .A(n257), .X(n254) );
  SEN_INV_S_0P5 U342 ( .A(n257), .X(n253) );
  SEN_INV_S_0P5 U343 ( .A(n220), .X(n230) );
  SEN_INV_S_0P5 U344 ( .A(n220), .X(n231) );
  SEN_INV_S_0P5 U345 ( .A(n220), .X(n232) );
  SEN_INV_S_0P5 U346 ( .A(n246), .X(n242) );
  SEN_INV_S_0P5 U347 ( .A(n246), .X(n243) );
  SEN_INV_S_0P5 U348 ( .A(n178), .X(n322) );
  SEN_INV_S_0P5 U349 ( .A(n246), .X(n244) );
  SEN_INV_S_0P5 U350 ( .A(n179), .X(n224) );
  SEN_INV_S_0P5 U351 ( .A(n179), .X(n225) );
  SEN_INV_S_0P5 U352 ( .A(n246), .X(n245) );
  SEN_INV_S_0P5 U353 ( .A(n179), .X(n226) );
  SEN_ND2_S_0P5 U354 ( .A1(n232), .A2(n234), .X(N188) );
  SEN_ND2_S_0P5 U355 ( .A1(n223), .A2(n234), .X(N189) );
  SEN_ND2_S_0P5 U356 ( .A1(n189), .A2(n200), .X(n178) );
  SEN_INV_S_0P5 U357 ( .A(n252), .X(n250) );
  SEN_INV_S_0P5 U358 ( .A(n252), .X(n251) );
  SEN_INV_S_0P5 U359 ( .A(n249), .X(n248) );
  SEN_INV_S_0P5 U360 ( .A(n249), .X(n247) );
  SEN_INV_S_0P5 U361 ( .A(n238), .X(n236) );
  SEN_INV_S_0P5 U362 ( .A(n238), .X(n237) );
  SEN_INV_S_0P5 U363 ( .A(n235), .X(n233) );
  SEN_INV_S_0P5 U364 ( .A(n217), .X(n222) );
  SEN_INV_S_0P5 U365 ( .A(n217), .X(n221) );
  SEN_INV_S_0P5 U366 ( .A(n229), .X(n228) );
  SEN_INV_S_0P5 U367 ( .A(n229), .X(n227) );
  SEN_INV_S_0P5 U368 ( .A(n203), .X(n330) );
  SEN_INV_S_0P5 U369 ( .A(n235), .X(n234) );
  SEN_INV_S_0P5 U370 ( .A(n217), .X(n223) );
  SEN_NR2B_V1_1 U371 ( .A(n199), .B(n191), .X(n85) );
  SEN_NR2B_V1_1 U372 ( .A(n188), .B(n189), .X(n83) );
  SEN_NR2_S_0P5 U373 ( .A1(n323), .A2(n327), .X(n189) );
  SEN_OAI221_0P5 U374 ( .A1(n184), .A2(n185), .B1(n186), .B2(n329), .C(n187), 
        .X(n183) );
  SEN_AOI22_0P5 U375 ( .A1(n290), .A2(n84), .B1(n250), .B2(adder_out[0]), .X(
        n187) );
  SEN_NR2_S_0P5 U376 ( .A1(n325), .A2(n326), .X(n200) );
  SEN_AO2BB2_0P5 U377 ( .A1(n191), .A2(n323), .B1(n198), .B2(n202), .X(n204)
         );
  SEN_INV_S_0P5 U378 ( .A(A[0]), .X(n290) );
  SEN_NR2B_V1_1 U379 ( .A(n190), .B(n191), .X(n84) );
  SEN_OAI22_S_0P5 U380 ( .A1(n329), .A2(n326), .B1(n325), .B2(n185), .X(n201)
         );
  SEN_OAI211_0P5 U381 ( .A1(n145), .A2(n321), .B1(n146), .B2(n147), .X(Z[1])
         );
  SEN_AOI22_0P5 U382 ( .A1(adder_out[1]), .A2(n250), .B1(n248), .B2(n288), .X(
        n147) );
  SEN_AOAI211_0P5 U383 ( .A1(n243), .A2(n321), .B(n239), .C(A[1]), .X(n146) );
  SEN_AOI221_0P5 U384 ( .A1(n244), .A2(n288), .B1(A[1]), .B2(n224), .C(n236), 
        .X(n145) );
  SEN_OAI211_0P5 U385 ( .A1(n112), .A2(n320), .B1(n113), .B2(n114), .X(Z[2])
         );
  SEN_AOI22_0P5 U386 ( .A1(adder_out[2]), .A2(n251), .B1(n247), .B2(n287), .X(
        n114) );
  SEN_AOAI211_0P5 U387 ( .A1(n242), .A2(n320), .B(n240), .C(A[2]), .X(n113) );
  SEN_AOI221_0P5 U388 ( .A1(n243), .A2(n287), .B1(A[2]), .B2(n225), .C(n237), 
        .X(n112) );
  SEN_OAI211_0P5 U389 ( .A1(n103), .A2(n319), .B1(n104), .B2(n105), .X(Z[3])
         );
  SEN_AOI22_0P5 U390 ( .A1(adder_out[3]), .A2(n251), .B1(n247), .B2(n286), .X(
        n105) );
  SEN_AOAI211_0P5 U391 ( .A1(n242), .A2(n319), .B(n240), .C(A[3]), .X(n104) );
  SEN_AOI221_0P5 U392 ( .A1(n245), .A2(n286), .B1(A[3]), .B2(n225), .C(n237), 
        .X(n103) );
  SEN_OAI211_0P5 U393 ( .A1(n100), .A2(n318), .B1(n101), .B2(n102), .X(Z[4])
         );
  SEN_AOI22_0P5 U394 ( .A1(adder_out[4]), .A2(n251), .B1(n247), .B2(n285), .X(
        n102) );
  SEN_AOAI211_0P5 U395 ( .A1(n242), .A2(n318), .B(n240), .C(A[4]), .X(n101) );
  SEN_AOI221_0P5 U396 ( .A1(n245), .A2(n285), .B1(A[4]), .B2(n225), .C(n237), 
        .X(n100) );
  SEN_OAI211_0P5 U397 ( .A1(n97), .A2(n317), .B1(n98), .B2(n99), .X(Z[5]) );
  SEN_AOI22_0P5 U398 ( .A1(adder_out[5]), .A2(n251), .B1(n247), .B2(n284), .X(
        n99) );
  SEN_AOAI211_0P5 U399 ( .A1(n242), .A2(n317), .B(n240), .C(A[5]), .X(n98) );
  SEN_AOI221_0P5 U400 ( .A1(n243), .A2(n284), .B1(A[5]), .B2(n225), .C(n237), 
        .X(n97) );
  SEN_OAI211_0P5 U401 ( .A1(n94), .A2(n316), .B1(n95), .B2(n96), .X(Z[6]) );
  SEN_AOI22_0P5 U402 ( .A1(adder_out[6]), .A2(n251), .B1(n247), .B2(n283), .X(
        n96) );
  SEN_AOAI211_0P5 U403 ( .A1(n242), .A2(n316), .B(n240), .C(A[6]), .X(n95) );
  SEN_AOI221_0P5 U404 ( .A1(n242), .A2(n283), .B1(A[6]), .B2(n225), .C(n237), 
        .X(n94) );
  SEN_OAI211_0P5 U405 ( .A1(n91), .A2(n315), .B1(n92), .B2(n93), .X(Z[7]) );
  SEN_AOI22_0P5 U406 ( .A1(adder_out[7]), .A2(n250), .B1(n247), .B2(n282), .X(
        n93) );
  SEN_AOAI211_0P5 U407 ( .A1(n242), .A2(n315), .B(n239), .C(A[7]), .X(n92) );
  SEN_AOI221_0P5 U408 ( .A1(n242), .A2(n282), .B1(A[7]), .B2(n226), .C(n236), 
        .X(n91) );
  SEN_OAI211_0P5 U409 ( .A1(n88), .A2(n314), .B1(n89), .B2(n90), .X(Z[8]) );
  SEN_AOI22_0P5 U410 ( .A1(adder_out[8]), .A2(n83), .B1(n247), .B2(n281), .X(
        n90) );
  SEN_AOAI211_0P5 U411 ( .A1(n242), .A2(n314), .B(n86), .C(A[8]), .X(n89) );
  SEN_AOI221_0P5 U412 ( .A1(n85), .A2(n281), .B1(A[8]), .B2(n226), .C(n237), 
        .X(n88) );
  SEN_OAI211_0P5 U413 ( .A1(n80), .A2(n313), .B1(n81), .B2(n82), .X(Z[9]) );
  SEN_AOI22_0P5 U414 ( .A1(adder_out[9]), .A2(n83), .B1(n247), .B2(n280), .X(
        n82) );
  SEN_AOAI211_0P5 U415 ( .A1(n243), .A2(n313), .B(n86), .C(A[9]), .X(n81) );
  SEN_AOI221_0P5 U416 ( .A1(n85), .A2(n280), .B1(n226), .B2(A[9]), .C(n87), 
        .X(n80) );
  SEN_OAI211_0P5 U417 ( .A1(n175), .A2(n312), .B1(n176), .B2(n177), .X(Z[10])
         );
  SEN_AOI22_0P5 U418 ( .A1(adder_out[10]), .A2(n250), .B1(n84), .B2(n279), .X(
        n177) );
  SEN_AOAI211_0P5 U419 ( .A1(n244), .A2(n312), .B(n239), .C(A[10]), .X(n176)
         );
  SEN_AOI221_0P5 U420 ( .A1(n85), .A2(n279), .B1(A[10]), .B2(n224), .C(n236), 
        .X(n175) );
  SEN_OAI211_0P5 U421 ( .A1(n172), .A2(n311), .B1(n173), .B2(n174), .X(Z[11])
         );
  SEN_AOI22_0P5 U422 ( .A1(adder_out[11]), .A2(n250), .B1(n84), .B2(n278), .X(
        n174) );
  SEN_AOAI211_0P5 U423 ( .A1(n244), .A2(n311), .B(n239), .C(A[11]), .X(n173)
         );
  SEN_AOI221_0P5 U424 ( .A1(n85), .A2(n278), .B1(A[11]), .B2(n224), .C(n236), 
        .X(n172) );
  SEN_OAI211_0P5 U425 ( .A1(n169), .A2(n310), .B1(n170), .B2(n171), .X(Z[12])
         );
  SEN_AOI22_0P5 U426 ( .A1(adder_out[12]), .A2(n250), .B1(n84), .B2(n277), .X(
        n171) );
  SEN_AOAI211_0P5 U427 ( .A1(n243), .A2(n310), .B(n239), .C(A[12]), .X(n170)
         );
  SEN_AOI221_0P5 U428 ( .A1(n245), .A2(n277), .B1(A[12]), .B2(n224), .C(n236), 
        .X(n169) );
  SEN_OAI211_0P5 U429 ( .A1(n166), .A2(n309), .B1(n167), .B2(n168), .X(Z[13])
         );
  SEN_AOI22_0P5 U430 ( .A1(adder_out[13]), .A2(n250), .B1(n84), .B2(n276), .X(
        n168) );
  SEN_AOAI211_0P5 U431 ( .A1(n244), .A2(n309), .B(n239), .C(A[13]), .X(n167)
         );
  SEN_AOI221_0P5 U432 ( .A1(n245), .A2(n276), .B1(A[13]), .B2(n224), .C(n236), 
        .X(n166) );
  SEN_OAI211_0P5 U433 ( .A1(n163), .A2(n308), .B1(n164), .B2(n165), .X(Z[14])
         );
  SEN_AOI22_0P5 U434 ( .A1(adder_out[14]), .A2(n250), .B1(n84), .B2(n275), .X(
        n165) );
  SEN_AOAI211_0P5 U435 ( .A1(n244), .A2(n308), .B(n239), .C(A[14]), .X(n164)
         );
  SEN_AOI221_0P5 U436 ( .A1(n245), .A2(n275), .B1(A[14]), .B2(n224), .C(n236), 
        .X(n163) );
  SEN_OAI211_0P5 U437 ( .A1(n160), .A2(n307), .B1(n161), .B2(n162), .X(Z[15])
         );
  SEN_AOI22_0P5 U438 ( .A1(adder_out[15]), .A2(n250), .B1(n248), .B2(n274), 
        .X(n162) );
  SEN_AOAI211_0P5 U439 ( .A1(n243), .A2(n307), .B(n239), .C(A[15]), .X(n161)
         );
  SEN_AOI221_0P5 U440 ( .A1(n245), .A2(n274), .B1(A[15]), .B2(n224), .C(n236), 
        .X(n160) );
  SEN_OAI211_0P5 U441 ( .A1(n157), .A2(n306), .B1(n158), .B2(n159), .X(Z[16])
         );
  SEN_AOI22_0P5 U442 ( .A1(adder_out[16]), .A2(n250), .B1(n248), .B2(n273), 
        .X(n159) );
  SEN_AOAI211_0P5 U443 ( .A1(n244), .A2(n306), .B(n239), .C(A[16]), .X(n158)
         );
  SEN_AOI221_0P5 U444 ( .A1(n245), .A2(n273), .B1(A[16]), .B2(n224), .C(n236), 
        .X(n157) );
  SEN_OAI211_0P5 U445 ( .A1(n154), .A2(n305), .B1(n155), .B2(n156), .X(Z[17])
         );
  SEN_AOI22_0P5 U446 ( .A1(adder_out[17]), .A2(n250), .B1(n248), .B2(n272), 
        .X(n156) );
  SEN_AOAI211_0P5 U447 ( .A1(n244), .A2(n305), .B(n239), .C(A[17]), .X(n155)
         );
  SEN_AOI221_0P5 U448 ( .A1(n245), .A2(n272), .B1(A[17]), .B2(n224), .C(n236), 
        .X(n154) );
  SEN_OAI211_0P5 U449 ( .A1(n151), .A2(n304), .B1(n152), .B2(n153), .X(Z[18])
         );
  SEN_AOI22_0P5 U450 ( .A1(adder_out[18]), .A2(n250), .B1(n248), .B2(n271), 
        .X(n153) );
  SEN_AOAI211_0P5 U451 ( .A1(n243), .A2(n304), .B(n239), .C(A[18]), .X(n152)
         );
  SEN_AOI221_0P5 U452 ( .A1(n244), .A2(n271), .B1(A[18]), .B2(n224), .C(n236), 
        .X(n151) );
  SEN_OAI211_0P5 U453 ( .A1(n148), .A2(n303), .B1(n149), .B2(n150), .X(Z[19])
         );
  SEN_AOI22_0P5 U454 ( .A1(adder_out[19]), .A2(n250), .B1(n248), .B2(n270), 
        .X(n150) );
  SEN_AOAI211_0P5 U455 ( .A1(n243), .A2(n303), .B(n239), .C(A[19]), .X(n149)
         );
  SEN_AOI221_0P5 U456 ( .A1(n245), .A2(n270), .B1(A[19]), .B2(n224), .C(n236), 
        .X(n148) );
  SEN_OAI211_0P5 U457 ( .A1(n142), .A2(n302), .B1(n143), .B2(n144), .X(Z[20])
         );
  SEN_AOI22_0P5 U458 ( .A1(adder_out[20]), .A2(n250), .B1(n248), .B2(n269), 
        .X(n144) );
  SEN_AOAI211_0P5 U459 ( .A1(n243), .A2(n302), .B(n239), .C(A[20]), .X(n143)
         );
  SEN_AOI221_0P5 U460 ( .A1(n244), .A2(n269), .B1(A[20]), .B2(n224), .C(n236), 
        .X(n142) );
  SEN_OAI211_0P5 U461 ( .A1(n139), .A2(n301), .B1(n140), .B2(n141), .X(Z[21])
         );
  SEN_AOI22_0P5 U462 ( .A1(adder_out[21]), .A2(n250), .B1(n248), .B2(n268), 
        .X(n141) );
  SEN_AOAI211_0P5 U463 ( .A1(n243), .A2(n301), .B(n239), .C(A[21]), .X(n140)
         );
  SEN_AOI221_0P5 U464 ( .A1(n244), .A2(n268), .B1(A[21]), .B2(n224), .C(n236), 
        .X(n139) );
  SEN_OAI211_0P5 U465 ( .A1(n136), .A2(n300), .B1(n137), .B2(n138), .X(Z[22])
         );
  SEN_AOI22_0P5 U466 ( .A1(adder_out[22]), .A2(n251), .B1(n248), .B2(n267), 
        .X(n138) );
  SEN_AOAI211_0P5 U467 ( .A1(n243), .A2(n300), .B(n240), .C(A[22]), .X(n137)
         );
  SEN_AOI221_0P5 U468 ( .A1(n244), .A2(n267), .B1(A[22]), .B2(n224), .C(n236), 
        .X(n136) );
  SEN_OAI211_0P5 U469 ( .A1(n133), .A2(n299), .B1(n134), .B2(n135), .X(Z[23])
         );
  SEN_AOI22_0P5 U470 ( .A1(adder_out[23]), .A2(n251), .B1(n248), .B2(n266), 
        .X(n135) );
  SEN_AOAI211_0P5 U471 ( .A1(n243), .A2(n299), .B(n240), .C(A[23]), .X(n134)
         );
  SEN_AOI221_0P5 U472 ( .A1(n244), .A2(n266), .B1(A[23]), .B2(n225), .C(n237), 
        .X(n133) );
  SEN_OAI211_0P5 U473 ( .A1(n130), .A2(n298), .B1(n131), .B2(n132), .X(Z[24])
         );
  SEN_AOI22_0P5 U474 ( .A1(adder_out[24]), .A2(n251), .B1(n248), .B2(n265), 
        .X(n132) );
  SEN_AOAI211_0P5 U475 ( .A1(n243), .A2(n298), .B(n240), .C(A[24]), .X(n131)
         );
  SEN_AOI221_0P5 U476 ( .A1(n244), .A2(n265), .B1(A[24]), .B2(n225), .C(n237), 
        .X(n130) );
  SEN_OAI211_0P5 U477 ( .A1(n127), .A2(n297), .B1(n128), .B2(n129), .X(Z[25])
         );
  SEN_AOI22_0P5 U478 ( .A1(adder_out[25]), .A2(n251), .B1(n248), .B2(n264), 
        .X(n129) );
  SEN_AOAI211_0P5 U479 ( .A1(n243), .A2(n297), .B(n240), .C(A[25]), .X(n128)
         );
  SEN_AOI221_0P5 U480 ( .A1(n244), .A2(n264), .B1(A[25]), .B2(n225), .C(n237), 
        .X(n127) );
  SEN_OAI211_0P5 U481 ( .A1(n124), .A2(n296), .B1(n125), .B2(n126), .X(Z[26])
         );
  SEN_AOI22_0P5 U482 ( .A1(adder_out[26]), .A2(n251), .B1(n248), .B2(n263), 
        .X(n126) );
  SEN_AOAI211_0P5 U483 ( .A1(n243), .A2(n296), .B(n240), .C(A[26]), .X(n125)
         );
  SEN_AOI221_0P5 U484 ( .A1(n245), .A2(n263), .B1(A[26]), .B2(n225), .C(n237), 
        .X(n124) );
  SEN_OAI211_0P5 U485 ( .A1(n121), .A2(n295), .B1(n122), .B2(n123), .X(Z[27])
         );
  SEN_AOAI211_0P5 U486 ( .A1(n242), .A2(n295), .B(n240), .C(A[27]), .X(n122)
         );
  SEN_AOI221_0P5 U487 ( .A1(n245), .A2(n262), .B1(A[27]), .B2(n225), .C(n237), 
        .X(n121) );
  SEN_OAI211_0P5 U488 ( .A1(n118), .A2(n294), .B1(n119), .B2(n120), .X(Z[28])
         );
  SEN_AOAI211_0P5 U489 ( .A1(n242), .A2(n294), .B(n240), .C(A[28]), .X(n119)
         );
  SEN_AOI221_0P5 U490 ( .A1(n245), .A2(n261), .B1(A[28]), .B2(n225), .C(n237), 
        .X(n118) );
  SEN_OAI211_0P5 U491 ( .A1(n115), .A2(n293), .B1(n116), .B2(n117), .X(Z[29])
         );
  SEN_AOAI211_0P5 U492 ( .A1(n242), .A2(n293), .B(n240), .C(A[29]), .X(n116)
         );
  SEN_AOI221_0P5 U493 ( .A1(n245), .A2(n260), .B1(A[29]), .B2(n225), .C(n237), 
        .X(n115) );
  SEN_OAI211_0P5 U494 ( .A1(n109), .A2(n292), .B1(n110), .B2(n111), .X(Z[30])
         );
  SEN_AOAI211_0P5 U495 ( .A1(n242), .A2(n292), .B(n240), .C(A[30]), .X(n110)
         );
  SEN_AOI221_0P5 U496 ( .A1(n245), .A2(n259), .B1(A[30]), .B2(n225), .C(n237), 
        .X(n109) );
  SEN_OAI211_0P5 U497 ( .A1(n106), .A2(n291), .B1(n107), .B2(n108), .X(Z[31])
         );
  SEN_AOAI211_0P5 U498 ( .A1(n242), .A2(n291), .B(n240), .C(A[31]), .X(n107)
         );
  SEN_AOI221_0P5 U499 ( .A1(n245), .A2(n258), .B1(A[31]), .B2(n225), .C(n237), 
        .X(n106) );
  SEN_ND2_S_0P5 U500 ( .A1(n189), .A2(n198), .X(n184) );
  SEN_INV_S_0P5 U501 ( .A(A[1]), .X(n288) );
  SEN_INV_S_0P5 U502 ( .A(A[2]), .X(n287) );
  SEN_INV_S_0P5 U503 ( .A(A[3]), .X(n286) );
  SEN_INV_S_0P5 U504 ( .A(A[4]), .X(n285) );
  SEN_INV_S_0P5 U505 ( .A(A[5]), .X(n284) );
  SEN_INV_S_0P5 U506 ( .A(A[6]), .X(n283) );
  SEN_INV_S_0P5 U507 ( .A(A[7]), .X(n282) );
  SEN_INV_S_0P5 U508 ( .A(A[8]), .X(n281) );
  SEN_INV_S_0P5 U509 ( .A(A[9]), .X(n280) );
  SEN_INV_S_0P5 U510 ( .A(A[10]), .X(n279) );
  SEN_INV_S_0P5 U511 ( .A(A[11]), .X(n278) );
  SEN_INV_S_0P5 U512 ( .A(A[12]), .X(n277) );
  SEN_INV_S_0P5 U513 ( .A(A[13]), .X(n276) );
  SEN_INV_S_0P5 U514 ( .A(A[14]), .X(n275) );
  SEN_INV_S_0P5 U515 ( .A(A[15]), .X(n274) );
  SEN_INV_S_0P5 U516 ( .A(A[16]), .X(n273) );
  SEN_INV_S_0P5 U517 ( .A(A[17]), .X(n272) );
  SEN_INV_S_0P5 U518 ( .A(A[18]), .X(n271) );
  SEN_INV_S_0P5 U519 ( .A(A[19]), .X(n270) );
  SEN_INV_S_0P5 U520 ( .A(A[20]), .X(n269) );
  SEN_INV_S_0P5 U521 ( .A(A[21]), .X(n268) );
  SEN_INV_S_0P5 U522 ( .A(A[22]), .X(n267) );
  SEN_INV_S_0P5 U523 ( .A(A[23]), .X(n266) );
  SEN_INV_S_0P5 U524 ( .A(A[24]), .X(n265) );
  SEN_INV_S_0P5 U525 ( .A(A[25]), .X(n264) );
  SEN_INV_S_0P5 U526 ( .A(A[26]), .X(n263) );
  SEN_INV_S_0P5 U527 ( .A(A[27]), .X(n262) );
  SEN_INV_S_0P5 U528 ( .A(A[28]), .X(n261) );
  SEN_INV_S_0P5 U529 ( .A(A[29]), .X(n260) );
  SEN_INV_S_0P5 U530 ( .A(A[30]), .X(n259) );
  SEN_INV_S_0P5 U531 ( .A(A[31]), .X(n258) );
  SEN_ND2_S_0P5 U532 ( .A1(n199), .A2(n200), .X(n194) );
  SEN_ND2_S_0P5 U533 ( .A1(n188), .A2(n189), .X(n186) );
  SEN_ND2_S_0P5 U534 ( .A1(n199), .A2(n198), .X(n179) );
  SEN_ND2_S_0P5 U535 ( .A1(n190), .A2(n198), .X(n195) );
  SEN_ND2_S_0P5 U536 ( .A1(n200), .A2(n190), .X(n193) );
  SEN_ND2_S_0P5 U537 ( .A1(n324), .A2(n178), .X(n87) );
  SEN_NR4_0P5 U538 ( .A1(adder_out[24]), .A2(adder_out[25]), .A3(adder_out[26]), .A4(adder_out[27]), .X(n213) );
  SEN_NR4_0P5 U539 ( .A1(adder_out[28]), .A2(adder_out[29]), .A3(adder_out[2]), 
        .A4(adder_out[30]), .X(n212) );
  SEN_NR4_0P5 U540 ( .A1(adder_out[31]), .A2(adder_out[3]), .A3(adder_out[4]), 
        .A4(adder_out[5]), .X(n211) );
  SEN_NR4_0P5 U541 ( .A1(adder_out[6]), .A2(adder_out[7]), .A3(adder_out[8]), 
        .A4(adder_out[9]), .X(n210) );
  SEN_NR4_0P5 U542 ( .A1(adder_out[16]), .A2(adder_out[15]), .A3(adder_out[14]), .A4(adder_out[13]), .X(n206) );
  SEN_AN4B_0P5 U543 ( .B1(n205), .B2(n206), .B3(n207), .A(n208), .X(n203) );
  SEN_AN4_0P5 U544 ( .A1(n210), .A2(n211), .A3(n212), .A4(n213), .X(n207) );
  SEN_OR5_1 U545 ( .A1(adder_out[17]), .A2(adder_out[18]), .A3(adder_out[19]), 
        .A4(adder_out[1]), .A5(n209), .X(n208) );
  SEN_NR4_0P5 U546 ( .A1(adder_out[12]), .A2(adder_out[11]), .A3(adder_out[10]), .A4(adder_out[0]), .X(n205) );
  SEN_INV_S_0P5 U547 ( .A(n185), .X(n329) );
  SEN_ND2_S_0P5 U548 ( .A1(n188), .A2(n199), .X(n216) );
  SEN_ND2_S_0P5 U549 ( .A1(n188), .A2(n190), .X(n214) );
  SEN_OAI22_S_0P5 U550 ( .A1(n230), .A2(n290), .B1(A[0]), .B2(n233), .X(N124)
         );
  SEN_OAI22_S_0P5 U551 ( .A1(n230), .A2(n288), .B1(A[1]), .B2(n233), .X(N125)
         );
  SEN_OAI22_S_0P5 U552 ( .A1(n230), .A2(n287), .B1(A[2]), .B2(n233), .X(N126)
         );
  SEN_OAI22_S_0P5 U553 ( .A1(n230), .A2(n286), .B1(A[3]), .B2(n233), .X(N127)
         );
  SEN_OAI22_S_0P5 U554 ( .A1(n230), .A2(n285), .B1(A[4]), .B2(n233), .X(N128)
         );
  SEN_OAI22_S_0P5 U555 ( .A1(n230), .A2(n284), .B1(A[5]), .B2(n233), .X(N129)
         );
  SEN_OAI22_S_0P5 U556 ( .A1(n230), .A2(n283), .B1(A[6]), .B2(n233), .X(N130)
         );
  SEN_OAI22_S_0P5 U557 ( .A1(n230), .A2(n282), .B1(A[7]), .B2(n233), .X(N131)
         );
  SEN_OAI22_S_0P5 U558 ( .A1(n230), .A2(n281), .B1(A[8]), .B2(n233), .X(N132)
         );
  SEN_OAI22_S_0P5 U559 ( .A1(n230), .A2(n280), .B1(A[9]), .B2(n233), .X(N133)
         );
  SEN_OAI22_S_0P5 U560 ( .A1(n230), .A2(n279), .B1(A[10]), .B2(n233), .X(N134)
         );
  SEN_OAI22_S_0P5 U561 ( .A1(n230), .A2(n278), .B1(A[11]), .B2(n233), .X(N135)
         );
  SEN_OAI22_S_0P5 U562 ( .A1(n230), .A2(n277), .B1(A[12]), .B2(n233), .X(N136)
         );
  SEN_OAI22_S_0P5 U563 ( .A1(n231), .A2(n276), .B1(A[13]), .B2(n214), .X(N137)
         );
  SEN_OAI22_S_0P5 U564 ( .A1(n231), .A2(n275), .B1(A[14]), .B2(n214), .X(N138)
         );
  SEN_OAI22_S_0P5 U565 ( .A1(n231), .A2(n274), .B1(A[15]), .B2(n214), .X(N139)
         );
  SEN_OAI22_S_0P5 U566 ( .A1(n231), .A2(n273), .B1(A[16]), .B2(n214), .X(N140)
         );
  SEN_OAI22_S_0P5 U567 ( .A1(n231), .A2(n272), .B1(A[17]), .B2(n214), .X(N141)
         );
  SEN_OAI22_S_0P5 U568 ( .A1(n231), .A2(n271), .B1(A[18]), .B2(n214), .X(N142)
         );
  SEN_OAI22_S_0P5 U569 ( .A1(n231), .A2(n270), .B1(A[19]), .B2(n214), .X(N143)
         );
  SEN_OAI22_S_0P5 U570 ( .A1(n231), .A2(n269), .B1(A[20]), .B2(n234), .X(N144)
         );
  SEN_OAI22_S_0P5 U571 ( .A1(n231), .A2(n268), .B1(A[21]), .B2(n214), .X(N145)
         );
  SEN_OAI22_S_0P5 U572 ( .A1(n231), .A2(n267), .B1(A[22]), .B2(n234), .X(N146)
         );
  SEN_OAI22_S_0P5 U573 ( .A1(n231), .A2(n266), .B1(A[23]), .B2(n214), .X(N147)
         );
  SEN_OAI22_S_0P5 U574 ( .A1(n231), .A2(n265), .B1(A[24]), .B2(n234), .X(N148)
         );
  SEN_OAI22_S_0P5 U575 ( .A1(n231), .A2(n264), .B1(A[25]), .B2(n214), .X(N149)
         );
  SEN_OAI22_S_0P5 U576 ( .A1(n232), .A2(n263), .B1(A[26]), .B2(n234), .X(N150)
         );
  SEN_OAI22_S_0P5 U577 ( .A1(n232), .A2(n262), .B1(A[27]), .B2(n234), .X(N151)
         );
  SEN_OAI22_S_0P5 U578 ( .A1(n232), .A2(n261), .B1(A[28]), .B2(n234), .X(N152)
         );
  SEN_OAI22_S_0P5 U579 ( .A1(n232), .A2(n260), .B1(A[29]), .B2(n234), .X(N153)
         );
  SEN_OAI22_S_0P5 U580 ( .A1(n232), .A2(n259), .B1(A[30]), .B2(n234), .X(N154)
         );
  SEN_OAI22_S_0P5 U581 ( .A1(n232), .A2(n258), .B1(A[31]), .B2(n234), .X(N155)
         );
  SEN_ND2_S_0P5 U582 ( .A1(INST[2]), .A2(n326), .X(n191) );
  SEN_NR2_S_0P5 U583 ( .A1(INST[2]), .A2(INST[1]), .X(n188) );
  SEN_INV_S_0P5 U584 ( .A(SEL), .X(n328) );
  SEN_NR2_S_0P5 U585 ( .A1(INST[3]), .A2(INST[0]), .X(n199) );
  SEN_NR2_S_0P5 U586 ( .A1(n326), .A2(INST[2]), .X(n198) );
  SEN_AOI22_0P5 U587 ( .A1(B[0]), .A2(n192), .B1(A[0]), .B2(n239), .X(n182) );
  SEN_OAI211_0P5 U588 ( .A1(n179), .A2(n290), .B1(n324), .B2(n196), .X(n192)
         );
  SEN_AOI22_0P5 U589 ( .A1(n322), .A2(n328), .B1(n244), .B2(n290), .X(n196) );
  SEN_NR2_S_0P5 U590 ( .A1(n327), .A2(INST[3]), .X(n190) );
  SEN_INV_S_0P5 U591 ( .A(INST[1]), .X(n326) );
  SEN_INV_S_0P5 U592 ( .A(INST[2]), .X(n325) );
  SEN_OAI2111_0P5 U593 ( .A1(B[0]), .A2(n180), .B1(n181), .B2(n182), .B3(n289), 
        .X(Z[0]) );
  SEN_AOI32_1 U594 ( .A1(n201), .A2(n330), .A3(n202), .B1(n203), .B2(n204), 
        .X(n181) );
  SEN_AOI22_0P5 U595 ( .A1(n322), .A2(SEL), .B1(A[0]), .B2(n242), .X(n180) );
  SEN_INV_S_0P5 U596 ( .A(n183), .X(n289) );
  SEN_OAI221_0P5 U597 ( .A1(n193), .A2(n328), .B1(SEL), .B2(n194), .C(n195), 
        .X(n86) );
  SEN_INV_S_0P5 U598 ( .A(B[1]), .X(n321) );
  SEN_INV_S_0P5 U599 ( .A(B[2]), .X(n320) );
  SEN_INV_S_0P5 U600 ( .A(B[3]), .X(n319) );
  SEN_INV_S_0P5 U601 ( .A(B[4]), .X(n318) );
  SEN_INV_S_0P5 U602 ( .A(B[5]), .X(n317) );
  SEN_INV_S_0P5 U603 ( .A(B[6]), .X(n316) );
  SEN_INV_S_0P5 U604 ( .A(B[7]), .X(n315) );
  SEN_INV_S_0P5 U605 ( .A(B[8]), .X(n314) );
  SEN_INV_S_0P5 U606 ( .A(B[9]), .X(n313) );
  SEN_INV_S_0P5 U607 ( .A(B[10]), .X(n312) );
  SEN_INV_S_0P5 U608 ( .A(B[11]), .X(n311) );
  SEN_INV_S_0P5 U609 ( .A(B[12]), .X(n310) );
  SEN_INV_S_0P5 U610 ( .A(B[13]), .X(n309) );
  SEN_INV_S_0P5 U611 ( .A(B[14]), .X(n308) );
  SEN_INV_S_0P5 U612 ( .A(B[15]), .X(n307) );
  SEN_INV_S_0P5 U613 ( .A(B[16]), .X(n306) );
  SEN_INV_S_0P5 U614 ( .A(B[17]), .X(n305) );
  SEN_INV_S_0P5 U615 ( .A(B[18]), .X(n304) );
  SEN_INV_S_0P5 U616 ( .A(B[19]), .X(n303) );
  SEN_INV_S_0P5 U617 ( .A(B[20]), .X(n302) );
  SEN_INV_S_0P5 U618 ( .A(B[21]), .X(n301) );
  SEN_INV_S_0P5 U619 ( .A(B[22]), .X(n300) );
  SEN_INV_S_0P5 U620 ( .A(B[23]), .X(n299) );
  SEN_INV_S_0P5 U621 ( .A(B[24]), .X(n298) );
  SEN_INV_S_0P5 U622 ( .A(B[25]), .X(n297) );
  SEN_INV_S_0P5 U623 ( .A(B[26]), .X(n296) );
  SEN_INV_S_0P5 U624 ( .A(B[27]), .X(n295) );
  SEN_INV_S_0P5 U625 ( .A(B[28]), .X(n294) );
  SEN_INV_S_0P5 U626 ( .A(B[29]), .X(n293) );
  SEN_INV_S_0P5 U627 ( .A(B[30]), .X(n292) );
  SEN_INV_S_0P5 U628 ( .A(B[31]), .X(n291) );
  SEN_INV_S_0P5 U629 ( .A(INST[0]), .X(n327) );
  SEN_INV_S_0P5 U630 ( .A(INST[3]), .X(n323) );
  SEN_NR2_S_0P5 U631 ( .A1(n323), .A2(INST[0]), .X(n202) );
  SEN_INV_S_0P5 U632 ( .A(n197), .X(n324) );
  SEN_OAI221_0P5 U633 ( .A1(SEL), .A2(n193), .B1(n328), .B2(n194), .C(n195), 
        .X(n197) );
  SEN_OAI22_S_0P5 U634 ( .A1(n321), .A2(n216), .B1(B[1]), .B2(n223), .X(N157)
         );
  SEN_OAI22_S_0P5 U635 ( .A1(n320), .A2(n216), .B1(B[2]), .B2(n223), .X(N158)
         );
  SEN_OAI22_S_0P5 U636 ( .A1(n319), .A2(n216), .B1(B[3]), .B2(n223), .X(N159)
         );
  SEN_OAI22_S_0P5 U637 ( .A1(n318), .A2(n216), .B1(B[4]), .B2(n223), .X(N160)
         );
  SEN_OAI22_S_0P5 U638 ( .A1(n317), .A2(n216), .B1(B[5]), .B2(n223), .X(N161)
         );
  SEN_OAI22_S_0P5 U639 ( .A1(n316), .A2(n228), .B1(B[6]), .B2(n222), .X(N162)
         );
  SEN_OAI22_S_0P5 U640 ( .A1(n315), .A2(n228), .B1(B[7]), .B2(n222), .X(N163)
         );
  SEN_OAI22_S_0P5 U641 ( .A1(n314), .A2(n228), .B1(B[8]), .B2(n222), .X(N164)
         );
  SEN_OAI22_S_0P5 U642 ( .A1(n313), .A2(n228), .B1(B[9]), .B2(n222), .X(N165)
         );
  SEN_OAI22_S_0P5 U643 ( .A1(n312), .A2(n228), .B1(B[10]), .B2(n222), .X(N166)
         );
  SEN_OAI22_S_0P5 U644 ( .A1(n311), .A2(n228), .B1(B[11]), .B2(n222), .X(N167)
         );
  SEN_OAI22_S_0P5 U645 ( .A1(n310), .A2(n228), .B1(B[12]), .B2(n222), .X(N168)
         );
  SEN_OAI22_S_0P5 U646 ( .A1(n309), .A2(n228), .B1(B[13]), .B2(n222), .X(N169)
         );
  SEN_OAI22_S_0P5 U647 ( .A1(n308), .A2(n228), .B1(B[14]), .B2(n222), .X(N170)
         );
  SEN_OAI22_S_0P5 U648 ( .A1(n307), .A2(n228), .B1(B[15]), .B2(n222), .X(N171)
         );
  SEN_OAI22_S_0P5 U649 ( .A1(n306), .A2(n228), .B1(B[16]), .B2(n222), .X(N172)
         );
  SEN_OAI22_S_0P5 U650 ( .A1(n305), .A2(n228), .B1(B[17]), .B2(n222), .X(N173)
         );
  SEN_OAI22_S_0P5 U651 ( .A1(n304), .A2(n228), .B1(B[18]), .B2(n221), .X(N174)
         );
  SEN_OAI22_S_0P5 U652 ( .A1(n303), .A2(n227), .B1(B[19]), .B2(n221), .X(N175)
         );
  SEN_OAI22_S_0P5 U653 ( .A1(n302), .A2(n227), .B1(B[20]), .B2(n221), .X(N176)
         );
  SEN_OAI22_S_0P5 U654 ( .A1(n301), .A2(n227), .B1(B[21]), .B2(n221), .X(N177)
         );
  SEN_OAI22_S_0P5 U655 ( .A1(n300), .A2(n227), .B1(B[22]), .B2(n221), .X(N178)
         );
  SEN_OAI22_S_0P5 U656 ( .A1(n299), .A2(n227), .B1(B[23]), .B2(n221), .X(N179)
         );
  SEN_OAI22_S_0P5 U657 ( .A1(n298), .A2(n227), .B1(B[24]), .B2(n222), .X(N180)
         );
  SEN_OAI22_S_0P5 U658 ( .A1(n297), .A2(n227), .B1(B[25]), .B2(n221), .X(N181)
         );
  SEN_OAI22_S_0P5 U659 ( .A1(n296), .A2(n227), .B1(B[26]), .B2(n221), .X(N182)
         );
  SEN_OAI22_S_0P5 U660 ( .A1(n295), .A2(n227), .B1(B[27]), .B2(n221), .X(N183)
         );
  SEN_OAI22_S_0P5 U661 ( .A1(n294), .A2(n227), .B1(B[28]), .B2(n221), .X(N184)
         );
  SEN_OAI22_S_0P5 U662 ( .A1(n293), .A2(n227), .B1(B[29]), .B2(n221), .X(N185)
         );
  SEN_OAI22_S_0P5 U663 ( .A1(n292), .A2(n227), .B1(B[30]), .B2(n221), .X(N186)
         );
  SEN_OAI22_S_0P5 U664 ( .A1(n291), .A2(n227), .B1(B[31]), .B2(n221), .X(N187)
         );
endmodule

