module MADD (
	CLK, 
	A, 
	B, 
	C, 
	Z);
   input CLK;
   input [31:0] A;
   input [31:0] B;
   input [31:0] C;
   output [31:0] Z;

   // Internal wires
   wire \dp_cluster_0/N32 ;
   wire \dp_cluster_0/N291 ;
   wire \dp_cluster_0/N290 ;
   wire \dp_cluster_0/N289 ;
   wire \dp_cluster_0/N288 ;
   wire \bmul/neg15 ;
   wire \bmul/neg14 ;
   wire \bmul/two14 ;
   wire \bmul/one14 ;
   wire \bmul/neg13 ;
   wire \bmul/two13 ;
   wire \bmul/one13 ;
   wire \bmul/neg12 ;
   wire \bmul/two12 ;
   wire \bmul/one12 ;
   wire \bmul/neg11 ;
   wire \bmul/two11 ;
   wire \bmul/one11 ;
   wire \bmul/neg10 ;
   wire \bmul/two10 ;
   wire \bmul/one10 ;
   wire \bmul/neg9 ;
   wire \bmul/two9 ;
   wire \bmul/one9 ;
   wire \bmul/neg8 ;
   wire \bmul/two8 ;
   wire \bmul/one8 ;
   wire \bmul/neg7 ;
   wire \bmul/two7 ;
   wire \bmul/one7 ;
   wire \bmul/neg6 ;
   wire \bmul/two6 ;
   wire \bmul/one6 ;
   wire \bmul/neg5 ;
   wire \bmul/two5 ;
   wire \bmul/one5 ;
   wire \bmul/neg4 ;
   wire \bmul/two4 ;
   wire \bmul/neg3 ;
   wire \bmul/two3 ;
   wire \bmul/neg2 ;
   wire \bmul/neg1 ;
   wire \bmul/ppgen0/n35 ;
   wire \bmul/ppgen0/n34 ;
   wire \bmul/ppgen0/n33 ;
   wire \bmul/ppgen0/n32 ;
   wire \bmul/ppgen0/n31 ;
   wire \bmul/ppgen0/n30 ;
   wire \bmul/ppgen0/n29 ;
   wire \bmul/ppgen0/n28 ;
   wire \bmul/ppgen0/n27 ;
   wire \bmul/ppgen0/n26 ;
   wire \bmul/ppgen0/n25 ;
   wire \bmul/ppgen0/n24 ;
   wire \bmul/ppgen0/n23 ;
   wire \bmul/ppgen0/n22 ;
   wire \bmul/ppgen0/n21 ;
   wire \bmul/ppgen0/n20 ;
   wire \bmul/ppgen0/n19 ;
   wire \bmul/ppgen0/n18 ;
   wire \bmul/ppgen0/n17 ;
   wire \bmul/ppgen0/n16 ;
   wire \bmul/ppgen0/n15 ;
   wire \bmul/ppgen0/n14 ;
   wire \bmul/ppgen0/n13 ;
   wire \bmul/ppgen0/n12 ;
   wire \bmul/ppgen0/n11 ;
   wire \bmul/ppgen0/n9 ;
   wire \bmul/ppgen0/n8 ;
   wire \bmul/ppgen0/n7 ;
   wire \bmul/ppgen0/n6 ;
   wire \bmul/ppgen0/n5 ;
   wire \bmul/ppgen0/n4 ;
   wire \bmul/ppgen0/n3 ;
   wire \bmul/ppgen1/n35 ;
   wire \bmul/ppgen1/n34 ;
   wire \bmul/ppgen1/n33 ;
   wire \bmul/ppgen1/n32 ;
   wire \bmul/ppgen1/n31 ;
   wire \bmul/ppgen1/n30 ;
   wire \bmul/ppgen1/n29 ;
   wire \bmul/ppgen1/n28 ;
   wire \bmul/ppgen1/n27 ;
   wire \bmul/ppgen1/n26 ;
   wire \bmul/ppgen1/n25 ;
   wire \bmul/ppgen1/n24 ;
   wire \bmul/ppgen1/n23 ;
   wire \bmul/ppgen1/n22 ;
   wire \bmul/ppgen1/n21 ;
   wire \bmul/ppgen1/n20 ;
   wire \bmul/ppgen1/n19 ;
   wire \bmul/ppgen1/n18 ;
   wire \bmul/ppgen1/n17 ;
   wire \bmul/ppgen1/n16 ;
   wire \bmul/ppgen1/n15 ;
   wire \bmul/ppgen1/n14 ;
   wire \bmul/ppgen1/n13 ;
   wire \bmul/ppgen1/n8 ;
   wire \bmul/ppgen1/n7 ;
   wire \bmul/ppgen1/n6 ;
   wire \bmul/ppgen1/n5 ;
   wire \bmul/ppgen1/n4 ;
   wire \bmul/ppgen1/n3 ;
   wire \bmul/ppgen1/n2 ;
   wire \bmul/ppgen14/n35 ;
   wire \bmul/ppgen14/n24 ;
   wire \bmul/ppgen15/twoscomp[0] ;
   wire net2259;
   wire net2268;
   wire net2269;
   wire net82058;
   wire net82063;
   wire net82066;
   wire net82067;
   wire net82068;
   wire net82069;
   wire net82070;
   wire net82071;
   wire net82080;
   wire net82082;
   wire net82084;
   wire net82091;
   wire net82098;
   wire net82100;
   wire net82102;
   wire net82125;
   wire net82130;
   wire net82137;
   wire net82141;
   wire net82142;
   wire net82161;
   wire net82162;
   wire net82163;
   wire net82165;
   wire net82166;
   wire net82167;
   wire net82171;
   wire net82179;
   wire net82180;
   wire net82181;
   wire net82182;
   wire net82183;
   wire net82202;
   wire net82203;
   wire net82206;
   wire net82207;
   wire net82209;
   wire net82210;
   wire net82233;
   wire net82234;
   wire net82235;
   wire net82236;
   wire net82237;
   wire net82238;
   wire net82241;
   wire net82247;
   wire net82248;
   wire net82251;
   wire net82260;
   wire net82280;
   wire net82284;
   wire net82285;
   wire net82308;
   wire net82320;
   wire net82321;
   wire net82322;
   wire net82323;
   wire net82324;
   wire net82332;
   wire net82333;
   wire net82334;
   wire net82347;
   wire net82348;
   wire net82349;
   wire net82354;
   wire net82376;
   wire net82385;
   wire net82386;
   wire net82387;
   wire net82394;
   wire net82395;
   wire net82404;
   wire net82420;
   wire net82426;
   wire net82427;
   wire net82428;
   wire net82429;
   wire net82430;
   wire net82431;
   wire net82432;
   wire net82436;
   wire net82455;
   wire net82460;
   wire net82462;
   wire net82466;
   wire net82467;
   wire net82486;
   wire net82499;
   wire net82503;
   wire net82508;
   wire net82510;
   wire net82511;
   wire net82512;
   wire net82513;
   wire net82514;
   wire net82520;
   wire net82521;
   wire net82522;
   wire net82523;
   wire net82525;
   wire net82527;
   wire net82550;
   wire net82555;
   wire net82565;
   wire net82581;
   wire net82582;
   wire net82583;
   wire net82586;
   wire net82587;
   wire net82595;
   wire net82616;
   wire net82636;
   wire net82638;
   wire net82641;
   wire net82658;
   wire net82659;
   wire net82701;
   wire net82702;
   wire net82703;
   wire net82705;
   wire net82706;
   wire net82717;
   wire net82721;
   wire net82734;
   wire net82736;
   wire net82741;
   wire net82743;
   wire net82745;
   wire net82758;
   wire net82768;
   wire net82770;
   wire net82771;
   wire net82772;
   wire net82773;
   wire net82798;
   wire net82819;
   wire net82820;
   wire net82821;
   wire net82823;
   wire net82824;
   wire net82829;
   wire net82839;
   wire net82842;
   wire net82843;
   wire net82845;
   wire net82846;
   wire net82847;
   wire net82850;
   wire net82875;
   wire net82876;
   wire net82878;
   wire net82879;
   wire net82884;
   wire net82889;
   wire net82899;
   wire net82901;
   wire net82902;
   wire net82903;
   wire net82930;
   wire net82931;
   wire net82932;
   wire net82934;
   wire net82941;
   wire net82946;
   wire net82962;
   wire net82965;
   wire net82970;
   wire net82972;
   wire net82973;
   wire net82975;
   wire net82976;
   wire net82977;
   wire net82980;
   wire net82981;
   wire net82982;
   wire net82983;
   wire net82997;
   wire net82998;
   wire net83001;
   wire net83018;
   wire net83019;
   wire net83025;
   wire net83036;
   wire net83064;
   wire net83071;
   wire net83077;
   wire net83090;
   wire net83094;
   wire net83095;
   wire net83096;
   wire net83097;
   wire net83098;
   wire net83103;
   wire net83105;
   wire net83108;
   wire net83111;
   wire net83114;
   wire net83127;
   wire net83152;
   wire net83156;
   wire net83157;
   wire net83158;
   wire net83159;
   wire net83163;
   wire net83164;
   wire net83166;
   wire net83170;
   wire net83171;
   wire net83172;
   wire net83174;
   wire net83175;
   wire net83176;
   wire net83189;
   wire net83192;
   wire net83197;
   wire net83203;
   wire net83204;
   wire net83205;
   wire net83206;
   wire net83209;
   wire net83214;
   wire net83220;
   wire net83223;
   wire net83224;
   wire net83292;
   wire net83293;
   wire net83295;
   wire net83298;
   wire net83299;
   wire net83300;
   wire net83302;
   wire net83303;
   wire net83304;
   wire net83308;
   wire net83309;
   wire net83332;
   wire net83333;
   wire net83334;
   wire net83359;
   wire net83369;
   wire net83371;
   wire net83372;
   wire net83373;
   wire net83374;
   wire net83376;
   wire net83380;
   wire net83381;
   wire net83382;
   wire net83383;
   wire net83384;
   wire net83385;
   wire net83389;
   wire net83390;
   wire net83392;
   wire net83395;
   wire net83397;
   wire net83414;
   wire net83415;
   wire net83418;
   wire net83422;
   wire net83424;
   wire net83431;
   wire net83434;
   wire net83435;
   wire net83436;
   wire net83437;
   wire net83451;
   wire net83452;
   wire net83453;
   wire net83455;
   wire net83459;
   wire net83461;
   wire net83462;
   wire net83494;
   wire net83495;
   wire net83496;
   wire net83505;
   wire net83506;
   wire net83507;
   wire net83510;
   wire net83512;
   wire net83516;
   wire net83520;
   wire net83521;
   wire net83522;
   wire net83526;
   wire net83527;
   wire net83528;
   wire net83530;
   wire net83540;
   wire net83541;
   wire net83544;
   wire net83546;
   wire net83549;
   wire net83550;
   wire net83552;
   wire net83555;
   wire net83556;
   wire net83559;
   wire net83570;
   wire net83571;
   wire net83572;
   wire net83574;
   wire net83577;
   wire net83581;
   wire net83583;
   wire net83584;
   wire net83585;
   wire net83608;
   wire net83609;
   wire net83610;
   wire net83611;
   wire net83612;
   wire net83614;
   wire net83615;
   wire net83617;
   wire net83626;
   wire net83631;
   wire net83634;
   wire net83636;
   wire net83639;
   wire net83640;
   wire net83642;
   wire net83644;
   wire net83645;
   wire net83646;
   wire net83647;
   wire net83648;
   wire net83676;
   wire net83677;
   wire net83678;
   wire net83679;
   wire net83681;
   wire net83684;
   wire net83685;
   wire net83689;
   wire net83721;
   wire net83722;
   wire net83723;
   wire net83724;
   wire net83729;
   wire net83730;
   wire net83731;
   wire net83733;
   wire net83735;
   wire net83741;
   wire net83743;
   wire net83777;
   wire net83778;
   wire net83781;
   wire net83782;
   wire net83786;
   wire net83787;
   wire net83789;
   wire net83790;
   wire net83792;
   wire net83796;
   wire net83798;
   wire net83813;
   wire net83814;
   wire net83815;
   wire net83816;
   wire net83817;
   wire net83820;
   wire net83825;
   wire net83826;
   wire net83828;
   wire net83829;
   wire net83833;
   wire net83843;
   wire net83844;
   wire net83845;
   wire net83851;
   wire net83852;
   wire net83862;
   wire net83870;
   wire net83875;
   wire net83885;
   wire net83887;
   wire net83889;
   wire net83890;
   wire net83891;
   wire net83918;
   wire net83919;
   wire net83933;
   wire net83936;
   wire net83951;
   wire net83952;
   wire net83953;
   wire net83954;
   wire net83958;
   wire net83960;
   wire net83961;
   wire net83962;
   wire net83989;
   wire net83991;
   wire net83993;
   wire net83998;
   wire net83999;
   wire net84000;
   wire net84002;
   wire net84003;
   wire net84004;
   wire net84005;
   wire net84006;
   wire net84007;
   wire net84008;
   wire net84009;
   wire net84011;
   wire net84012;
   wire net84013;
   wire net84025;
   wire net84026;
   wire net84028;
   wire net84029;
   wire net84040;
   wire net84042;
   wire net84045;
   wire net84046;
   wire net84047;
   wire net84056;
   wire net84057;
   wire net84058;
   wire net84063;
   wire net84066;
   wire net84067;
   wire net84068;
   wire net84081;
   wire net84106;
   wire net84108;
   wire net84111;
   wire net84115;
   wire net84116;
   wire net84117;
   wire net84118;
   wire net84119;
   wire net84121;
   wire net84146;
   wire net84147;
   wire net84148;
   wire net84150;
   wire net84152;
   wire net84153;
   wire net84156;
   wire net84157;
   wire net84160;
   wire net84177;
   wire net84186;
   wire net84187;
   wire net84189;
   wire net84191;
   wire net84192;
   wire net84193;
   wire net84200;
   wire net84208;
   wire net84217;
   wire net84218;
   wire net84220;
   wire net84221;
   wire net84223;
   wire net84226;
   wire net84229;
   wire net84230;
   wire net84231;
   wire net84232;
   wire net84233;
   wire net84235;
   wire net84236;
   wire net84237;
   wire net84238;
   wire net84239;
   wire net84241;
   wire net84246;
   wire net84248;
   wire net84271;
   wire net84272;
   wire net84276;
   wire net84281;
   wire net84284;
   wire net84286;
   wire net84358;
   wire net84359;
   wire net84362;
   wire net84364;
   wire net84365;
   wire net84366;
   wire net84370;
   wire net84371;
   wire net84372;
   wire net84378;
   wire net84384;
   wire net84385;
   wire net84395;
   wire net84404;
   wire net84405;
   wire net84407;
   wire net84408;
   wire net84409;
   wire net84411;
   wire net84412;
   wire net84413;
   wire net84414;
   wire net84415;
   wire net84425;
   wire net84433;
   wire net84435;
   wire net84437;
   wire net84441;
   wire net84442;
   wire net84445;
   wire net84448;
   wire net84449;
   wire net84451;
   wire net84471;
   wire net84592;
   wire net84588;
   wire net84586;
   wire net84600;
   wire net84634;
   wire net84636;
   wire net84650;
   wire net84654;
   wire net84734;
   wire net85046;
   wire net85071;
   wire net85334;
   wire net85748;
   wire net85815;
   wire net85838;
   wire net85837;
   wire net85880;
   wire net85897;
   wire net85926;
   wire net85984;
   wire net86002;
   wire net86010;
   wire net86023;
   wire net86022;
   wire net86076;
   wire net86086;
   wire net86124;
   wire net86213;
   wire net86258;
   wire net86257;
   wire net86273;
   wire net86274;
   wire net86279;
   wire net86299;
   wire net86306;
   wire net86321;
   wire net86332;
   wire net86333;
   wire net86390;
   wire net86455;
   wire net86454;
   wire net86459;
   wire net86466;
   wire net86491;
   wire net86494;
   wire net86493;
   wire net86517;
   wire net86534;
   wire net86655;
   wire net86698;
   wire net86699;
   wire net87351;
   wire net87543;
   wire net87542;
   wire net87541;
   wire net87547;
   wire net87546;
   wire net87549;
   wire net87627;
   wire net87761;
   wire net87763;
   wire net87762;
   wire net87769;
   wire net87787;
   wire net87786;
   wire net87791;
   wire net87790;
   wire net87795;
   wire net87800;
   wire net87799;
   wire net87814;
   wire net87813;
   wire net87822;
   wire net87821;
   wire net87828;
   wire net87827;
   wire net87846;
   wire net87845;
   wire net87844;
   wire net87990;
   wire net88056;
   wire net88080;
   wire net88079;
   wire net88078;
   wire net88089;
   wire net88108;
   wire net88113;
   wire net87837;
   wire net86446;
   wire net82822;
   wire net82640;
   wire net87836;
   wire net85257;
   wire net82859;
   wire net82858;
   wire net82856;
   wire net82855;
   wire net82854;
   wire net83632;
   wire net83513;
   wire net83387;
   wire net83370;
   wire net83169;
   wire net86078;
   wire net85173;
   wire net84450;
   wire net84410;
   wire net84391;
   wire net83830;
   wire net83740;
   wire net82999;
   wire net89933;
   wire net89992;
   wire net90258;
   wire net90316;
   wire net90615;
   wire net90631;
   wire net90705;
   wire net90704;
   wire net90746;
   wire net90814;
   wire net90815;
   wire net90868;
   wire net90880;
   wire net90884;
   wire net90917;
   wire net90993;
   wire net91024;
   wire net91053;
   wire net91065;
   wire net91110;
   wire net91120;
   wire net91426;
   wire net91419;
   wire net91418;
   wire net91410;
   wire net91408;
   wire net91406;
   wire net91390;
   wire net91386;
   wire net91363;
   wire net91564;
   wire net84059;
   wire net83301;
   wire net83534;
   wire net83454;
   wire net82201;
   wire net82061;
   wire net82060;
   wire net87798;
   wire net87797;
   wire net91415;
   wire net91407;
   wire net87101;
   wire net82674;
   wire net82516;
   wire net82515;
   wire net82197;
   wire net82196;
   wire net82195;
   wire net82193;
   wire net84202;
   wire net84201;
   wire net83965;
   wire net83578;
   wire net87796;
   wire net86477;
   wire net83607;
   wire net83331;
   wire net83329;
   wire net87100;
   wire net82390;
   wire net82389;
   wire net82194;
   wire net82190;
   wire net82189;
   wire net82188;
   wire net82187;
   wire net82186;
   wire net82075;
   wire net85252;
   wire net82336;
   wire net82335;
   wire net82055;
   wire net86385;
   wire net83547;
   wire net83538;
   wire net83537;
   wire net83535;
   wire net83297;
   wire net84251;
   wire net84073;
   wire net84001;
   wire net94064;
   wire net94058;
   wire net94057;
   wire net94132;
   wire net94217;
   wire net94287;
   wire net94314;
   wire net94322;
   wire net94321;
   wire net94359;
   wire net94383;
   wire net84288;
   wire net84274;
   wire net83153;
   wire net82939;
   wire net82938;
   wire net82936;
   wire net82935;
   wire net84361;
   wire net84357;
   wire net84356;
   wire net84355;
   wire net84353;
   wire net84352;
   wire net84351;
   wire net84350;
   wire net84227;
   wire net84418;
   wire net84417;
   wire net84393;
   wire net84392;
   wire net84354;
   wire net84730;
   wire net84322;
   wire net84283;
   wire net84228;
   wire net84159;
   wire net95575;
   wire net95563;
   wire net95561;
   wire net95559;
   wire net95557;
   wire net95543;
   wire net95536;
   wire net95509;
   wire net95748;
   wire net95774;
   wire net95817;
   wire net95846;
   wire net95872;
   wire net95928;
   wire net95993;
   wire net83964;
   wire net83582;
   wire net83566;
   wire net83565;
   wire net85351;
   wire net83580;
   wire net83573;
   wire net97222;
   wire net97350;
   wire net97377;
   wire net97397;
   wire net91392;
   wire net82564;
   wire net82562;
   wire net82457;
   wire net82079;
   wire net82078;
   wire net82077;
   wire net82076;
   wire net82074;
   wire net91413;
   wire net82454;
   wire net82246;
   wire net82243;
   wire net91405;
   wire net91399;
   wire net91398;
   wire net91397;
   wire net91396;
   wire net90740;
   wire net90738;
   wire net90737;
   wire net86266;
   wire net85931;
   wire net82245;
   wire net82244;
   wire net82173;
   wire net82083;
   wire net82057;
   wire net98319;
   wire net98293;
   wire net84732;
   wire net84394;
   wire net94176;
   wire net86483;
   wire net82831;
   wire net83863;
   wire net83168;
   wire net84443;
   wire net86498;
   wire net86382;
   wire net86381;
   wire net82383;
   wire net82302;
   wire net96981;
   wire net83498;
   wire net83497;
   wire net83413;
   wire net83412;
   wire net83408;
   wire net82967;
   wire net89993;
   wire net84275;
   wire net84273;
   wire net84196;
   wire net84183;
   wire net83861;
   wire net90668;
   wire net88104;
   wire net88103;
   wire net86553;
   wire net86518;
   wire net82836;
   wire net82833;
   wire net82827;
   wire net82634;
   wire net82317;
   wire net82315;
   wire net82313;
   wire net82309;
   wire net82062;
   wire net82059;
   wire net82056;
   wire net83849;
   wire net83848;
   wire net83846;
   wire net83630;
   wire net83629;
   wire net83627;
   wire net83508;
   wire net83499;
   wire net100921;
   wire net100928;
   wire net101248;
   wire net101261;
   wire net101269;
   wire net82124;
   wire net82123;
   wire net82114;
   wire net102542;
   wire net102677;
   wire net103418;
   wire net88015;
   wire net88014;
   wire net87948;
   wire net87947;
   wire net87946;
   wire net87944;
   wire net87943;
   wire net86468;
   wire net82639;
   wire net82319;
   wire net82316;
   wire net82311;
   wire net82310;
   wire net82306;
   wire net82305;
   wire net82304;
   wire net82065;
   wire net82052;
   wire net82051;
   wire net82050;
   wire net82049;
   wire net82047;
   wire net82046;
   wire net82044;
   wire net82043;
   wire net82042;
   wire net82041;
   wire net86557;
   wire net86556;
   wire net83076;
   wire net83072;
   wire net82937;
   wire net82857;
   wire net82838;
   wire net82742;
   wire net83165;
   wire net83070;
   wire net86560;
   wire net86559;
   wire net84110;
   wire net84107;
   wire net83649;
   wire net83525;
   wire net83524;
   wire net83523;
   wire net83000;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;
   wire n890;
   wire n891;
   wire n892;
   wire n893;
   wire n894;
   wire n895;
   wire n896;
   wire n897;
   wire n898;
   wire n899;
   wire n900;
   wire n901;
   wire n902;
   wire n903;
   wire n904;
   wire n905;
   wire n906;
   wire n907;
   wire n908;
   wire n909;
   wire n910;
   wire n911;
   wire n912;
   wire n913;
   wire n914;
   wire n915;
   wire n916;
   wire n917;
   wire n918;
   wire n919;
   wire n920;
   wire n921;
   wire n922;
   wire n923;
   wire n924;
   wire n925;
   wire n926;
   wire n927;
   wire n928;
   wire n929;
   wire n930;
   wire n931;
   wire n932;
   wire n933;
   wire n934;
   wire n935;
   wire n936;
   wire n937;
   wire n938;
   wire n939;
   wire n940;
   wire n941;
   wire n942;
   wire n943;
   wire n944;
   wire n945;
   wire n946;
   wire n947;
   wire n948;
   wire n949;
   wire n950;
   wire n951;
   wire n952;
   wire n953;
   wire n954;
   wire n955;
   wire n956;
   wire n957;
   wire n958;
   wire n959;
   wire n960;
   wire n961;
   wire n962;
   wire n963;
   wire n964;
   wire n965;
   wire n966;
   wire n967;
   wire n968;
   wire n969;
   wire n970;
   wire n971;
   wire n972;
   wire n973;
   wire n974;
   wire n975;
   wire n976;
   wire n977;
   wire n978;
   wire n979;
   wire n980;
   wire n981;
   wire n982;
   wire n983;
   wire n984;
   wire n985;
   wire n986;
   wire n987;
   wire n988;
   wire n989;
   wire n990;
   wire n991;
   wire n992;
   wire n993;
   wire n994;
   wire n995;
   wire n996;
   wire n997;
   wire n998;
   wire n999;
   wire n1000;
   wire n1001;
   wire n1002;
   wire n1003;
   wire n1004;
   wire n1005;
   wire n1006;
   wire n1007;
   wire n1008;
   wire n1009;
   wire n1010;
   wire n1011;
   wire n1012;
   wire n1013;
   wire n1014;
   wire n1015;
   wire n1016;
   wire n1017;
   wire n1018;
   wire n1019;
   wire n1020;
   wire n1021;
   wire n1022;
   wire n1023;
   wire n1024;
   wire n1025;
   wire n1026;
   wire n1027;
   wire n1028;
   wire n1029;
   wire n1030;
   wire n1031;
   wire n1032;
   wire n1033;
   wire n1034;
   wire n1035;
   wire n1036;
   wire n1037;
   wire n1038;
   wire n1039;
   wire n1040;
   wire n1041;
   wire n1042;
   wire n1043;
   wire n1044;
   wire n1045;
   wire n1046;
   wire n1047;
   wire n1048;
   wire n1049;
   wire n1050;
   wire n1051;
   wire n1052;
   wire n1053;
   wire n1054;
   wire n1055;
   wire n1056;
   wire n1057;
   wire n1058;
   wire n1059;
   wire n1060;
   wire n1061;
   wire n1062;
   wire n1063;
   wire n1064;
   wire n1065;
   wire n1066;
   wire n1067;
   wire n1068;
   wire n1069;
   wire n1070;
   wire n1071;
   wire n1072;
   wire n1073;
   wire n1074;
   wire n1075;
   wire n1076;
   wire n1077;
   wire n1078;
   wire n1079;
   wire n1080;
   wire n1081;
   wire n1082;
   wire n1083;
   wire n1084;
   wire n1085;
   wire n1086;
   wire n1087;
   wire n1088;
   wire n1089;
   wire n1090;
   wire n1091;
   wire n1092;
   wire n1093;
   wire n1094;
   wire n1095;
   wire n1096;
   wire n1097;
   wire n1098;
   wire n1099;
   wire n1100;
   wire n1101;
   wire n1102;
   wire n1103;
   wire n1104;
   wire n1105;
   wire n1106;
   wire n1107;
   wire n1108;
   wire n1109;
   wire n1110;
   wire n1111;
   wire n1112;
   wire n1113;
   wire n1114;
   wire n1115;
   wire n1116;
   wire n1117;
   wire n1118;
   wire n1119;
   wire n1120;
   wire n1121;
   wire n1122;
   wire n1123;
   wire n1124;
   wire n1125;
   wire n1126;
   wire n1127;
   wire n1128;
   wire n1129;
   wire n1130;
   wire n1131;
   wire n1132;
   wire n1133;
   wire n1134;
   wire n1135;
   wire n1136;
   wire n1137;
   wire n1138;
   wire n1139;
   wire n1140;
   wire n1141;
   wire n1142;
   wire n1143;
   wire n1144;
   wire n1145;
   wire n1146;
   wire n1147;
   wire n1148;
   wire n1149;
   wire n1150;
   wire n1151;
   wire n1152;
   wire n1153;
   wire n1154;
   wire n1155;
   wire n1156;
   wire n1157;
   wire n1158;
   wire n1159;
   wire n1160;
   wire n1161;
   wire n1162;
   wire n1163;
   wire n1164;
   wire n1165;
   wire n1166;
   wire n1167;
   wire n1168;
   wire n1169;
   wire n1170;
   wire n1171;
   wire n1172;
   wire n1173;
   wire n1174;
   wire n1175;
   wire n1176;
   wire n1177;
   wire n1178;
   wire n1179;
   wire n1180;
   wire n1181;
   wire n1182;
   wire n1183;
   wire n1184;
   wire n1185;
   wire n1186;
   wire n1187;
   wire n1188;
   wire n1189;
   wire n1190;
   wire n1191;
   wire n1192;
   wire n1193;
   wire n1194;
   wire n1195;
   wire n1196;
   wire n1197;
   wire n1198;
   wire n1199;
   wire n1200;
   wire n1201;
   wire n1202;
   wire n1203;
   wire n1204;
   wire n1205;
   wire n1206;
   wire n1207;
   wire n1208;
   wire n1209;
   wire n1210;
   wire n1211;
   wire n1212;
   wire n1213;
   wire n1214;
   wire n1215;
   wire n1216;
   wire n1217;
   wire n1218;
   wire n1219;
   wire n1220;
   wire n1221;
   wire n1222;
   wire n1223;
   wire n1224;
   wire n1225;
   wire n1226;
   wire n1227;
   wire n1228;
   wire n1229;
   wire n1230;
   wire n1231;
   wire n1232;
   wire n1233;
   wire n1234;
   wire n1235;
   wire n1236;
   wire n1237;
   wire n1238;
   wire n1239;
   wire n1240;
   wire n1241;
   wire n1242;
   wire n1243;
   wire n1244;
   wire n1245;
   wire n1246;
   wire n1247;
   wire n1248;
   wire n1249;
   wire n1250;
   wire n1251;
   wire n1252;
   wire n1253;
   wire n1254;
   wire n1255;
   wire n1256;
   wire n1257;
   wire n1258;
   wire n1259;
   wire n1260;
   wire n1261;
   wire n1262;
   wire n1263;
   wire n1264;
   wire n1265;
   wire n1266;
   wire n1267;
   wire n1268;
   wire n1269;
   wire n1270;
   wire n1271;
   wire n1272;
   wire n1273;
   wire n1274;
   wire n1275;
   wire n1276;
   wire n1277;
   wire n1278;
   wire n1279;
   wire n1280;
   wire n1281;
   wire n1282;
   wire n1283;
   wire n1284;
   wire n1285;
   wire n1286;
   wire n1287;
   wire n1288;
   wire n1289;
   wire n1290;
   wire n1291;
   wire n1292;
   wire n1293;
   wire n1294;
   wire n1295;
   wire n1296;
   wire n1297;
   wire n1298;
   wire n1299;
   wire n1300;
   wire n1301;
   wire n1302;
   wire n1303;
   wire n1304;
   wire n1305;
   wire n1306;
   wire n1307;
   wire n1308;
   wire n1309;
   wire n1310;
   wire n1311;
   wire n1312;
   wire n1313;
   wire n1314;
   wire n1315;
   wire n1316;
   wire n1317;
   wire n1318;
   wire n1319;
   wire n1320;
   wire n1321;
   wire n1322;
   wire n1323;
   wire n1324;
   wire n1325;
   wire n1326;
   wire n1327;
   wire n1328;
   wire n1329;
   wire n1330;
   wire n1331;
   wire n1332;
   wire n1333;
   wire n1334;
   wire n1335;
   wire n1336;
   wire n1337;
   wire n1338;
   wire n1339;
   wire n1340;
   wire n1341;
   wire n1342;
   wire n1343;
   wire n1344;
   wire n1345;
   wire n1346;
   wire n1347;
   wire n1348;
   wire n1349;
   wire n1350;
   wire n1351;
   wire n1352;
   wire n1353;
   wire n1354;
   wire n1355;
   wire n1356;
   wire n1357;
   wire n1358;
   wire n1359;
   wire n1360;
   wire n1361;
   wire n1362;
   wire n1363;
   wire n1364;
   wire n1365;
   wire n1366;
   wire n1367;
   wire n1368;
   wire n1369;
   wire n1370;
   wire n1371;
   wire n1372;
   wire n1373;
   wire n1374;
   wire n1375;
   wire n1376;
   wire n1377;
   wire n1378;
   wire n1379;
   wire n1380;
   wire n1381;
   wire n1382;
   wire n1383;
   wire n1384;
   wire n1385;
   wire n1386;
   wire n1387;
   wire n1388;
   wire n1389;
   wire n1390;
   wire n1391;
   wire n1392;
   wire n1393;
   wire n1394;
   wire n1395;
   wire n1396;
   wire n1397;
   wire n1398;
   wire n1399;
   wire n1400;
   wire n1401;
   wire n1402;
   wire n1403;
   wire n1404;
   wire n1405;
   wire n1406;
   wire n1407;
   wire n1408;
   wire n1409;
   wire n1410;
   wire n1411;
   wire n1412;
   wire n1413;
   wire n1414;
   wire n1415;
   wire n1416;
   wire n1417;
   wire n1418;
   wire n1419;
   wire n1420;
   wire n1421;
   wire n1422;
   wire n1423;
   wire n1424;
   wire n1425;
   wire n1426;
   wire n1427;
   wire n1428;
   wire n1429;
   wire n1430;
   wire n1431;
   wire n1432;
   wire n1433;
   wire n1434;
   wire n1435;
   wire n1436;
   wire n1437;
   wire n1438;
   wire n1439;
   wire n1440;
   wire n1441;
   wire n1442;
   wire n1443;
   wire n1444;
   wire n1445;
   wire n1446;
   wire n1447;
   wire n1448;
   wire n1449;
   wire n1450;
   wire n1451;
   wire n1452;
   wire n1453;
   wire n1454;
   wire n1455;
   wire n1456;
   wire n1457;
   wire n1458;
   wire n1459;
   wire n1460;
   wire n1461;
   wire n1462;
   wire n1463;
   wire n1464;
   wire n1465;
   wire n1466;
   wire n1467;
   wire n1468;
   wire n1469;
   wire n1470;
   wire n1471;
   wire n1472;
   wire n1473;
   wire n1474;
   wire n1475;
   wire n1476;
   wire n1477;
   wire n1478;
   wire n1479;
   wire n1480;
   wire n1481;
   wire n1482;
   wire n1483;
   wire n1484;
   wire n1485;
   wire n1486;
   wire n1487;
   wire n1488;
   wire n1489;
   wire n1490;
   wire n1491;
   wire n1492;
   wire n1493;
   wire n1494;
   wire n1495;
   wire n1496;
   wire n1497;
   wire n1498;
   wire n1499;
   wire n1500;
   wire n1501;
   wire n1502;
   wire n1503;
   wire n1504;
   wire n1505;
   wire n1506;
   wire n1507;
   wire n1508;
   wire n1509;
   wire n1510;
   wire n1511;
   wire n1512;
   wire n1513;
   wire n1514;
   wire n1515;
   wire n1517;
   wire n1518;
   wire n1519;
   wire n1520;
   wire n1521;
   wire n1522;
   wire n1523;
   wire n1524;
   wire n1525;
   wire n1526;
   wire n1527;
   wire n1528;
   wire n1529;
   wire n1530;
   wire n1531;
   wire n1532;
   wire n1533;
   wire n1534;
   wire n1535;
   wire n1536;
   wire n1537;
   wire n1538;
   wire n1539;
   wire n1540;
   wire n1541;
   wire n1542;
   wire n1543;
   wire n1544;
   wire n1545;
   wire n1546;
   wire n1547;
   wire n1548;
   wire n1549;
   wire n1550;
   wire n1551;
   wire n1552;
   wire n1553;
   wire n1554;
   wire n1555;
   wire n1556;
   wire n1557;
   wire n1558;
   wire n1559;
   wire n1560;
   wire n1561;
   wire n1562;
   wire n1563;
   wire n1564;
   wire n1565;
   wire n1566;
   wire n1572;
   wire n1573;
   wire n1574;
   wire n1575;
   wire n1576;
   wire n1577;
   wire n1578;
   wire n1579;
   wire n1580;
   wire n1581;
   wire n1582;
   wire n1583;
   wire n1584;
   wire n1585;
   wire n1586;
   wire n1587;
   wire n1588;
   wire n1589;
   wire n1590;
   wire n1591;
   wire n1592;
   wire n1593;
   wire n1594;
   wire n1595;
   wire n1596;
   wire n1597;
   wire n1598;
   wire n1599;
   wire n1600;
   wire n1601;
   wire n1602;
   wire n1603;
   wire n1604;
   wire n1605;
   wire n1607;
   wire n1608;
   wire n1609;
   wire n1610;
   wire n1611;
   wire n1612;
   wire n1613;
   wire n1614;
   wire n1619;
   wire n1620;
   wire n1621;
   wire n1622;
   wire n1623;
   wire n1624;
   wire n1625;
   wire n1626;
   wire n1627;
   wire n1628;
   wire n1629;
   wire n1630;
   wire n1631;
   wire n1632;
   wire n1633;
   wire n1634;
   wire n1635;
   wire n1636;
   wire n1637;
   wire n1638;
   wire n1639;
   wire n1640;
   wire n1641;
   wire n1642;
   wire n1643;
   wire n1644;
   wire n1645;
   wire n1646;
   wire n1647;
   wire n1648;
   wire n1649;
   wire n1650;
   wire n1651;
   wire n1652;
   wire n1653;
   wire n1654;
   wire n1655;
   wire n1656;
   wire n1657;
   wire n1658;
   wire n1659;
   wire n1660;
   wire n1661;
   wire n1662;
   wire n1663;
   wire n1664;
   wire n1665;
   wire n1666;
   wire n1667;
   wire n1668;
   wire n1669;
   wire n1671;
   wire n1672;
   wire n1673;
   wire n1674;
   wire n1675;
   wire n1676;
   wire n1677;
   wire n1678;
   wire n1679;
   wire n1680;
   wire n1681;
   wire n1682;
   wire n1683;
   wire n1684;
   wire n1685;
   wire n1686;
   wire n1687;
   wire n1688;
   wire n1689;
   wire n1690;
   wire n1691;
   wire n1692;
   wire n1693;
   wire n1694;
   wire n1695;
   wire n1696;
   wire n1697;
   wire n1698;
   wire n1699;
   wire n1700;
   wire n1701;
   wire n1702;
   wire n1703;
   wire n1704;
   wire n1705;
   wire n1706;
   wire n1707;
   wire n1708;
   wire n1709;
   wire n1710;
   wire n1711;
   wire n1712;
   wire n1713;
   wire n1714;
   wire n1715;
   wire n1716;
   wire n1717;
   wire n1718;
   wire n1719;
   wire n1720;
   wire n1721;
   wire n1722;
   wire n1723;
   wire n1724;
   wire n1725;
   wire n1726;
   wire n1727;
   wire n1728;
   wire n1729;
   wire n1730;
   wire n1731;
   wire n1732;
   wire n1733;
   wire n1734;
   wire n1735;
   wire n1736;
   wire n1737;
   wire n1738;
   wire n1739;
   wire n1740;
   wire n1741;
   wire n1742;
   wire n1743;
   wire n1744;
   wire n1745;
   wire n1746;
   wire n1747;
   wire n1748;
   wire n1749;
   wire n1750;
   wire n1751;
   wire n1752;
   wire n1753;
   wire n1754;
   wire n1755;
   wire n1756;
   wire n1757;
   wire n1758;
   wire n1759;
   wire n1760;
   wire n1761;
   wire n1762;
   wire n1763;
   wire n1764;
   wire n1765;
   wire n1766;
   wire n1767;
   wire n1768;
   wire n1769;
   wire n1770;
   wire n1771;
   wire n1772;
   wire n1773;
   wire n1774;
   wire n1775;
   wire n1776;
   wire n1777;
   wire n1778;
   wire n1779;
   wire n1780;
   wire n1781;
   wire n1782;
   wire n1783;
   wire n1784;
   wire n1785;
   wire n1786;
   wire n1787;
   wire n1788;
   wire n1789;
   wire n1790;
   wire n1791;
   wire n1792;
   wire n1793;
   wire n1794;
   wire n1795;
   wire n1796;
   wire n1797;
   wire n1798;
   wire n1799;
   wire n1800;
   wire n1801;
   wire n1802;
   wire n1803;
   wire n1804;
   wire n1805;
   wire n1806;
   wire n1807;
   wire n1808;
   wire n1809;
   wire n1810;
   wire n1811;
   wire n1812;
   wire n1813;
   wire n1814;
   wire n1815;
   wire n1816;
   wire n1817;
   wire n1836;
   wire n1837;
   wire n1838;
   wire n1839;
   wire n1840;
   wire n1841;
   wire n1842;
   wire n1843;
   wire n1844;
   wire n1845;
   wire n1846;
   wire n1847;
   wire n1848;
   wire n1849;
   wire n1850;
   wire n1851;
   wire n1852;
   wire n1853;
   wire n1854;
   wire n1855;
   wire n1856;
   wire n1857;
   wire n1858;
   wire n1859;
   wire n1860;
   wire n1861;
   wire n1862;
   wire n1863;
   wire n1864;
   wire n1865;
   wire n1866;
   wire n1867;
   wire n1868;
   wire n1869;
   wire n1870;
   wire n1871;
   wire n1872;
   wire n1873;
   wire n1874;
   wire n1875;
   wire n1876;
   wire n1877;
   wire n1878;
   wire n1879;
   wire n1880;
   wire n1881;
   wire n1882;
   wire n1883;
   wire n1884;
   wire n1885;
   wire n1886;
   wire n1887;
   wire n1888;
   wire n1889;
   wire n1890;
   wire n1891;
   wire n1892;
   wire n1893;
   wire n1894;
   wire n1895;
   wire n1896;
   wire n1897;
   wire n1898;
   wire n1899;
   wire n1900;
   wire n1901;
   wire n1902;
   wire n1903;
   wire n1904;
   wire n1905;
   wire n1906;
   wire n1907;
   wire n1908;
   wire n1909;
   wire n1910;
   wire n1911;
   wire n1912;
   wire n1913;
   wire n1914;
   wire n1915;
   wire n1916;
   wire n1917;
   wire n1918;
   wire n1919;
   wire n1920;
   wire n1921;
   wire n1922;
   wire n1923;
   wire n1924;
   wire n1925;
   wire n1926;
   wire n1927;
   wire n1928;
   wire n1929;
   wire n1930;
   wire n1931;
   wire n1932;
   wire n1933;
   wire n1934;
   wire n1935;
   wire n1936;
   wire n1937;
   wire n1938;
   wire n1939;
   wire n1940;
   wire n1941;
   wire n1942;
   wire n1943;
   wire n1944;
   wire n1945;
   wire n1946;
   wire n1947;
   wire n1948;
   wire n1949;
   wire n1950;
   wire n1951;
   wire n1952;
   wire n1953;
   wire n1954;
   wire n1955;
   wire n1956;
   wire n1957;
   wire n1958;
   wire n1959;
   wire n1960;
   wire n1961;
   wire n1962;
   wire n1963;
   wire n1964;
   wire n1965;
   wire n1966;
   wire n1967;
   wire n1968;
   wire n1969;
   wire n1970;
   wire n1971;
   wire n1972;
   wire n1973;
   wire n1974;
   wire n1975;
   wire n1976;
   wire n1977;
   wire n1978;
   wire n1979;
   wire n1980;
   wire n1981;
   wire n1982;
   wire n1983;
   wire n1984;
   wire n1985;
   wire n1986;
   wire n1987;
   wire n1988;
   wire n1989;
   wire n1990;
   wire n1991;
   wire n1992;
   wire n1993;
   wire n1994;
   wire n1995;
   wire n1996;
   wire n1997;
   wire n1998;
   wire n1999;
   wire n2000;
   wire n2001;
   wire n2002;
   wire n2003;
   wire n2004;
   wire n2005;
   wire n2006;
   wire n2007;
   wire n2008;
   wire n2009;
   wire n2010;
   wire n2011;
   wire n2012;
   wire n2013;
   wire n2014;
   wire n2015;
   wire n2016;
   wire n2017;
   wire n2018;
   wire n2019;
   wire n2020;
   wire n2021;
   wire n2022;
   wire n2023;
   wire n2024;
   wire n2025;
   wire n2026;
   wire n2027;
   wire n2028;
   wire n2029;
   wire n2030;
   wire n2031;
   wire n2032;
   wire n2033;
   wire n2034;
   wire n2035;
   wire net91394;
   wire net82122;
   wire net82119;
   wire net90456;
   wire net82120;
   wire net82116;
   wire net82115;
   wire net82088;
   wire net82087;
   wire net82085;
   wire net82073;
   wire net82072;
   wire net82064;
   wire n178;
   wire n177;
   wire n176;
   wire n175;
   wire n174;
   wire n173;
   wire n172;
   wire n171;
   wire n170;
   wire n169;
   wire n168;
   wire n167;
   wire n166;
   wire n165;
   wire n164;
   wire n163;
   wire n2036;
   wire n2037;
   wire n2038;
   wire n2039;
   wire n2040;
   wire n2041;
   wire n2042;
   wire n2043;
   wire n2044;
   wire n2045;
   wire n2046;
   wire n2047;
   wire n2048;
   wire n2049;
   wire n2050;
   wire n2051;
   wire n2052;
   wire n2053;
   wire n2054;
   wire n2055;
   wire n2056;
   wire n2057;
   wire n2058;
   wire n2059;
   wire n2060;
   wire n2061;
   wire n2062;
   wire n2063;
   wire n2064;
   wire n2065;
   wire n2066;
   wire n2067;
   wire n2068;
   wire n2069;
   wire n2070;
   wire n2071;
   wire n2072;
   wire n2073;
   wire n2074;
   wire n2075;
   wire n2076;
   wire n2077;
   wire n2078;
   wire n2079;
   wire n2080;
   wire n2081;
   wire n2082;
   wire n2083;
   wire n2084;
   wire n2085;
   wire n2086;
   wire n2087;
   wire n2088;
   wire n2089;
   wire n2090;
   wire n2091;
   wire n2092;
   wire n2093;
   wire n2094;
   wire n2095;
   wire n2096;
   wire n2097;
   wire n2098;
   wire n2099;
   wire n2100;
   wire n2101;
   wire [35:0] pprow0;
   wire [34:0] pprow1;
   wire [34:0] pprow2;
   wire [34:0] pprow3;
   wire [34:0] pprow4;
   wire [34:0] pprow5;
   wire [34:0] pprow6;
   wire [34:0] pprow7;
   wire [34:0] pprow8;
   wire [34:0] pprow9;
   wire [34:0] pprow10;
   wire [34:0] pprow11;
   wire [34:0] pprow12;
   wire [34:0] pprow13;
   wire [35:0] pprow14;
   wire [31:0] pprow0_qual;
   wire [29:0] pprow1_qual;
   wire [25:0] pprow2_qual;
   wire [23:0] pprow3_qual;
   wire [21:0] pprow4_qual;
   wire [19:0] pprow5_qual;
   wire [17:0] pprow6_qual;
   wire [15:0] pprow7_qual;
   wire [13:0] pprow8_qual;
   wire [11:0] pprow9_qual;
   wire [9:0] pprow10_qual;
   wire [7:0] pprow11_qual;
   wire [5:0] pprow12_qual;
   wire [3:0] pprow13_qual;
   wire [1:0] pprow14_qual;

   assign \dp_cluster_0/N32  = A[1] ;
   assign Z[3] = \dp_cluster_0/N291  ;
   assign Z[2] = \dp_cluster_0/N290  ;
   assign Z[1] = \dp_cluster_0/N289  ;
   assign Z[0] = \dp_cluster_0/N288  ;
   assign \bmul/neg15  = A[31] ;
   assign \bmul/neg14  = A[29] ;
   assign \bmul/neg13  = A[27] ;
   assign \bmul/neg12  = A[25] ;
   assign \bmul/neg11  = A[23] ;
   assign \bmul/neg10  = A[21] ;
   assign \bmul/neg9  = A[19] ;
   assign \bmul/neg8  = A[17] ;
   assign \bmul/neg7  = A[15] ;
   assign \bmul/neg6  = A[13] ;
   assign \bmul/neg5  = A[11] ;
   assign \bmul/neg4  = A[9] ;
   assign \bmul/neg3  = A[7] ;
   assign \bmul/neg2  = A[5] ;
   assign \bmul/neg1  = A[3] ;
   assign \bmul/ppgen15/twoscomp[0]  = B[0] ;

   SEN_FDPQ_4 \pprow1_qual_reg[15]  (.Q(pprow1_qual[15]), 
	.D(pprow1[15]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[13]  (.Q(pprow1_qual[13]), 
	.D(pprow1[13]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[12]  (.Q(pprow1_qual[12]), 
	.D(pprow1[12]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[9]  (.Q(pprow1_qual[9]), 
	.D(pprow1[9]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[8]  (.Q(pprow1_qual[8]), 
	.D(pprow1[8]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[4]  (.Q(pprow1_qual[4]), 
	.D(pprow1[4]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[3]  (.Q(pprow1_qual[3]), 
	.D(pprow1[3]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[2]  (.Q(pprow1_qual[2]), 
	.D(pprow1[2]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[0]  (.Q(pprow1_qual[0]), 
	.D(pprow1[0]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[6]  (.Q(pprow2_qual[6]), 
	.D(pprow2[6]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[5]  (.Q(pprow2_qual[5]), 
	.D(pprow2[5]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[4]  (.Q(pprow2_qual[4]), 
	.D(pprow2[4]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[3]  (.Q(pprow2_qual[3]), 
	.D(pprow2[3]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow3_qual_reg[5]  (.Q(pprow3_qual[5]), 
	.D(pprow3[5]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow3_qual_reg[3]  (.Q(pprow3_qual[3]), 
	.D(pprow3[3]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow3_qual_reg[1]  (.Q(pprow3_qual[1]), 
	.D(pprow3[1]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow3_qual_reg[0]  (.Q(pprow3_qual[0]), 
	.D(pprow3[0]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow5_qual_reg[5]  (.Q(pprow5_qual[5]), 
	.D(pprow5[5]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow5_qual_reg[3]  (.Q(pprow5_qual[3]), 
	.D(pprow5[3]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow5_qual_reg[0]  (.Q(pprow5_qual[0]), 
	.D(pprow5[0]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow6_qual_reg[2]  (.Q(pprow6_qual[2]), 
	.D(pprow6[2]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow6_qual_reg[0]  (.Q(pprow6_qual[0]), 
	.D(pprow6[0]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow7_qual_reg[0]  (.Q(pprow7_qual[0]), 
	.D(pprow7[0]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow3_qual_reg[2]  (.Q(pprow3_qual[2]), 
	.D(pprow3[2]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[11]  (.Q(pprow1_qual[11]), 
	.D(pprow1[11]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[10]  (.Q(pprow1_qual[10]), 
	.D(pprow1[10]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow5_qual_reg[1]  (.Q(pprow5_qual[1]), 
	.D(pprow5[1]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[1]  (.Q(pprow1_qual[1]), 
	.D(pprow1[1]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[6]  (.Q(pprow1_qual[6]), 
	.D(pprow1[6]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow3_qual_reg[4]  (.Q(pprow3_qual[4]), 
	.D(pprow3[4]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[5]  (.Q(pprow1_qual[5]), 
	.D(pprow1[5]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow1_qual_reg[7]  (.Q(pprow1_qual[7]), 
	.D(pprow1[7]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[25]  (.Q(pprow2_qual[25]), 
	.D(pprow2[25]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[23]  (.Q(pprow3_qual[23]), 
	.D(pprow3[23]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[17]  (.Q(pprow6_qual[17]), 
	.D(pprow6[17]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[11]  (.Q(pprow9_qual[11]), 
	.D(pprow9[11]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow12_qual_reg[5]  (.Q(pprow12_qual[5]), 
	.D(pprow12[5]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[31]  (.Q(pprow0_qual[31]), 
	.D(pprow0[31]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[21]  (.Q(pprow4_qual[21]), 
	.D(pprow4[21]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[15]  (.Q(pprow7_qual[15]), 
	.D(pprow7[15]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[9]  (.Q(pprow10_qual[9]), 
	.D(pprow10[9]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow13_qual_reg[3]  (.Q(pprow13_qual[3]), 
	.D(pprow13[3]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[29]  (.Q(pprow1_qual[29]), 
	.D(pprow1[29]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[19]  (.Q(pprow5_qual[19]), 
	.D(pprow5[19]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[13]  (.Q(pprow8_qual[13]), 
	.D(pprow8[13]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow11_qual_reg[7]  (.Q(pprow11_qual[7]), 
	.D(pprow11[7]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow14_qual_reg[1]  (.Q(pprow14_qual[1]), 
	.D(pprow14[1]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[20]  (.Q(pprow4_qual[20]), 
	.D(pprow4[20]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[28]  (.Q(pprow0_qual[28]), 
	.D(pprow0[28]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[26]  (.Q(pprow0_qual[26]), 
	.D(pprow0[26]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[20]  (.Q(pprow3_qual[20]), 
	.D(pprow3[20]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[18]  (.Q(pprow3_qual[18]), 
	.D(pprow3[18]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[16]  (.Q(pprow3_qual[16]), 
	.D(pprow3[16]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[11]  (.Q(pprow3_qual[11]), 
	.D(pprow3[11]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[17]  (.Q(pprow5_qual[17]), 
	.D(pprow5[17]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[14]  (.Q(pprow5_qual[14]), 
	.D(pprow5[14]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[13]  (.Q(pprow5_qual[13]), 
	.D(pprow5[13]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow12_qual_reg[1]  (.Q(pprow12_qual[1]), 
	.D(pprow12[1]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[30]  (.Q(pprow0_qual[30]), 
	.D(pprow0[30]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[29]  (.Q(pprow0_qual[29]), 
	.D(pprow0[29]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[22]  (.Q(pprow2_qual[22]), 
	.D(pprow2[22]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[20]  (.Q(pprow2_qual[20]), 
	.D(pprow2[20]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[18]  (.Q(pprow2_qual[18]), 
	.D(pprow2[18]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[13]  (.Q(pprow2_qual[13]), 
	.D(pprow2[13]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[19]  (.Q(pprow4_qual[19]), 
	.D(pprow4[19]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[16]  (.Q(pprow4_qual[16]), 
	.D(pprow4[16]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[15]  (.Q(pprow4_qual[15]), 
	.D(pprow4[15]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow12_qual_reg[0]  (.Q(pprow12_qual[0]), 
	.D(pprow12[0]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow14_qual_reg[0]  (.Q(pprow14_qual[0]), 
	.D(pprow14[0]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[18]  (.Q(pprow5_qual[18]), 
	.D(pprow5[18]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[21]  (.Q(pprow3_qual[21]), 
	.D(pprow3[21]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[23]  (.Q(pprow2_qual[23]), 
	.D(pprow2[23]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[24]  (.Q(pprow0_qual[24]), 
	.D(pprow0[24]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[27]  (.Q(pprow0_qual[27]), 
	.D(pprow0[27]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[25]  (.Q(pprow0_qual[25]), 
	.D(pprow0[25]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[24]  (.Q(pprow2_qual[24]), 
	.D(pprow2[24]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[17]  (.Q(pprow2_qual[17]), 
	.D(pprow2[17]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[16]  (.Q(pprow2_qual[16]), 
	.D(pprow2[16]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[14]  (.Q(pprow2_qual[14]), 
	.D(pprow2[14]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[16]  (.Q(pprow6_qual[16]), 
	.D(pprow6[16]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[7]  (.Q(pprow8_qual[7]), 
	.D(pprow8[7]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow12_qual_reg[2]  (.Q(pprow12_qual[2]), 
	.D(pprow12[2]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[18]  (.Q(pprow4_qual[18]), 
	.D(pprow4[18]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[14]  (.Q(pprow6_qual[14]), 
	.D(pprow6[14]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[12]  (.Q(pprow6_qual[12]), 
	.D(pprow6[12]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[9]  (.Q(pprow8_qual[9]), 
	.D(pprow8[9]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[6]  (.Q(pprow10_qual[6]), 
	.D(pprow10[6]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow11_qual_reg[6]  (.Q(pprow11_qual[6]), 
	.D(pprow11[6]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[19]  (.Q(pprow2_qual[19]), 
	.D(pprow2[19]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[22]  (.Q(pprow3_qual[22]), 
	.D(pprow3[22]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[15]  (.Q(pprow3_qual[15]), 
	.D(pprow3[15]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[14]  (.Q(pprow3_qual[14]), 
	.D(pprow3[14]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[12]  (.Q(pprow3_qual[12]), 
	.D(pprow3[12]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[14]  (.Q(pprow7_qual[14]), 
	.D(pprow7[14]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[5]  (.Q(pprow9_qual[5]), 
	.D(pprow9[5]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow13_qual_reg[0]  (.Q(pprow13_qual[0]), 
	.D(pprow13[0]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[11]  (.Q(pprow5_qual[11]), 
	.D(pprow5[11]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[10]  (.Q(pprow5_qual[10]), 
	.D(pprow5[10]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[6]  (.Q(pprow7_qual[6]), 
	.D(pprow7[6]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[3]  (.Q(pprow9_qual[3]), 
	.D(pprow9[3]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[10]  (.Q(pprow9_qual[10]), 
	.D(pprow9[10]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow13_qual_reg[2]  (.Q(pprow13_qual[2]), 
	.D(pprow13[2]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[28]  (.Q(pprow1_qual[28]), 
	.D(pprow1[28]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[8]  (.Q(pprow10_qual[8]), 
	.D(pprow10[8]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[13]  (.Q(pprow4_qual[13]), 
	.D(pprow4[13]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[12]  (.Q(pprow4_qual[12]), 
	.D(pprow4[12]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[8]  (.Q(pprow6_qual[8]), 
	.D(pprow6[8]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[5]  (.Q(pprow8_qual[5]), 
	.D(pprow8[5]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[16]  (.Q(pprow5_qual[16]), 
	.D(pprow5[16]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[12]  (.Q(pprow7_qual[12]), 
	.D(pprow7[12]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[10]  (.Q(pprow7_qual[10]), 
	.D(pprow7[10]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[7]  (.Q(pprow9_qual[7]), 
	.D(pprow9[7]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow11_qual_reg[4]  (.Q(pprow11_qual[4]), 
	.D(pprow11[4]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[9]  (.Q(pprow9_qual[9]), 
	.D(pprow9[9]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[19]  (.Q(pprow3_qual[19]), 
	.D(pprow3[19]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[21]  (.Q(pprow2_qual[21]), 
	.D(pprow2[21]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[12]  (.Q(pprow8_qual[12]), 
	.D(pprow8[12]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow12_qual_reg[4]  (.Q(pprow12_qual[4]), 
	.D(pprow12[4]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[10]  (.Q(pprow6_qual[10]), 
	.D(pprow6[10]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[11]  (.Q(pprow8_qual[11]), 
	.D(pprow8[11]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[7]  (.Q(pprow10_qual[7]), 
	.D(pprow10[7]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow12_qual_reg[3]  (.Q(pprow12_qual[3]), 
	.D(pprow12[3]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[8]  (.Q(pprow7_qual[8]), 
	.D(pprow7[8]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[17]  (.Q(pprow3_qual[17]), 
	.D(pprow3[17]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[10]  (.Q(pprow8_qual[10]), 
	.D(pprow8[10]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[8]  (.Q(pprow8_qual[8]), 
	.D(pprow8[8]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[6]  (.Q(pprow8_qual[6]), 
	.D(pprow8[6]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow11_qual_reg[5]  (.Q(pprow11_qual[5]), 
	.D(pprow11[5]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow13_qual_reg[1]  (.Q(pprow13_qual[1]), 
	.D(pprow13[1]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[17]  (.Q(pprow4_qual[17]), 
	.D(pprow4[17]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[14]  (.Q(pprow4_qual[14]), 
	.D(pprow4[14]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[23]  (.Q(pprow0_qual[23]), 
	.D(pprow0[23]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[13]  (.Q(pprow6_qual[13]), 
	.D(pprow6[13]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[27]  (.Q(pprow1_qual[27]), 
	.D(pprow1[27]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[8]  (.Q(pprow9_qual[8]), 
	.D(pprow9[8]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[6]  (.Q(pprow9_qual[6]), 
	.D(pprow9[6]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[4]  (.Q(pprow9_qual[4]), 
	.D(pprow9[4]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[15]  (.Q(pprow5_qual[15]), 
	.D(pprow5[15]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[12]  (.Q(pprow5_qual[12]), 
	.D(pprow5[12]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow2_qual_reg[15]  (.Q(pprow2_qual[15]), 
	.D(pprow2[15]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[11]  (.Q(pprow7_qual[11]), 
	.D(pprow7[11]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[13]  (.Q(pprow3_qual[13]), 
	.D(pprow3[13]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[15]  (.Q(pprow6_qual[15]), 
	.D(pprow6[15]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[11]  (.Q(pprow6_qual[11]), 
	.D(pprow6[11]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[26]  (.Q(pprow1_qual[26]), 
	.D(pprow1[26]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[13]  (.Q(pprow7_qual[13]), 
	.D(pprow7[13]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[9]  (.Q(pprow7_qual[9]), 
	.D(pprow7[9]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[24]  (.Q(pprow1_qual[24]), 
	.D(pprow1[24]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[23]  (.Q(pprow1_qual[23]), 
	.D(pprow1[23]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[22]  (.Q(pprow1_qual[22]), 
	.D(pprow1[22]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[21]  (.Q(pprow1_qual[21]), 
	.D(pprow1[21]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[20]  (.Q(pprow1_qual[20]), 
	.D(pprow1[20]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[25]  (.Q(pprow1_qual[25]), 
	.D(pprow1[25]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[7]  (.Q(pprow2_qual[7]), 
	.D(pprow2[7]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[5]  (.Q(pprow6_qual[5]), 
	.D(pprow6[5]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[2]  (.Q(pprow8_qual[2]), 
	.D(pprow8[2]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[1]  (.Q(pprow8_qual[1]), 
	.D(pprow8[1]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[2]  (.Q(pprow10_qual[2]), 
	.D(pprow10[2]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[0]  (.Q(pprow9_qual[0]), 
	.D(pprow9[0]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow11_qual_reg[1]  (.Q(pprow11_qual[1]), 
	.D(pprow11[1]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[18]  (.Q(pprow1_qual[18]), 
	.D(pprow1[18]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow5_qual_reg[2]  (.Q(pprow5_qual[2]), 
	.D(pprow5[2]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow4_qual_reg[4]  (.Q(pprow4_qual[4]), 
	.D(pprow4[4]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[2]  (.Q(pprow2_qual[2]), 
	.D(pprow2[2]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow3_qual_reg[6]  (.Q(pprow3_qual[6]), 
	.D(pprow3[6]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[1]  (.Q(pprow2_qual[1]), 
	.D(pprow2[1]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow7_qual_reg[1]  (.Q(pprow7_qual[1]), 
	.D(pprow7[1]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow6_qual_reg[3]  (.Q(pprow6_qual[3]), 
	.D(pprow6[3]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow4_qual_reg[5]  (.Q(pprow4_qual[5]), 
	.D(pprow4[5]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[0]  (.Q(pprow2_qual[0]), 
	.D(pprow2[0]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow6_qual_reg[1]  (.Q(pprow6_qual[1]), 
	.D(pprow6[1]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow3_qual_reg[7]  (.Q(pprow3_qual[7]), 
	.D(pprow3[7]), 
	.CK(CLK));
   SEN_FDPQ_D_2 \pprow3_qual_reg[9]  (.Q(pprow3_qual[9]), 
	.D(pprow3[9]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow11_qual_reg[0]  (.Q(pprow11_qual[0]), 
	.D(pprow11[0]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow0_qual_reg[8]  (.Q(pprow0_qual[8]), 
	.D(pprow0[8]), 
	.CK(CLK));
   SEN_ND2_4 net101362 (.X(net84063), 
	.A2(net84073), 
	.A1(n128));
   SEN_FDPQ_D_4 \pprow0_qual_reg[1]  (.Q(pprow0_qual[1]), 
	.D(pprow0[1]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow1_qual_reg[14]  (.Q(pprow1_qual[14]), 
	.D(pprow1[14]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow4_qual_reg[7]  (.Q(pprow4_qual[7]), 
	.D(pprow4[7]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow4_qual_reg[2]  (.Q(pprow4_qual[2]), 
	.D(pprow4[2]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow4_qual_reg[1]  (.Q(pprow4_qual[1]), 
	.D(pprow4[1]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[20]  (.Q(pprow0_qual[20]), 
	.D(pprow0[20]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[21]  (.Q(pprow0_qual[21]), 
	.D(pprow0[21]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[17]  (.Q(pprow0_qual[17]), 
	.D(pprow0[17]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow0_qual_reg[16]  (.Q(pprow0_qual[16]), 
	.D(pprow0[16]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[19]  (.Q(pprow0_qual[19]), 
	.D(pprow0[19]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[4]  (.Q(pprow10_qual[4]), 
	.D(pprow10[4]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[10]  (.Q(pprow4_qual[10]), 
	.D(pprow4[10]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[9]  (.Q(pprow6_qual[9]), 
	.D(pprow6[9]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[15]  (.Q(pprow0_qual[15]), 
	.D(pprow0[15]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[3]  (.Q(pprow10_qual[3]), 
	.D(pprow10[3]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[6]  (.Q(pprow6_qual[6]), 
	.D(pprow6[6]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[8]  (.Q(pprow5_qual[8]), 
	.D(pprow5[8]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[7]  (.Q(pprow7_qual[7]), 
	.D(pprow7[7]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow11_qual_reg[2]  (.Q(pprow11_qual[2]), 
	.D(pprow11[2]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[5]  (.Q(pprow10_qual[5]), 
	.D(pprow10[5]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[4]  (.Q(pprow7_qual[4]), 
	.D(pprow7[4]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[3]  (.Q(pprow8_qual[3]), 
	.D(pprow8[3]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow11_qual_reg[3]  (.Q(pprow11_qual[3]), 
	.D(pprow11[3]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[1]  (.Q(pprow9_qual[1]), 
	.D(pprow9[1]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow8_qual_reg[4]  (.Q(pprow8_qual[4]), 
	.D(pprow8[4]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow6_qual_reg[7]  (.Q(pprow6_qual[7]), 
	.D(pprow6[7]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow4_qual_reg[11]  (.Q(pprow4_qual[11]), 
	.D(pprow4[11]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow9_qual_reg[2]  (.Q(pprow9_qual[2]), 
	.D(pprow9[2]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[5]  (.Q(pprow7_qual[5]), 
	.D(pprow7[5]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow5_qual_reg[9]  (.Q(pprow5_qual[9]), 
	.D(pprow5[9]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow3_qual_reg[10]  (.Q(pprow3_qual[10]), 
	.D(pprow3[10]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow1_qual_reg[19]  (.Q(pprow1_qual[19]), 
	.D(pprow1[19]), 
	.CK(CLK));
   SEN_FDPQ_D_2 \pprow2_qual_reg[12]  (.Q(pprow2_qual[12]), 
	.D(pprow2[12]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[22]  (.Q(pprow0_qual[22]), 
	.D(pprow0[22]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[0]  (.Q(pprow10_qual[0]), 
	.D(pprow10[0]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow10_qual_reg[1]  (.Q(pprow10_qual[1]), 
	.D(pprow10[1]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow0_qual_reg[0]  (.Q(pprow0_qual[0]), 
	.D(pprow0[0]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow0_qual_reg[5]  (.Q(pprow0_qual[5]), 
	.D(pprow0[5]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow5_qual_reg[6]  (.Q(pprow5_qual[6]), 
	.D(pprow5[6]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow2_qual_reg[8]  (.Q(pprow2_qual[8]), 
	.D(pprow2[8]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow0_qual_reg[4]  (.Q(pprow0_qual[4]), 
	.D(pprow0[4]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow1_qual_reg[17]  (.Q(pprow1_qual[17]), 
	.D(pprow1[17]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[12]  (.Q(pprow0_qual[12]), 
	.D(pprow0[12]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow4_qual_reg[0]  (.Q(pprow4_qual[0]), 
	.D(pprow4[0]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow7_qual_reg[3]  (.Q(pprow7_qual[3]), 
	.D(pprow7[3]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[14]  (.Q(pprow0_qual[14]), 
	.D(pprow0[14]), 
	.CK(CLK));
   SEN_FDPQ_D_2 \pprow0_qual_reg[11]  (.Q(pprow0_qual[11]), 
	.D(pprow0[11]), 
	.CK(CLK));
   SEN_FDPQ_D_2 \pprow0_qual_reg[9]  (.Q(pprow0_qual[9]), 
	.D(pprow0[9]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow2_qual_reg[10]  (.Q(pprow2_qual[10]), 
	.D(pprow2[10]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[18]  (.Q(pprow0_qual[18]), 
	.D(pprow0[18]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[13]  (.Q(pprow0_qual[13]), 
	.D(pprow0[13]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow2_qual_reg[9]  (.Q(pprow2_qual[9]), 
	.D(pprow2[9]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow5_qual_reg[7]  (.Q(pprow5_qual[7]), 
	.D(pprow5[7]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow4_qual_reg[9]  (.Q(pprow4_qual[9]), 
	.D(pprow4[9]), 
	.CK(CLK));
   SEN_FDPQ_D_2 \pprow7_qual_reg[2]  (.Q(pprow7_qual[2]), 
	.D(pprow7[2]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow3_qual_reg[8]  (.Q(pprow3_qual[8]), 
	.D(pprow3[8]), 
	.CK(CLK));
   SEN_FDPQ_D_1 \pprow0_qual_reg[6]  (.Q(pprow0_qual[6]), 
	.D(pprow0[6]), 
	.CK(CLK));
   SEN_FDPQ_D_2 \pprow0_qual_reg[10]  (.Q(pprow0_qual[10]), 
	.D(pprow0[10]), 
	.CK(CLK));
   SEN_FDPQ_D_2 \pprow8_qual_reg[0]  (.Q(pprow8_qual[0]), 
	.D(pprow8[0]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow6_qual_reg[4]  (.Q(pprow6_qual[4]), 
	.D(pprow6[4]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow0_qual_reg[7]  (.Q(pprow0_qual[7]), 
	.D(pprow0[7]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow1_qual_reg[16]  (.Q(pprow1_qual[16]), 
	.D(pprow1[16]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow5_qual_reg[4]  (.Q(pprow5_qual[4]), 
	.D(pprow5[4]), 
	.CK(CLK));
   SEN_FDPQ_2 \pprow4_qual_reg[8]  (.Q(pprow4_qual[8]), 
	.D(pprow4[8]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow4_qual_reg[6]  (.Q(pprow4_qual[6]), 
	.D(pprow4[6]), 
	.CK(CLK));
   SEN_FDPQ_1 \pprow0_qual_reg[3]  (.Q(pprow0_qual[3]), 
	.D(pprow0[3]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow4_qual_reg[3]  (.Q(pprow4_qual[3]), 
	.D(pprow4[3]), 
	.CK(CLK));
   SEN_ND2B_1 U23 (.X(net82819), 
	.B(net102677), 
	.A(net82634));
   SEN_ND2_G_3 U24 (.X(n1578), 
	.A2(n1526), 
	.A1(n1527));
   SEN_ND2_T_5 U25 (.X(net84196), 
	.A2(net84221), 
	.A1(net90868));
   SEN_ND2_1P5 U26 (.X(n1030), 
	.A2(pprow4_qual[0]), 
	.A1(n810));
   SEN_OAI21_S_1 U27 (.X(n1139), 
	.B(n1175), 
	.A2(n1180), 
	.A1(n810));
   SEN_INV_4 U28 (.X(n511), 
	.A(net84208));
   SEN_OR2_2 U29 (.X(n705), 
	.A2(n267), 
	.A1(n1523));
   SEN_EN2_S_4 U31 (.X(n1738), 
	.A2(n1736), 
	.A1(n1737));
   SEN_NR2_6 U33 (.X(n18), 
	.A2(n1603), 
	.A1(n1604));
   SEN_NR2_G_4 U35 (.X(n1098), 
	.A2(net83552), 
	.A1(n2045));
   SEN_INV_2P5 U38 (.X(n899), 
	.A(n901));
   SEN_EO2_S_3 U39 (.X(n901), 
	.A2(n730), 
	.A1(n729));
   SEN_INV_4 U41 (.X(net88078), 
	.A(net82429));
   SEN_BUF_1 U42 (.X(n19), 
	.A(net82522));
   SEN_INV_S_1 U43 (.X(n20), 
	.A(n1781));
   SEN_EN2_1 U44 (.X(n1777), 
	.A2(n1785), 
	.A1(n719));
   SEN_INV_2 U45 (.X(n540), 
	.A(n897));
   SEN_NR2B_2 U46 (.X(n894), 
	.B(n893), 
	.A(n897));
   SEN_ND2_T_1 U47 (.X(net82210), 
	.A2(n1735), 
	.A1(n1734));
   SEN_INV_1 U48 (.X(n274), 
	.A(n285));
   SEN_EO2_S_6 U50 (.X(n701), 
	.A2(n31), 
	.A1(net82091));
   SEN_AO21_DG_4 U52 (.X(n21), 
	.B(n1544), 
	.A2(pprow0_qual[24]), 
	.A1(C[24]));
   SEN_ND2B_S_4 U53 (.X(n1619), 
	.B(n1572), 
	.A(n1574));
   SEN_ND2_T_2 U54 (.X(n1621), 
	.A2(n1573), 
	.A1(n1574));
   SEN_OAI21_5 U55 (.X(net82057), 
	.B(net82245), 
	.A2(net82244), 
	.A1(net82243));
   SEN_EO2_S_6 U56 (.X(net82334), 
	.A2(net82243), 
	.A1(net90631));
   SEN_BUF_D_3 U57 (.X(net91564), 
	.A(net82280));
   SEN_ND2_0P8 U58 (.X(n776), 
	.A2(n1741), 
	.A1(n1742));
   SEN_OAI21_G_6 U59 (.X(n1445), 
	.B(n1441), 
	.A2(net82962), 
	.A1(n1442));
   SEN_ND2_T_8 U61 (.X(net83609), 
	.A2(n1185), 
	.A1(n1186));
   SEN_INV_S_8 U62 (.X(n1802), 
	.A(n1730));
   SEN_NR2_G_3 U63 (.X(n1715), 
	.A2(n81), 
	.A1(n1710));
   SEN_INV_1 U64 (.X(n81), 
	.A(n384));
   SEN_INV_S_3 U65 (.X(n1710), 
	.A(n1767));
   SEN_EO2_4 U68 (.X(n1020), 
	.A2(net84106), 
	.A1(n993));
   SEN_AN3B_4 U69 (.X(net84106), 
	.B2(net84029), 
	.B1(net83741), 
	.A(n49));
   SEN_ND2_T_8 U71 (.X(net82936), 
	.A2(net91120), 
	.A1(net83153));
   SEN_ND4_2 U73 (.X(n22), 
	.A4(net83385), 
	.A3(net85046), 
	.A2(net83172), 
	.A1(n45));
   SEN_ND4_1 U74 (.X(net83204), 
	.A4(net83385), 
	.A3(net85046), 
	.A2(net83172), 
	.A1(n45));
   SEN_INV_1 U76 (.X(n1749), 
	.A(n1745));
   SEN_ND2_G_1 U77 (.X(n1747), 
	.A2(n1745), 
	.A1(n1746));
   SEN_EN2_S_2 U78 (.X(n1745), 
	.A2(n1756), 
	.A1(n1695));
   SEN_INV_S_0P5 U79 (.X(n23), 
	.A(net88078));
   SEN_BUF_4 U80 (.X(n204), 
	.A(n566));
   SEN_NR2_T_3 U81 (.X(n1494), 
	.A2(n1492), 
	.A1(n1493));
   SEN_ND2_2 U82 (.X(net82235), 
	.A2(net82237), 
	.A1(net82236));
   SEN_EO2_3 U83 (.X(net82236), 
	.A2(n739), 
	.A1(n1793));
   SEN_EO2_2 U84 (.X(n24), 
	.A2(n1028), 
	.A1(n1027));
   SEN_EO2_S_3 U85 (.X(net83918), 
	.A2(n1028), 
	.A1(n1027));
   SEN_ND2_2 U86 (.X(n1028), 
	.A2(n1065), 
	.A1(n1106));
   SEN_ND2B_V1_8 U87 (.X(net84186), 
	.B(n900), 
	.A(n899));
   SEN_ND2B_6 U88 (.X(n25), 
	.B(net83540), 
	.A(net83541));
   SEN_ND2B_4 U89 (.X(net83297), 
	.B(net83540), 
	.A(net83541));
   SEN_EO2_4 U90 (.X(net83541), 
	.A2(net86023), 
	.A1(net86022));
   SEN_ND2_S_8 U91 (.X(n283), 
	.A2(net91110), 
	.A1(net85837));
   SEN_INV_3 U93 (.X(n67), 
	.A(net86273));
   SEN_AOI21B_4 U95 (.X(n1348), 
	.B(n1379), 
	.A2(n604), 
	.A1(n1345));
   SEN_INV_5 U97 (.X(net83961), 
	.A(net84650));
   SEN_EN2_S_2 U98 (.X(n1045), 
	.A2(n1043), 
	.A1(n1044));
   SEN_NR2B_V1DG_2 U99 (.X(net86390), 
	.B(n987), 
	.A(n985));
   SEN_ND2_2 U100 (.X(net86266), 
	.A2(net90740), 
	.A1(n358));
   SEN_BUF_1 U101 (.X(n26), 
	.A(net83632));
   SEN_ND2B_S_4 U103 (.X(n639), 
	.B(net83689), 
	.A(n638));
   SEN_INV_1P25 U104 (.X(net88089), 
	.A(n457));
   SEN_INV_S_2 U105 (.X(n471), 
	.A(net83333));
   SEN_AN2_4 U107 (.X(net87795), 
	.A2(n25), 
	.A1(n480));
   SEN_ND2_T_6 U108 (.X(net84372), 
	.A2(n881), 
	.A1(n882));
   SEN_OAI21_G_2 U109 (.X(n1249), 
	.B(n557), 
	.A2(n1273), 
	.A1(n669));
   SEN_ND2_3 U110 (.X(net87351), 
	.A2(n214), 
	.A1(net83111));
   SEN_EO2_3 U112 (.X(n867), 
	.A2(net86699), 
	.A1(n458));
   SEN_EO2_DG_1 U113 (.X(n458), 
	.A2(n524), 
	.A1(n872));
   SEN_INV_1P5 U114 (.X(n1085), 
	.A(n1138));
   SEN_INV_1 U115 (.X(net83989), 
	.A(net83952));
   SEN_EN2_S_6 U116 (.X(n992), 
	.A2(n544), 
	.A1(n27));
   SEN_EO2_DG_8 U117 (.X(n27), 
	.A2(n48), 
	.A1(net84117));
   SEN_OAI21_4 U118 (.X(net82742), 
	.B(net83072), 
	.A2(net83071), 
	.A1(net83070));
   SEN_BUF_D_1 U119 (.X(n515), 
	.A(n1476));
   SEN_AO21B_8 U120 (.X(n1476), 
	.B(n1411), 
	.A2(n748), 
	.A1(n1410));
   SEN_ND2_T_2 U123 (.X(n878), 
	.A2(pprow0_qual[4]), 
	.A1(C[4]));
   SEN_EO2_6 U124 (.X(net83505), 
	.A2(n29), 
	.A1(n28));
   SEN_EN2_DG_8 U125 (.X(n28), 
	.A2(C[17]), 
	.A1(net83516));
   SEN_AO31_4 U126 (.X(n29), 
	.B(net83526), 
	.A3(net83522), 
	.A2(net101269), 
	.A1(net83639));
   SEN_INV_6 U127 (.X(n57), 
	.A(n56));
   SEN_BUF_1 U128 (.X(net101248), 
	.A(n56));
   SEN_ND2_T_4 U129 (.X(net83333), 
	.A2(net83455), 
	.A1(net83454));
   SEN_ND2_G_4 U130 (.X(n1759), 
	.A2(net88113), 
	.A1(n571));
   SEN_INV_1P5 U132 (.X(n1742), 
	.A(n1740));
   SEN_EN2_2 U133 (.X(net83076), 
	.A2(net98319), 
	.A1(net83090));
   SEN_NR2_T_0P5 U134 (.X(n331), 
	.A2(pprow1_qual[17]), 
	.A1(net83090));
   SEN_INV_S_6 U135 (.X(net98293), 
	.A(net83090));
   SEN_BUF_2 U136 (.X(n30), 
	.A(net83993));
   SEN_ND2_4 U137 (.X(net83952), 
	.A2(net83991), 
	.A1(n1035));
   SEN_NR2_2 U138 (.X(n193), 
	.A2(net87549), 
	.A1(net84650));
   SEN_ND2_6 U140 (.X(net84007), 
	.A2(n940), 
	.A1(n941));
   SEN_ND2_T_2 U141 (.X(net84157), 
	.A2(pprow0_qual[8]), 
	.A1(C[8]));
   SEN_ND2B_V1_2 U142 (.X(net84153), 
	.B(net84288), 
	.A(C[8]));
   SEN_ND2_T_1 U143 (.X(n88), 
	.A2(pprow0_qual[7]), 
	.A1(C[8]));
   SEN_NR2_T_2 U144 (.X(net84417), 
	.A2(net84394), 
	.A1(net84451));
   SEN_NR2_T_1P5 U145 (.X(net84451), 
	.A2(pprow0_qual[1]), 
	.A1(net84734));
   SEN_OA21_2 U146 (.X(n45), 
	.B(n55), 
	.A2(net83389), 
	.A1(net83390));
   SEN_BUF_S_6 U147 (.X(n249), 
	.A(net84228));
   SEN_ND2B_V1_3 U148 (.X(n265), 
	.B(net83614), 
	.A(net83611));
   SEN_INV_6 U149 (.X(n1084), 
	.A(n1173));
   SEN_NR2_S_1 U150 (.X(net83998), 
	.A2(net84011), 
	.A1(net83580));
   SEN_INV_S_2 U151 (.X(net84011), 
	.A(net83965));
   SEN_OAOI211_1 U153 (.X(n562), 
	.C(n1375), 
	.B(n386), 
	.A2(n1377), 
	.A1(n1378));
   SEN_INV_S_2 U154 (.X(net83105), 
	.A(net83097));
   SEN_ND2_4 U156 (.X(net83103), 
	.A2(n1351), 
	.A1(n1352));
   SEN_ND2_T_4 U157 (.X(net82586), 
	.A2(n1588), 
	.A1(n1587));
   SEN_AOI21_T_1 U159 (.X(n1555), 
	.B(net82820), 
	.A2(net82819), 
	.A1(net82638));
   SEN_OAOI211_G_4 U160 (.X(n32), 
	.C(n1607), 
	.B(n1608), 
	.A2(pprow8_qual[8]), 
	.A1(pprow9_qual[6]));
   SEN_BUF_1 U161 (.X(n33), 
	.A(n1033));
   SEN_EO2_DG_1 U162 (.X(n675), 
	.A2(n1163), 
	.A1(n236));
   SEN_ND2_S_3 U163 (.X(n1439), 
	.A2(n1163), 
	.A1(n236));
   SEN_ND2B_V1_2 U164 (.X(n1334), 
	.B(n1301), 
	.A(pprow6_qual[5]));
   SEN_INV_6 U165 (.X(n1184), 
	.A(n1188));
   SEN_EO2_G_1 U167 (.X(n1117), 
	.A2(net83721), 
	.A1(n467));
   SEN_INV_S_4 U168 (.X(net83724), 
	.A(net83721));
   SEN_BUF_1 U171 (.X(n34), 
	.A(net82137));
   SEN_INV_S_0P5 U172 (.X(n35), 
	.A(n1779));
   SEN_INV_1P25 U175 (.X(net87762), 
	.A(net82936));
   SEN_ND2_4 U176 (.X(n1131), 
	.A2(net83685), 
	.A1(n629));
   SEN_INV_8 U177 (.X(net84273), 
	.A(net84274));
   SEN_INV_2P5 U178 (.X(n592), 
	.A(n1118));
   SEN_OAI21_G_2 U180 (.X(net83538), 
	.B(n25), 
	.A2(n487), 
	.A1(n480));
   SEN_ND2_S_6 U181 (.X(n1309), 
	.A2(n1173), 
	.A1(n1179));
   SEN_ND3_T_6 U182 (.X(n1173), 
	.A3(n1051), 
	.A2(n1049), 
	.A1(n1050));
   SEN_ND2_4 U183 (.X(net84004), 
	.A2(net84002), 
	.A1(net84008));
   SEN_ND3_T_4 U184 (.X(n318), 
	.A3(net83814), 
	.A2(net83815), 
	.A1(net83816));
   SEN_ND2_T_6 U186 (.X(n1725), 
	.A2(n586), 
	.A1(n1722));
   SEN_ND2_G_3 U187 (.X(net83376), 
	.A2(n958), 
	.A1(n959));
   SEN_ND3_T_2 U188 (.X(n295), 
	.A3(n296), 
	.A2(net83852), 
	.A1(n301));
   SEN_INV_S_4 U189 (.X(n296), 
	.A(net83376));
   SEN_ND2_T_6 U190 (.X(net84040), 
	.A2(n296), 
	.A1(net87828));
   SEN_AOI31_T_2 U191 (.X(n948), 
	.B(n947), 
	.A3(net84218), 
	.A2(n959), 
	.A1(net97377));
   SEN_INV_4 U193 (.X(n399), 
	.A(n1842));
   SEN_ND2_S_2 U194 (.X(n211), 
	.A2(n1173), 
	.A1(n1179));
   SEN_BUF_2 U195 (.X(n38), 
	.A(n1179));
   SEN_AOI21B_4 U197 (.X(net84081), 
	.B(net84042), 
	.A2(n301), 
	.A1(net84121));
   SEN_ND2_S_4 U198 (.X(net84121), 
	.A2(net84040), 
	.A1(n80));
   SEN_EO2_DG_1 U200 (.X(net86002), 
	.A2(net84361), 
	.A1(C[6]));
   SEN_INV_4 U201 (.X(n36), 
	.A(net83778));
   SEN_INV_S_6 U202 (.X(net83778), 
	.A(net83584));
   SEN_INV_S_6 U204 (.X(net86274), 
	.A(n199));
   SEN_EN2_8 U205 (.X(net83389), 
	.A2(net86655), 
	.A1(n37));
   SEN_EO2_DG_8 U206 (.X(n37), 
	.A2(C[19]), 
	.A1(n1289));
   SEN_EO2_1 U207 (.X(net83451), 
	.A2(net83334), 
	.A1(net87796));
   SEN_ND2_T_6 U209 (.X(net83555), 
	.A2(n1096), 
	.A1(n1097));
   SEN_INV_6 U211 (.X(net83387), 
	.A(net83370));
   SEN_EO2_5 U212 (.X(net83415), 
	.A2(n210), 
	.A1(n695));
   SEN_OAI21_T_4 U213 (.X(n1344), 
	.B(n1319), 
	.A2(n1320), 
	.A1(n1321));
   SEN_ND2_G_1 U214 (.X(n1666), 
	.A2(net82426), 
	.A1(net82431));
   SEN_BUF_AS_3 U215 (.X(n557), 
	.A(n1274));
   SEN_EN2_8 U216 (.X(net82241), 
	.A2(net82058), 
	.A1(net82056));
   SEN_ND2_T_2 U217 (.X(n1106), 
	.A2(n1019), 
	.A1(n1020));
   SEN_INV_6 U218 (.X(n1021), 
	.A(n1020));
   SEN_EN2_DG_1 U219 (.X(net83627), 
	.A2(net83506), 
	.A1(net83505));
   SEN_ND2_2 U222 (.X(n444), 
	.A2(net84284), 
	.A1(net84228));
   SEN_OAOI211_8 U223 (.X(n1756), 
	.C(n1693), 
	.B(n1694), 
	.A2(pprow10_qual[5]), 
	.A1(pprow11_qual[3]));
   SEN_INV_S_6 U224 (.X(net84358), 
	.A(net84359));
   SEN_BUF_S_4 U225 (.X(n39), 
	.A(net83165));
   SEN_ND2_G_4 U226 (.X(n1082), 
	.A2(pprow5_qual[1]), 
	.A1(pprow4_qual[3]));
   SEN_OAI21_8 U227 (.X(n1308), 
	.B(n1082), 
	.A2(n1083), 
	.A1(n1052));
   SEN_ND2_T_3 U229 (.X(n473), 
	.A2(net94064), 
	.A1(n477));
   SEN_NR2_G_4 U230 (.X(net84229), 
	.A2(net84235), 
	.A1(n945));
   SEN_EO2_0P5 U233 (.X(net86306), 
	.A2(n26), 
	.A1(net83634));
   SEN_ND2_3 U234 (.X(n196), 
	.A2(net84001), 
	.A1(n193));
   SEN_ND2_T_6 U236 (.X(net94064), 
	.A2(n241), 
	.A1(net83609));
   SEN_ND2B_V1_6 U237 (.X(net82238), 
	.B(n1725), 
	.A(n547));
   SEN_ND2_S_6 U239 (.X(n384), 
	.A2(n1660), 
	.A1(n661));
   SEN_EO2_8 U240 (.X(net86498), 
	.A2(net82305), 
	.A1(net82304));
   SEN_AOI21_S_4 U241 (.X(net84353), 
	.B(net84356), 
	.A2(net84355), 
	.A1(net84354));
   SEN_ND2_T_1 U244 (.X(n1011), 
	.A2(n1050), 
	.A1(n810));
   SEN_INV_1 U245 (.X(net83224), 
	.A(net83220));
   SEN_EN2_DG_4 U246 (.X(n205), 
	.A2(net91065), 
	.A1(net83220));
   SEN_ND2_T_2 U247 (.X(n1379), 
	.A2(net83224), 
	.A1(net83223));
   SEN_ND2_T_2 U248 (.X(n600), 
	.A2(n604), 
	.A1(net83127));
   SEN_ND2_2 U249 (.X(n1483), 
	.A2(n1386), 
	.A1(n1387));
   SEN_INV_6 U250 (.X(net95563), 
	.A(net95575));
   SEN_ND2_S_4 U251 (.X(n506), 
	.A2(net84068), 
	.A1(net84067));
   SEN_INV_S_4 U252 (.X(n320), 
	.A(n319));
   SEN_ND2_T_4 U253 (.X(n319), 
	.A2(net83813), 
	.A1(n317));
   SEN_ND2_T_5 U254 (.X(net83813), 
	.A2(net84046), 
	.A1(net84047));
   SEN_ND2_T_8 U256 (.X(net83418), 
	.A2(net83508), 
	.A1(net83507));
   SEN_ND3_T_8 U257 (.X(net84443), 
	.A3(n277), 
	.A2(n276), 
	.A1(n275));
   SEN_ND2B_6 U258 (.X(n277), 
	.B(n283), 
	.A(n83));
   SEN_INV_1P25 U259 (.X(n271), 
	.A(net84734));
   SEN_NR2_T_4 U260 (.X(net87100), 
	.A2(n501), 
	.A1(n493));
   SEN_INV_6 U261 (.X(net83677), 
	.A(net83308));
   SEN_INV_3 U262 (.X(n78), 
	.A(net82309));
   SEN_ND2_T_6 U264 (.X(net86556), 
	.A2(n69), 
	.A1(net82742));
   SEN_INV_6 U265 (.X(net83843), 
	.A(net83845));
   SEN_EO2_3 U266 (.X(net86491), 
	.A2(n663), 
	.A1(n671));
   SEN_OAI21_T_3 U267 (.X(n1371), 
	.B(n1370), 
	.A2(pprow8_qual[3]), 
	.A1(pprow9_qual[1]));
   SEN_OAI21_5 U268 (.X(n1499), 
	.B(n1466), 
	.A2(n1467), 
	.A1(n1468));
   SEN_OAOI211_8 U269 (.X(n1468), 
	.C(n1400), 
	.B(n1401), 
	.A2(pprow8_qual[4]), 
	.A1(pprow9_qual[2]));
   SEN_OA2BB2_4 U270 (.X(net83825), 
	.B2(n114), 
	.B1(net83733), 
	.A2(net82999), 
	.A1(net83826));
   SEN_ND2_4 U271 (.X(n1241), 
	.A2(n552), 
	.A1(n703));
   SEN_AO21B_4 U272 (.X(n1388), 
	.B(n382), 
	.A2(n381), 
	.A1(n1344));
   SEN_INV_S_6 U273 (.X(n484), 
	.A(net83953));
   SEN_AOI22_T_1P5 U275 (.X(net82124), 
	.B2(pprow10_qual[8]), 
	.B1(pprow11_qual[6]), 
	.A2(n119), 
	.A1(net82125));
   SEN_ND2_T_2 U276 (.X(n1159), 
	.A2(n1157), 
	.A1(n1158));
   SEN_ND2B_V1_3 U277 (.X(n1157), 
	.B(net83936), 
	.A(C[13]));
   SEN_AOA211_DG_1 U278 (.X(n114), 
	.C(n1158), 
	.B(net83828), 
	.A2(n1157), 
	.A1(n1156));
   SEN_AN2_S_0P5 U279 (.X(net100921), 
	.A2(n1157), 
	.A1(n1156));
   SEN_INV_2 U281 (.X(net82997), 
	.A(net83001));
   SEN_INV_10 U282 (.X(net82336), 
	.A(net82334));
   SEN_AN2_6 U284 (.X(n1092), 
	.A2(n631), 
	.A1(net87791));
   SEN_ND3_T_6 U285 (.X(net82847), 
	.A3(n1453), 
	.A2(n1454), 
	.A1(n1455));
   SEN_ND3_T_3 U286 (.X(net87791), 
	.A3(net83887), 
	.A2(net83559), 
	.A1(net83885));
   SEN_INV_S_4 U288 (.X(net82824), 
	.A(net82822));
   SEN_AN2_S_1P5 U289 (.X(n577), 
	.A2(n1395), 
	.A1(net86332));
   SEN_INV_S_6 U290 (.X(n1179), 
	.A(n1174));
   SEN_INV_4 U291 (.X(net84442), 
	.A(net84445));
   SEN_ND2_4 U292 (.X(n1649), 
	.A2(n1603), 
	.A1(n1604));
   SEN_OAI22_4 U293 (.X(net83556), 
	.B2(n485), 
	.B1(net86274), 
	.A2(n484), 
	.A1(net86274));
   SEN_ND2_T_4 U294 (.X(net83870), 
	.A2(n482), 
	.A1(net83550));
   SEN_NR2_G_3 U295 (.X(net83826), 
	.A2(net83525), 
	.A1(net83740));
   SEN_INV_S_3 U296 (.X(net82827), 
	.A(net82838));
   SEN_NR2_S_5 U297 (.X(net83072), 
	.A2(net86086), 
	.A1(n68));
   SEN_ND2_4 U298 (.X(net83408), 
	.A2(n320), 
	.A1(n318));
   SEN_AO21B_2 U299 (.X(n947), 
	.B(n777), 
	.A2(n959), 
	.A1(net84220));
   SEN_ND2_S_3 U300 (.X(net87546), 
	.A2(n265), 
	.A1(net83607));
   SEN_ND2_T_3 U302 (.X(n470), 
	.A2(net83612), 
	.A1(net83611));
   SEN_NR2B_V1_4 U303 (.X(n1214), 
	.B(n1213), 
	.A(n1215));
   SEN_OR2_5 U304 (.X(n1215), 
	.A2(pprow7_qual[1]), 
	.A1(pprow6_qual[3]));
   SEN_ND2_T_8 U305 (.X(n1333), 
	.A2(n1237), 
	.A1(n1236));
   SEN_ND2_6 U306 (.X(n1236), 
	.A2(n257), 
	.A1(n1235));
   SEN_AOI21_S_8 U307 (.X(n1217), 
	.B(n1214), 
	.A2(pprow7_qual[1]), 
	.A1(pprow6_qual[3]));
   SEN_INV_4 U308 (.X(net82316), 
	.A(net82319));
   SEN_NR2_4 U309 (.X(net91110), 
	.A2(n1843), 
	.A1(n861));
   SEN_INV_1 U310 (.X(n1843), 
	.A(n808));
   SEN_EO2_S_3 U311 (.X(net83792), 
	.A2(n1086), 
	.A1(n1087));
   SEN_ND2_G_3 U312 (.X(n1183), 
	.A2(net83792), 
	.A1(n1129));
   SEN_INV_5 U313 (.X(net83681), 
	.A(net83792));
   SEN_INV_6 U314 (.X(n1451), 
	.A(n1327));
   SEN_ND2_S_4 U315 (.X(net84191), 
	.A2(net84189), 
	.A1(net84187));
   SEN_BUF_1 U316 (.X(n40), 
	.A(n314));
   SEN_OAI21B_2 U318 (.X(n452), 
	.B(net91120), 
	.A2(net2268), 
	.A1(n453));
   SEN_INV_6 U320 (.X(n315), 
	.A(n310));
   SEN_ND2_1P5 U321 (.X(n1441), 
	.A2(net83414), 
	.A1(net83415));
   SEN_EN2_0P5 U322 (.X(net83494), 
	.A2(n40), 
	.A1(n313));
   SEN_EO2_DG_1 U323 (.X(net83615), 
	.A2(net83497), 
	.A1(net83499));
   SEN_EN2_3 U325 (.X(n190), 
	.A2(n186), 
	.A1(n191));
   SEN_ND2_T_5 U326 (.X(n1035), 
	.A2(net87800), 
	.A1(net87799));
   SEN_ND2_6 U327 (.X(net83862), 
	.A2(n1066), 
	.A1(n1067));
   SEN_EN2_6 U328 (.X(n1066), 
	.A2(n1026), 
	.A1(n538));
   SEN_ND2_G_6 U329 (.X(n1105), 
	.A2(n1068), 
	.A1(n1069));
   SEN_INV_1P25 U330 (.X(n1842), 
	.A(n810));
   SEN_ND2_8 U334 (.X(net83453), 
	.A2(net87547), 
	.A1(net83608));
   SEN_AOI21B_0P5 U336 (.X(n42), 
	.B(n1161), 
	.A2(n467), 
	.A1(net83724));
   SEN_ND2_6 U337 (.X(n1161), 
	.A2(net83844), 
	.A1(net83843));
   SEN_INV_6 U338 (.X(net82234), 
	.A(net82238));
   SEN_EN2_3 U341 (.X(net84208), 
	.A2(n810), 
	.A1(pprow4_qual[0]));
   SEN_EN2_DG_8 U343 (.X(n43), 
	.A2(pprow14_qual[1]), 
	.A1(pprow13_qual[3]));
   SEN_ND2_S_2 U344 (.X(n861), 
	.A2(n619), 
	.A1(net87846));
   SEN_BUF_D_2 U346 (.X(n461), 
	.A(net83462));
   SEN_AO21B_8 U347 (.X(net86023), 
	.B(net83565), 
	.A2(net83583), 
	.A1(net83689));
   SEN_NR2_S_0P65 U348 (.X(n189), 
	.A2(pprow2_qual[6]), 
	.A1(pprow3_qual[4]));
   SEN_ND2_4 U349 (.X(net83574), 
	.A2(pprow2_qual[6]), 
	.A1(pprow3_qual[4]));
   SEN_INV_4 U350 (.X(n479), 
	.A(net83544));
   SEN_ND2_4 U351 (.X(net83544), 
	.A2(net83679), 
	.A1(net83678));
   SEN_ND3_S_2 U353 (.X(n1464), 
	.A3(n1583), 
	.A2(n1582), 
	.A1(n1463));
   SEN_EN2_S_2 U354 (.X(n1460), 
	.A2(n1463), 
	.A1(n670));
   SEN_ND2B_6 U355 (.X(n472), 
	.B(n476), 
	.A(net83454));
   SEN_INV_S_0P5 U356 (.X(n44), 
	.A(n882));
   SEN_EO2_S_3 U357 (.X(n1145), 
	.A2(n1143), 
	.A1(n746));
   SEN_ND2_S_3 U358 (.X(n1143), 
	.A2(n1166), 
	.A1(n812));
   SEN_EO2_S_3 U359 (.X(net84272), 
	.A2(n911), 
	.A1(n912));
   SEN_ND2_T_5 U363 (.X(net83168), 
	.A2(net83863), 
	.A1(net83862));
   SEN_ND2_T_2 U364 (.X(net83863), 
	.A2(n323), 
	.A1(net83845));
   SEN_ND2_T_2 U365 (.X(net82879), 
	.A2(net83158), 
	.A1(net83166));
   SEN_AOAI211_6 U367 (.X(net84227), 
	.C(net84353), 
	.B(net84352), 
	.A2(net84351), 
	.A1(net84350));
   SEN_EO2_0P5 U368 (.X(n680), 
	.A2(n1406), 
	.A1(n1405));
   SEN_ND2_T_1 U369 (.X(n1407), 
	.A2(n1405), 
	.A1(n1406));
   SEN_NR2_T_2 U370 (.X(n1408), 
	.A2(n1406), 
	.A1(n1405));
   SEN_NR2B_4 U371 (.X(n1036), 
	.B(net83951), 
	.A(n1055));
   SEN_INV_5 U372 (.X(net82354), 
	.A(net82349));
   SEN_EO2_S_6 U374 (.X(n1076), 
	.A2(n1057), 
	.A1(n47));
   SEN_EN2_DG_8 U375 (.X(n47), 
	.A2(n1094), 
	.A1(n1095));
   SEN_INV_S_4 U376 (.X(n251), 
	.A(n1184));
   SEN_AN2_6 U377 (.X(n1472), 
	.A2(n1475), 
	.A1(n1474));
   SEN_BUF_1 U378 (.X(n48), 
	.A(C[11]));
   SEN_BUF_1 U379 (.X(n49), 
	.A(n51));
   SEN_OAI21_5 U380 (.X(n51), 
	.B(n53), 
	.A2(net84108), 
	.A1(net84107));
   SEN_NR2_T_2 U382 (.X(net83523), 
	.A2(net83527), 
	.A1(net83528));
   SEN_AO2BB2_8 U383 (.X(net83528), 
	.B2(net84115), 
	.B1(net86698), 
	.A2(net84118), 
	.A1(net84119));
   SEN_ND2_G_1 U384 (.X(net83527), 
	.A2(net84110), 
	.A1(net84116));
   SEN_NR3_T_4 U386 (.X(net86559), 
	.A3(net83526), 
	.A2(net83524), 
	.A1(net83525));
   SEN_ND2_S_4 U387 (.X(net83525), 
	.A2(net83645), 
	.A1(net83649));
   SEN_INV_S_1 U388 (.X(net83524), 
	.A(net83646));
   SEN_INV_S_1 U389 (.X(net83526), 
	.A(net83520));
   SEN_AOI21B_8 U390 (.X(net86332), 
	.B(net83001), 
	.A2(net83000), 
	.A1(net82999));
   SEN_NR2_T_6 U392 (.X(net83649), 
	.A2(n50), 
	.A1(n51));
   SEN_ND2_1P5 U393 (.X(net83645), 
	.A2(pprow0_qual[14]), 
	.A1(C[14]));
   SEN_NR2_T_1P5 U394 (.X(net90704), 
	.A2(net83524), 
	.A1(net83525));
   SEN_ND2_T_3 U395 (.X(n50), 
	.A2(n52), 
	.A1(net83735));
   SEN_ND2_2 U396 (.X(net83735), 
	.A2(pprow0_qual[13]), 
	.A1(C[13]));
   SEN_ND2_G_1 U397 (.X(n52), 
	.A2(pprow0_qual[12]), 
	.A1(C[12]));
   SEN_OA2BB2_8 U398 (.X(net83933), 
	.B2(net100921), 
	.B1(net83828), 
	.A2(net83649), 
	.A1(net95928));
   SEN_AOI21B_3 U399 (.X(net83642), 
	.B(net83649), 
	.A2(net83648), 
	.A1(net83647));
   SEN_INV_S_6 U400 (.X(net84107), 
	.A(net84110));
   SEN_ND2B_S_4 U401 (.X(net84110), 
	.B(net84117), 
	.A(C[11]));
   SEN_ND2_T_2 U402 (.X(net84108), 
	.A2(pprow0_qual[10]), 
	.A1(C[10]));
   SEN_NR2B_V1_1 U404 (.X(net84025), 
	.B(n49), 
	.A(n52));
   SEN_INV_S_2 U405 (.X(net84117), 
	.A(pprow0_qual[11]));
   SEN_AN3B_8 U406 (.X(net86213), 
	.B2(net84110), 
	.B1(net86124), 
	.A(net84115));
   SEN_ND2_4 U407 (.X(net83070), 
	.A2(net83166), 
	.A1(net83165));
   SEN_INV_1 U409 (.X(net83159), 
	.A(net83070));
   SEN_OR4B_4 U410 (.X(net83205), 
	.B3(net83369), 
	.B2(n39), 
	.B1(net94359), 
	.A(net95846));
   SEN_EO2_8 U411 (.X(n56), 
	.A2(n59), 
	.A1(n58));
   SEN_INV_S_6 U412 (.X(n54), 
	.A(net83424));
   SEN_EN2_5 U413 (.X(net83424), 
	.A2(net83530), 
	.A1(net86010));
   SEN_INV_S_0P5 U414 (.X(net83422), 
	.A(n55));
   SEN_EN2_DG_8 U415 (.X(n58), 
	.A2(C[18]), 
	.A1(net83435));
   SEN_INV_2 U416 (.X(net83435), 
	.A(pprow0_qual[18]));
   SEN_AO21B_6 U417 (.X(n59), 
	.B(net83431), 
	.A2(net83434), 
	.A1(net86332));
   SEN_ND2B_V1_2 U418 (.X(net83434), 
	.B(net83516), 
	.A(C[17]));
   SEN_ND2_2 U419 (.X(net83431), 
	.A2(pprow0_qual[17]), 
	.A1(C[17]));
   SEN_AO21B_6 U421 (.X(net83001), 
	.B(net83520), 
	.A2(net83521), 
	.A1(net83522));
   SEN_EN3_DG_4 U422 (.X(net82838), 
	.A3(net82859), 
	.A2(net85257), 
	.A1(net82857));
   SEN_EN2_S_6 U424 (.X(net85257), 
	.A2(net82975), 
	.A1(net86279));
   SEN_AO21_DG_1 U425 (.X(net82859), 
	.B(net82884), 
	.A2(net82973), 
	.A1(net82972));
   SEN_OR2_2 U426 (.X(net82639), 
	.A2(net82829), 
	.A1(net82838));
   SEN_EN2_0P5 U428 (.X(n60), 
	.A2(net84634), 
	.A1(pprow10_qual[0]));
   SEN_ND2_8 U429 (.X(n61), 
	.A2(net82939), 
	.A1(n62));
   SEN_INV_1 U431 (.X(net82939), 
	.A(n60));
   SEN_AOAI211_6 U432 (.X(net82854), 
	.C(net82858), 
	.B(net82857), 
	.A2(net82856), 
	.A1(net82855));
   SEN_ND2B_V1_6 U433 (.X(n65), 
	.B(net82937), 
	.A(n67));
   SEN_AN2_12 U434 (.X(net82937), 
	.A2(net86556), 
	.A1(net86557));
   SEN_ND2_T_16 U435 (.X(n66), 
	.A2(n67), 
	.A1(n64));
   SEN_ND3B_V1DG_8 U436 (.X(net86557), 
	.B2(n70), 
	.B1(net94217), 
	.A(net95543));
   SEN_ND2B_V1_4 U437 (.X(net95543), 
	.B(net95561), 
	.A(net83174));
   SEN_NR2_T_8 U439 (.X(n70), 
	.A2(net95575), 
	.A1(n71));
   SEN_ND2_12 U441 (.X(net90814), 
	.A2(net83172), 
	.A1(net94132));
   SEN_NR2_S_5 U442 (.X(net95575), 
	.A2(net95557), 
	.A1(net95559));
   SEN_ND2_S_1 U443 (.X(n69), 
	.A2(net83076), 
	.A1(net83077));
   SEN_EO2_3 U444 (.X(net83077), 
	.A2(net83176), 
	.A1(net83175));
   SEN_EN2_S_2 U445 (.X(net82935), 
	.A2(net82938), 
	.A1(net82937));
   SEN_INV_0P8 U446 (.X(net82736), 
	.A(net82742));
   SEN_INV_2 U447 (.X(net83071), 
	.A(net83158));
   SEN_NR2B_V1_2 U448 (.X(n68), 
	.B(net83077), 
	.A(net95557));
   SEN_INV_4 U449 (.X(net95557), 
	.A(net83076));
   SEN_NR2_G_4 U450 (.X(net86086), 
	.A2(net83163), 
	.A1(net83164));
   SEN_AOI21_2 U451 (.X(net82875), 
	.B(net82743), 
	.A2(net102542), 
	.A1(net82742));
   SEN_NR2_1 U452 (.X(net82976), 
	.A2(net82742), 
	.A1(net82977));
   SEN_EO2_2 U453 (.X(Z[31]), 
	.A2(net82042), 
	.A1(net82041));
   SEN_ND2_T_2 U454 (.X(net82041), 
	.A2(n79), 
	.A1(net87948));
   SEN_INV_3 U457 (.X(net87947), 
	.A(net82065));
   SEN_AOAI211_6 U458 (.X(net82065), 
	.C(net82067), 
	.B(net82062), 
	.A2(net82059), 
	.A1(net82066));
   SEN_ND2_4 U459 (.X(n79), 
	.A2(net82065), 
	.A1(net87946));
   SEN_OA2BB2_4 U461 (.X(net82042), 
	.B2(net82046), 
	.B1(net86493), 
	.A2(net82044), 
	.A1(net82043));
   SEN_OAI21_5 U462 (.X(net82043), 
	.B(n75), 
	.A2(n74), 
	.A1(n73));
   SEN_EO2_S_6 U463 (.X(net82044), 
	.A2(n72), 
	.A1(net82047));
   SEN_ND2_T_4 U464 (.X(net82047), 
	.A2(net82062), 
	.A1(net82046));
   SEN_INV_5 U465 (.X(net82046), 
	.A(net82063));
   SEN_INV_8 U466 (.X(net82062), 
	.A(net82070));
   SEN_EO2_6 U467 (.X(n72), 
	.A2(net82050), 
	.A1(net82049));
   SEN_NR2_6 U468 (.X(net82049), 
	.A2(net82059), 
	.A1(net82052));
   SEN_EN2_5 U469 (.X(net82052), 
	.A2(net82075), 
	.A1(net82060));
   SEN_INV_1 U470 (.X(net82059), 
	.A(net82069));
   SEN_NR2_4 U471 (.X(net82050), 
	.A2(net82051), 
	.A1(net82052));
   SEN_EN3_6 U472 (.X(net82051), 
	.A3(net82055), 
	.A2(net95872), 
	.A1(net86468));
   SEN_EO2_S_3 U473 (.X(net86468), 
	.A2(net82057), 
	.A1(net82056));
   SEN_INV_S_1 U474 (.X(net82056), 
	.A(net82181));
   SEN_ND2_6 U475 (.X(net95872), 
	.A2(net82335), 
	.A1(net82336));
   SEN_EN3_6 U476 (.X(net82055), 
	.A3(net82179), 
	.A2(net85252), 
	.A1(net85931));
   SEN_ND2_T_4 U477 (.X(net86493), 
	.A2(net87543), 
	.A1(net87542));
   SEN_NR2_T_6 U478 (.X(n73), 
	.A2(n76), 
	.A1(net82306));
   SEN_NR2_T_4 U479 (.X(net82306), 
	.A2(net82311), 
	.A1(net88015));
   SEN_NR2B_V1DG_8 U480 (.X(net88015), 
	.B(net88014), 
	.A(net82309));
   SEN_ND2_T_4 U482 (.X(net82310), 
	.A2(net82430), 
	.A1(net88080));
   SEN_ND2_4 U483 (.X(net88080), 
	.A2(net88079), 
	.A1(net88078));
   SEN_ND2_T_3 U484 (.X(net82430), 
	.A2(net82523), 
	.A1(net82522));
   SEN_NR3_T_8 U485 (.X(net82311), 
	.A3(n78), 
	.A2(net82313), 
	.A1(n77));
   SEN_AN2_6 U486 (.X(n77), 
	.A2(net87944), 
	.A1(net87943));
   SEN_ND3_T_4 U487 (.X(net87943), 
	.A3(net82317), 
	.A2(net82316), 
	.A1(net82315));
   SEN_ND2_T_4 U488 (.X(net82315), 
	.A2(net82833), 
	.A1(net86553));
   SEN_OAI211_4 U489 (.X(net82317), 
	.B2(net82836), 
	.B1(net82827), 
	.A2(net82831), 
	.A1(net94176));
   SEN_INV_4 U490 (.X(net87944), 
	.A(net86518));
   SEN_OAI21_S_8 U491 (.X(net86518), 
	.B(net82638), 
	.A2(net91053), 
	.A1(net82636));
   SEN_ND2_T_6 U492 (.X(net82313), 
	.A2(net82431), 
	.A1(net82432));
   SEN_INV_S_4 U493 (.X(n76), 
	.A(net82308));
   SEN_ND2_4 U494 (.X(net82308), 
	.A2(net82324), 
	.A1(net82323));
   SEN_OAI21_5 U495 (.X(n74), 
	.B(net82302), 
	.A2(net86381), 
	.A1(net86498));
   SEN_EO2_8 U496 (.X(net82304), 
	.A2(net82285), 
	.A1(net82284));
   SEN_ND2_T_5 U497 (.X(net82305), 
	.A2(net91564), 
	.A1(net82376));
   SEN_EO2_S_6 U498 (.X(net86381), 
	.A2(net86382), 
	.A1(net82383));
   SEN_ND2B_V1_6 U499 (.X(net82302), 
	.B(net86491), 
	.A(net82323));
   SEN_ND2_2 U500 (.X(n75), 
	.A2(net86381), 
	.A1(net86498));
   SEN_EN2_S_1 U501 (.X(Z[30]), 
	.A2(net90316), 
	.A1(net82043));
   SEN_ND2_T_4 U502 (.X(net82319), 
	.A2(net82640), 
	.A1(net82639));
   SEN_ND2_4 U503 (.X(net82640), 
	.A2(net82821), 
	.A1(net82822));
   SEN_INV_S_0P5 U504 (.X(net90668), 
	.A(net82316));
   SEN_EO2_2 U505 (.X(net82829), 
	.A2(net83019), 
	.A1(net83018));
   SEN_BUF_1 U506 (.X(net102677), 
	.A(net82639));
   SEN_AOAI211_6 U507 (.X(n1300), 
	.C(n1229), 
	.B(n1230), 
	.A2(n1231), 
	.A1(n1232));
   SEN_ND2B_V1_3 U508 (.X(n1230), 
	.B(n1169), 
	.A(n1171));
   SEN_ND2B_V1_2 U509 (.X(n863), 
	.B(n377), 
	.A(n869));
   SEN_ND2_T_2 U510 (.X(n869), 
	.A2(pprow1_qual[0]), 
	.A1(n291));
   SEN_ND2_S_2 U511 (.X(n1620), 
	.A2(n1523), 
	.A1(n1524));
   SEN_INV_S_0P5 U512 (.X(n1102), 
	.A(n1125));
   SEN_ND2_6 U513 (.X(n310), 
	.A2(net83497), 
	.A1(net83498));
   SEN_ND2_6 U514 (.X(n579), 
	.A2(net83851), 
	.A1(n1103));
   SEN_ND2_6 U515 (.X(net82822), 
	.A2(n568), 
	.A1(net87837));
   SEN_OR2_2 U516 (.X(n266), 
	.A2(n1484), 
	.A1(net82889));
   SEN_ND2_T_6 U517 (.X(n1519), 
	.A2(n1484), 
	.A1(net82889));
   SEN_EN2_S_1 U518 (.X(n1420), 
	.A2(n1484), 
	.A1(net82889));
   SEN_EO2_6 U519 (.X(net82889), 
	.A2(net82703), 
	.A1(n125));
   SEN_ND3_S_8 U520 (.X(net83382), 
	.A3(net84365), 
	.A2(net84366), 
	.A1(net84364));
   SEN_INV_4 U521 (.X(net82745), 
	.A(net82741));
   SEN_NR3_T_4 U522 (.X(n336), 
	.A3(n339), 
	.A2(n338), 
	.A1(n337));
   SEN_INV_1P5 U523 (.X(n338), 
	.A(n352));
   SEN_AOI31_4 U524 (.X(n1142), 
	.B(n1130), 
	.A3(net83790), 
	.A2(net83789), 
	.A1(n1131));
   SEN_ND2_T_2 U525 (.X(net84239), 
	.A2(n89), 
	.A1(net84730));
   SEN_OAI211_4 U526 (.X(net84217), 
	.B2(net84191), 
	.B1(n306), 
	.A2(net83382), 
	.A1(net84362));
   SEN_ND3_T_6 U528 (.X(net83550), 
	.A3(n508), 
	.A2(n507), 
	.A1(n506));
   SEN_OAI221_2 U530 (.X(n508), 
	.C(n509), 
	.B2(net84059), 
	.B1(net84058), 
	.A2(net84057), 
	.A1(net84056));
   SEN_NR2_T_1P5 U531 (.X(net84412), 
	.A2(net84395), 
	.A1(net84413));
   SEN_AOAI211_8 U535 (.X(n1125), 
	.C(n1078), 
	.B(n1079), 
	.A2(n1080), 
	.A1(n1081));
   SEN_EN2_S_4 U536 (.X(net83611), 
	.A2(net83676), 
	.A1(n389));
   SEN_AN2_S_8 U538 (.X(net86321), 
	.A2(n487), 
	.A1(net83297));
   SEN_ND2_4 U541 (.X(net83848), 
	.A2(n295), 
	.A1(net83849));
   SEN_ND2B_V1_8 U542 (.X(net84183), 
	.B(net83383), 
	.A(net83382));
   SEN_ND2_T_2 U543 (.X(net84365), 
	.A2(n246), 
	.A1(n880));
   SEN_ND2_T_8 U544 (.X(net83512), 
	.A2(net83722), 
	.A1(net83721));
   SEN_ND2_T_2 U546 (.X(net82734), 
	.A2(net82983), 
	.A1(net94217));
   SEN_AOAI211_6 U547 (.X(n950), 
	.C(n918), 
	.B(n919), 
	.A2(n920), 
	.A1(n921));
   SEN_OAOI211_G_4 U548 (.X(n919), 
	.C(n894), 
	.B(n895), 
	.A2(n896), 
	.A1(n541));
   SEN_INV_6 U549 (.X(n898), 
	.A(n900));
   SEN_ND2_S_8 U550 (.X(net82973), 
	.A2(pprow10_qual[0]), 
	.A1(net84634));
   SEN_BUF_6 U551 (.X(net84634), 
	.A(\bmul/neg11 ));
   SEN_OAI21_4 U552 (.X(n1786), 
	.B(n1785), 
	.A2(pprow10_qual[7]), 
	.A1(pprow11_qual[5]));
   SEN_ND2B_V1DG_4 U553 (.X(n276), 
	.B(n85), 
	.A(n282));
   SEN_EO2_G_2 U554 (.X(n279), 
	.A2(pprow0_qual[2]), 
	.A1(net84732));
   SEN_ND2_4 U555 (.X(net82432), 
	.A2(net82520), 
	.A1(net82521));
   SEN_AO21_4 U556 (.X(n1065), 
	.B(n1269), 
	.A2(net84040), 
	.A1(n660));
   SEN_ND2_8 U557 (.X(net89993), 
	.A2(net84272), 
	.A1(net84273));
   SEN_EO2_4 U558 (.X(n1120), 
	.A2(n235), 
	.A1(n234));
   SEN_AN2_S_4 U559 (.X(net86124), 
	.A2(net84116), 
	.A1(net84159));
   SEN_ND2B_V1_6 U560 (.X(net84159), 
	.B(net84361), 
	.A(C[6]));
   SEN_INV_1 U561 (.X(net84356), 
	.A(net84159));
   SEN_OAI21_5 U562 (.X(n1816), 
	.B(n1794), 
	.A2(n1795), 
	.A1(n1796));
   SEN_OAOI211_G_8 U563 (.X(n1557), 
	.C(n1498), 
	.B(n1499), 
	.A2(pprow8_qual[6]), 
	.A1(pprow9_qual[4]));
   SEN_BUF_1 U566 (.X(n80), 
	.A(n1018));
   SEN_ND2_T_1 U567 (.X(n958), 
	.A2(n543), 
	.A1(n957));
   SEN_AO21B_6 U569 (.X(n1403), 
	.B(n1374), 
	.A2(n750), 
	.A1(n1373));
   SEN_INV_2 U570 (.X(n631), 
	.A(n1091));
   SEN_AOAI211_G_2 U571 (.X(n1091), 
	.C(net83572), 
	.B(net83889), 
	.A2(net83777), 
	.A1(n1135));
   SEN_EO2_6 U572 (.X(net87796), 
	.A2(net83459), 
	.A1(n385));
   SEN_EO2_0P5 U573 (.X(n677), 
	.A2(n1120), 
	.A1(n1121));
   SEN_ND2_T_1 U574 (.X(n1264), 
	.A2(n1121), 
	.A1(n1120));
   SEN_ND4_S_4 U575 (.X(net83639), 
	.A4(net83644), 
	.A3(n563), 
	.A2(net87761), 
	.A1(net83642));
   SEN_ND3_S_2 U576 (.X(n390), 
	.A3(n1714), 
	.A2(n1659), 
	.A1(net82436));
   SEN_INV_4 U577 (.X(n1643), 
	.A(n1647));
   SEN_ND2_T_6 U578 (.X(n92), 
	.A2(n91), 
	.A1(n90));
   SEN_INV_1P25 U579 (.X(n91), 
	.A(n698));
   SEN_OAI21_S_1P5 U580 (.X(net84220), 
	.B(net89993), 
	.A2(net84186), 
	.A1(net84192));
   SEN_EO2_S_6 U581 (.X(n1740), 
	.A2(n583), 
	.A1(n1759));
   SEN_ND2B_8 U582 (.X(net84350), 
	.B(n451), 
	.A(C[5]));
   SEN_ND2_2 U583 (.X(net83203), 
	.A2(net83174), 
	.A1(n45));
   SEN_ND2_T_3 U584 (.X(net84067), 
	.A2(n939), 
	.A1(n937));
   SEN_OAI21_3 U585 (.X(n1038), 
	.B(net84068), 
	.A2(net84067), 
	.A1(n955));
   SEN_ND2_T_1 U586 (.X(n1043), 
	.A2(net83951), 
	.A1(net83550));
   SEN_NR2_T_4 U587 (.X(n143), 
	.A2(n144), 
	.A1(n140));
   SEN_NR2_G_3 U588 (.X(n140), 
	.A2(n142), 
	.A1(n141));
   SEN_NR2_3 U589 (.X(n142), 
	.A2(n148), 
	.A1(net82721));
   SEN_EN2_S_4 U590 (.X(net85815), 
	.A2(n143), 
	.A1(n87));
   SEN_BUF_D_3 U591 (.X(n364), 
	.A(net82347));
   SEN_ND2_S_1P5 U592 (.X(n571), 
	.A2(net82347), 
	.A1(net82348));
   SEN_BUF_D_2 U593 (.X(net101269), 
	.A(net83521));
   SEN_INV_S_1P5 U594 (.X(net83936), 
	.A(pprow0_qual[13]));
   SEN_NR2_T_12 U595 (.X(net86477), 
	.A2(n502), 
	.A1(n242));
   SEN_INV_6 U597 (.X(net82983), 
	.A(net83170));
   SEN_ND2B_S_2 U598 (.X(net83607), 
	.B(n470), 
	.A(net83610));
   SEN_ND2_8 U599 (.X(net83559), 
	.A2(net83964), 
	.A1(n432));
   SEN_AO21B_6 U600 (.X(n1410), 
	.B(n1389), 
	.A2(n749), 
	.A1(n1388));
   SEN_ND2_2 U602 (.X(n994), 
	.A2(pprow1_qual[8]), 
	.A1(pprow1_qual[6]));
   SEN_OAI21_G_6 U603 (.X(n1007), 
	.B(n994), 
	.A2(n995), 
	.A1(n704));
   SEN_ND2_2 U604 (.X(n358), 
	.A2(net90738), 
	.A1(net82179));
   SEN_NR2_T_2 U605 (.X(net90738), 
	.A2(net91399), 
	.A1(net91396));
   SEN_EN2_3 U606 (.X(n661), 
	.A2(n1658), 
	.A1(n1657));
   SEN_INV_8 U607 (.X(net83647), 
	.A(net83528));
   SEN_AOAI211_3 U609 (.X(net82322), 
	.C(net82309), 
	.B(n393), 
	.A2(net82427), 
	.A1(net82426));
   SEN_INV_S_1P5 U610 (.X(n864), 
	.A(n863));
   SEN_ND2_S_4 U611 (.X(net83331), 
	.A2(net83332), 
	.A1(net83333));
   SEN_INV_8 U612 (.X(net83849), 
	.A(n207));
   SEN_EO3_DG_4 U614 (.X(net82082), 
	.A3(net85897), 
	.A2(net82102), 
	.A1(net82100));
   SEN_ND2_T_1 U615 (.X(n1562), 
	.A2(n1561), 
	.A1(net82717));
   SEN_NR2_S_3 U617 (.X(net83157), 
	.A2(net86086), 
	.A1(net83159));
   SEN_OAOI211_8 U618 (.X(n1511), 
	.C(n1472), 
	.B(n1473), 
	.A2(n1474), 
	.A1(n1475));
   SEN_EN2_5 U619 (.X(net82324), 
	.A2(n663), 
	.A1(n671));
   SEN_AO21B_8 U620 (.X(net83169), 
	.B(net83373), 
	.A2(net83372), 
	.A1(net83371));
   SEN_INV_1P25 U621 (.X(net84286), 
	.A(net84153));
   SEN_OAI21_G_4 U622 (.X(n1652), 
	.B(n1595), 
	.A2(n1596), 
	.A1(n1597));
   SEN_INV_S_1P5 U623 (.X(n1493), 
	.A(n1545));
   SEN_ND2_8 U625 (.X(n1104), 
	.A2(n580), 
	.A1(net83852));
   SEN_INV_S_4 U626 (.X(net84393), 
	.A(net84394));
   SEN_INV_S_6 U628 (.X(net103418), 
	.A(net82062));
   SEN_ND2_G_3 U630 (.X(n556), 
	.A2(n1006), 
	.A1(n1005));
   SEN_AOI211_G_3 U631 (.X(n1006), 
	.B2(n1198), 
	.B1(n1000), 
	.A2(n1001), 
	.A1(n1002));
   SEN_ND2_G_1 U632 (.X(net85838), 
	.A2(n582), 
	.A1(net94287));
   SEN_ND3_T_6 U633 (.X(n207), 
	.A3(n1104), 
	.A2(n1105), 
	.A1(n1106));
   SEN_INV_4 U634 (.X(n585), 
	.A(n584));
   SEN_INV_5 U635 (.X(n293), 
	.A(net83631));
   SEN_EO2_DG_1 U636 (.X(net83097), 
	.A2(n685), 
	.A1(n1376));
   SEN_ND2_4 U639 (.X(net82376), 
	.A2(n585), 
	.A1(n776));
   SEN_OR4_4 U640 (.X(n1147), 
	.A4(n998), 
	.A3(n1199), 
	.A2(n1193), 
	.A1(n554));
   SEN_INV_1P5 U641 (.X(n554), 
	.A(n1201));
   SEN_ND2_S_4 U642 (.X(n998), 
	.A2(n999), 
	.A1(n923));
   SEN_ND3_S_2 U643 (.X(n1155), 
	.A3(n1147), 
	.A2(n1190), 
	.A1(n620));
   SEN_OAI21_5 U645 (.X(n232), 
	.B(n230), 
	.A2(n135), 
	.A1(net85351));
   SEN_NR2_2 U648 (.X(n230), 
	.A2(n221), 
	.A1(n219));
   SEN_OR2_2 U649 (.X(n99), 
	.A2(n1490), 
	.A1(net82876));
   SEN_ND2_S_4 U650 (.X(n1593), 
	.A2(n1490), 
	.A1(net82876));
   SEN_EO3_4 U651 (.X(n1490), 
	.A3(pprow0_qual[23]), 
	.A2(C[23]), 
	.A1(n1491));
   SEN_ND2_4 U653 (.X(n1482), 
	.A2(n1414), 
	.A1(n1412));
   SEN_AOI211_12 U654 (.X(net94314), 
	.B2(n1391), 
	.B1(net83108), 
	.A2(pprow3_qual[13]), 
	.A1(pprow2_qual[15]));
   SEN_ND2_S_3 U655 (.X(net84394), 
	.A2(pprow0_qual[0]), 
	.A1(C[0]));
   SEN_ND2B_V1_6 U656 (.X(n568), 
	.B(net87836), 
	.A(net86446));
   SEN_ND2_6 U657 (.X(net82638), 
	.A2(net82823), 
	.A1(net82824));
   SEN_INV_S_0P5 U658 (.X(n1436), 
	.A(n1490));
   SEN_INV_3 U659 (.X(net87828), 
	.A(net87827));
   SEN_INV_4 U660 (.X(net83722), 
	.A(net83723));
   SEN_ND2B_S_0P5 U661 (.X(n395), 
	.B(n1725), 
	.A(n547));
   SEN_EO2_G_2 U662 (.X(net82386), 
	.A2(n696), 
	.A1(n1722));
   SEN_ND2_G_1 U663 (.X(net82245), 
	.A2(net82247), 
	.A1(net82246));
   SEN_EO2_8 U665 (.X(net83454), 
	.A2(net83535), 
	.A1(net83534));
   SEN_AOI21_6 U666 (.X(net83535), 
	.B(net83538), 
	.A2(net83537), 
	.A1(n481));
   SEN_NR2_S_3 U667 (.X(net83537), 
	.A2(net86385), 
	.A1(net83547));
   SEN_ND3_T_8 U668 (.X(n486), 
	.A3(net83952), 
	.A2(net83552), 
	.A1(net83951));
   SEN_INV_6 U669 (.X(net91397), 
	.A(net91418));
   SEN_EN2_3 U670 (.X(net90631), 
	.A2(net91418), 
	.A1(n517));
   SEN_AOAI211_8 U671 (.X(net91418), 
	.C(net91419), 
	.B(net91426), 
	.A2(net91390), 
	.A1(net91392));
   SEN_ND2B_S_8 U672 (.X(net83385), 
	.B(net83510), 
	.A(net83505));
   SEN_ND2_4 U673 (.X(n1268), 
	.A2(net83506), 
	.A1(net83505));
   SEN_ND2_T_2 U674 (.X(net83369), 
	.A2(net83385), 
	.A1(net83384));
   SEN_ND2_6 U675 (.X(net83679), 
	.A2(n640), 
	.A1(n639));
   SEN_NR2_T_6 U676 (.X(n325), 
	.A2(n326), 
	.A1(net82847));
   SEN_ND2_T_3 U677 (.X(net84275), 
	.A2(net84193), 
	.A1(net84276));
   SEN_ND2_6 U678 (.X(n1714), 
	.A2(net82773), 
	.A1(net82772));
   SEN_INV_S_1P5 U679 (.X(net84418), 
	.A(net84392));
   SEN_ND2_T_6 U680 (.X(n1413), 
	.A2(n1483), 
	.A1(n1481));
   SEN_OAI21_5 U682 (.X(n1345), 
	.B(n1305), 
	.A2(net83293), 
	.A1(net83292));
   SEN_ND2B_V1DG_4 U683 (.X(n1583), 
	.B(n1421), 
	.A(n1423));
   SEN_INV_0P65 U684 (.X(net83547), 
	.A(net83302));
   SEN_AN4B_4 U685 (.X(net83292), 
	.B3(net83302), 
	.B2(net83301), 
	.B1(net83300), 
	.A(net83303));
   SEN_ND2_T_3 U687 (.X(net83304), 
	.A2(net87790), 
	.A1(net83681));
   SEN_ND2_T_8 U688 (.X(net83172), 
	.A2(n237), 
	.A1(n1205));
   SEN_INV_S_6 U690 (.X(n1342), 
	.A(n1339));
   SEN_EO2_5 U692 (.X(net82581), 
	.A2(n1577), 
	.A1(n250));
   SEN_EN2_3 U693 (.X(net82595), 
	.A2(n404), 
	.A1(n413));
   SEN_NR2_S_0P8 U694 (.X(n1260), 
	.A2(net85071), 
	.A1(net83422));
   SEN_ND2_S_3 U695 (.X(net82980), 
	.A2(net82982), 
	.A1(net82981));
   SEN_OA2BB2_4 U696 (.X(n1319), 
	.B2(n1315), 
	.B1(n1316), 
	.A2(n1317), 
	.A1(n1318));
   SEN_ND2B_S_2 U697 (.X(n1317), 
	.B(n1313), 
	.A(n1314));
   SEN_INV_3 U698 (.X(n1318), 
	.A(n1320));
   SEN_OAI211_4 U699 (.X(n1321), 
	.B2(n1306), 
	.B1(n1307), 
	.A2(n1308), 
	.A1(n1309));
   SEN_EO2_DG_2 U700 (.X(n1588), 
	.A2(n682), 
	.A1(n1560));
   SEN_ND2_S_4 U702 (.X(n643), 
	.A2(n391), 
	.A1(n390));
   SEN_ND2_T_2 U703 (.X(net83299), 
	.A2(net83461), 
	.A1(net83462));
   SEN_ND2_T_8 U704 (.X(n1520), 
	.A2(n647), 
	.A1(n1481));
   SEN_AOI31_4 U705 (.X(n1486), 
	.B(n1485), 
	.A3(n1520), 
	.A2(n245), 
	.A1(n1518));
   SEN_ND2_T_8 U706 (.X(n298), 
	.A2(net84196), 
	.A1(net89993));
   SEN_ND2_4 U708 (.X(n1078), 
	.A2(n1077), 
	.A1(n1076));
   SEN_EN2_S_8 U709 (.X(net82060), 
	.A2(n505), 
	.A1(net82082));
   SEN_ND2B_V1_3 U711 (.X(net82965), 
	.B(net83499), 
	.A(net83497));
   SEN_INV_4 U713 (.X(n1067), 
	.A(n1069));
   SEN_AOAI211_8 U714 (.X(net82243), 
	.C(n362), 
	.B(net82349), 
	.A2(net82348), 
	.A1(n364));
   SEN_OAI21_S_8 U715 (.X(n480), 
	.B(n2048), 
	.A2(n479), 
	.A1(net86333));
   SEN_INV_3 U717 (.X(net84251), 
	.A(net84007));
   SEN_INV_6 U718 (.X(net82436), 
	.A(net82854));
   SEN_INV_1 U719 (.X(n228), 
	.A(n232));
   SEN_EO2_S_3 U720 (.X(n1387), 
	.A2(net87351), 
	.A1(n649));
   SEN_ND2_4 U721 (.X(n500), 
	.A2(net82586), 
	.A1(net82587));
   SEN_AO21B_1 U723 (.X(net83993), 
	.B(n1011), 
	.A2(n1030), 
	.A1(n1029));
   SEN_NR2_T_3 U724 (.X(n1031), 
	.A2(n1029), 
	.A1(n1030));
   SEN_BUF_1 U725 (.X(n819), 
	.A(n1842));
   SEN_INV_S_0P5 U726 (.X(net84218), 
	.A(net84275));
   SEN_ND2_1P5 U727 (.X(n450), 
	.A2(n442), 
	.A1(net84228));
   SEN_ND2B_1 U728 (.X(n1465), 
	.B(n1582), 
	.A(n1579));
   SEN_EO2_S_1 U729 (.X(n670), 
	.A2(n1423), 
	.A1(n1421));
   SEN_ND2_T_1 U730 (.X(n1579), 
	.A2(n1422), 
	.A1(n1423));
   SEN_AO21B_6 U731 (.X(net82457), 
	.B(net82564), 
	.A2(n371), 
	.A1(net82565));
   SEN_OAI21_S_8 U732 (.X(net82565), 
	.B(net82658), 
	.A2(n111), 
	.A1(n350));
   SEN_OA2BB2_2 U733 (.X(net82083), 
	.B2(net85931), 
	.B1(net86266), 
	.A2(net82173), 
	.A1(net82057));
   SEN_ND2_S_2 U734 (.X(net82173), 
	.A2(net86266), 
	.A1(net85931));
   SEN_EO2_4 U735 (.X(net82513), 
	.A2(n664), 
	.A1(n1674));
   SEN_EO2_8 U736 (.X(n505), 
	.A2(net91024), 
	.A1(net82201));
   SEN_ND2_T_5 U737 (.X(n1582), 
	.A2(n1580), 
	.A1(n1581));
   SEN_INV_4 U738 (.X(n1418), 
	.A(n1413));
   SEN_BUF_3 U739 (.X(n289), 
	.A(C[0]));
   SEN_INV_0P65 U740 (.X(net87845), 
	.A(n289));
   SEN_ND2B_V1_4 U744 (.X(net84276), 
	.B(net84274), 
	.A(net84272));
   SEN_ND2_S_2 U745 (.X(n1809), 
	.A2(n1808), 
	.A1(n701));
   SEN_NR2_S_4 U746 (.X(n537), 
	.A2(n1152), 
	.A1(n1150));
   SEN_EO3_4 U747 (.X(n920), 
	.A3(net84272), 
	.A2(net89992), 
	.A1(n699));
   SEN_EN2_2 U748 (.X(n1734), 
	.A2(n1671), 
	.A1(n1727));
   SEN_EO2_5 U749 (.X(n1095), 
	.A2(n757), 
	.A1(n756));
   SEN_ND2_T_3 U750 (.X(net83685), 
	.A2(n1095), 
	.A1(n1094));
   SEN_AOAI211_8 U751 (.X(net83308), 
	.C(net83870), 
	.B(n1098), 
	.A2(net83555), 
	.A1(net83556));
   SEN_OR4B_2 U752 (.X(n1491), 
	.B3(n1433), 
	.B2(n1434), 
	.B1(n1435), 
	.A(n1432));
   SEN_ND2_2 U753 (.X(net82460), 
	.A2(net82462), 
	.A1(n370));
   SEN_ND2_2 U754 (.X(net84435), 
	.A2(n879), 
	.A1(net84437));
   SEN_INV_S_6 U758 (.X(n580), 
	.A(n579));
   SEN_ND2B_V1_6 U759 (.X(net83852), 
	.B(n1021), 
	.A(n1019));
   SEN_AOAI211_3 U760 (.X(n1775), 
	.C(n1747), 
	.B(n1748), 
	.A2(n1749), 
	.A1(n1750));
   SEN_INV_3 U761 (.X(n1748), 
	.A(n1744));
   SEN_EN2_4 U762 (.X(n1628), 
	.A2(n1591), 
	.A1(n520));
   SEN_NR2_T_4 U763 (.X(n1245), 
	.A2(net87795), 
	.A1(n630));
   SEN_AN2_3 U764 (.X(n630), 
	.A2(net86321), 
	.A1(net83308));
   SEN_EO2_DG_8 U765 (.X(n82), 
	.A2(pprow1_qual[12]), 
	.A1(pprow1_qual[14]));
   SEN_EN2_S_2 U767 (.X(net82189), 
	.A2(n498), 
	.A1(n395));
   SEN_NR3_T_4 U768 (.X(n272), 
	.A3(n274), 
	.A2(n270), 
	.A1(n273));
   SEN_OAOI211_4 U770 (.X(net83676), 
	.C(n479), 
	.B(net86333), 
	.A2(net83546), 
	.A1(net83677));
   SEN_EN2_5 U771 (.X(n1033), 
	.A2(net84066), 
	.A1(net85880));
   SEN_NR2_T_6 U772 (.X(net84066), 
	.A2(net84200), 
	.A1(n651));
   SEN_INV_S_3 U774 (.X(n1135), 
	.A(n1090));
   SEN_AN2_5 U775 (.X(n469), 
	.A2(net83094), 
	.A1(net83103));
   SEN_NR2_T_4 U776 (.X(net86553), 
	.A2(net88104), 
	.A1(net88103));
   SEN_ND2_2 U778 (.X(n1455), 
	.A2(n1328), 
	.A1(n1451));
   SEN_NR2_T_4 U779 (.X(net83731), 
	.A2(net83733), 
	.A1(n1160));
   SEN_ND2_8 U780 (.X(n1701), 
	.A2(n1699), 
	.A1(n92));
   SEN_ND2_4 U781 (.X(net84000), 
	.A2(pprow3_qual[1]), 
	.A1(pprow2_qual[3]));
   SEN_INV_5 U782 (.X(n940), 
	.A(pprow3_qual[1]));
   SEN_ND2B_4 U783 (.X(n198), 
	.B(net84001), 
	.A(net87549));
   SEN_INV_1P25 U784 (.X(net84248), 
	.A(net87549));
   SEN_AOAI211_6 U786 (.X(n1793), 
	.C(n1719), 
	.B(net82420), 
	.A2(n1720), 
	.A1(n1721));
   SEN_AOAI211_6 U787 (.X(net82142), 
	.C(n1812), 
	.B(n1813), 
	.A2(n1814), 
	.A1(n1815));
   SEN_EO2_4 U788 (.X(net82102), 
	.A2(n733), 
	.A1(n1813));
   SEN_AOAI211_2 U789 (.X(n84), 
	.C(n322), 
	.B(net84443), 
	.A2(net84442), 
	.A1(net94322));
   SEN_OR2_5 U791 (.X(n645), 
	.A2(n1660), 
	.A1(n1661));
   SEN_EN2_S_3 U792 (.X(n1661), 
	.A2(n1657), 
	.A1(n1658));
   SEN_AOAI211_6 U793 (.X(n321), 
	.C(n322), 
	.B(net84443), 
	.A2(net84442), 
	.A1(net94322));
   SEN_ND2_12 U794 (.X(n1805), 
	.A2(net82394), 
	.A1(net82395));
   SEN_ND2_4 U795 (.X(net83631), 
	.A2(net83634), 
	.A1(net83636));
   SEN_ND2_6 U797 (.X(n1453), 
	.A2(n2039), 
	.A1(n1450));
   SEN_AOI21_T_4 U799 (.X(n1419), 
	.B(n1417), 
	.A2(n1418), 
	.A1(n1482));
   SEN_ND3_T_3 U800 (.X(n1530), 
	.A3(n536), 
	.A2(n1465), 
	.A1(n1464));
   SEN_AOAI211_8 U802 (.X(n1718), 
	.C(n1681), 
	.B(n1682), 
	.A2(n1683), 
	.A1(n1684));
   SEN_ND2_4 U803 (.X(n1401), 
	.A2(n1371), 
	.A1(n1372));
   SEN_INV_S_6 U805 (.X(net84119), 
	.A(net84147));
   SEN_INV_4 U806 (.X(net84241), 
	.A(net84157));
   SEN_EN2_S_3 U807 (.X(n957), 
	.A2(net84226), 
	.A1(n531));
   SEN_EN2_DG_8 U808 (.X(n370), 
	.A2(net82457), 
	.A1(n372));
   SEN_AO21B_6 U809 (.X(n350), 
	.B(n351), 
	.A2(net82758), 
	.A1(n349));
   SEN_INV_S_3 U810 (.X(net87547), 
	.A(net87546));
   SEN_AOI21B_8 U812 (.X(n1205), 
	.B(n1161), 
	.A2(n467), 
	.A1(net83724));
   SEN_INV_AS_5 U813 (.X(net82455), 
	.A(net82457));
   SEN_OR3_6 U814 (.X(net86257), 
	.A3(net83585), 
	.A2(n1134), 
	.A1(net83778));
   SEN_INV_4 U816 (.X(n312), 
	.A(net83408));
   SEN_ND2_4 U817 (.X(n918), 
	.A2(n916), 
	.A1(n917));
   SEN_INV_S_6 U818 (.X(net84362), 
	.A(net83383));
   SEN_ND2_S_2 U819 (.X(n100), 
	.A2(net83559), 
	.A1(n423));
   SEN_AOI211_8 U820 (.X(n1478), 
	.B2(n1391), 
	.B1(net83108), 
	.A2(pprow3_qual[13]), 
	.A1(pprow2_qual[15]));
   SEN_INV_4 U821 (.X(net83108), 
	.A(n231));
   SEN_ND2_G_3 U822 (.X(net82197), 
	.A2(net82582), 
	.A1(net82581));
   SEN_EO2_DG_2 U823 (.X(n685), 
	.A2(n1377), 
	.A1(n1378));
   SEN_ND2_T_4 U824 (.X(n440), 
	.A2(net95563), 
	.A1(net90814));
   SEN_AO21B_4 U826 (.X(n210), 
	.B(n1268), 
	.A2(n2042), 
	.A1(net83418));
   SEN_ND2_4 U827 (.X(n354), 
	.A2(pprow1_qual[19]), 
	.A1(n353));
   SEN_AN3_S_2 U828 (.X(n94), 
	.A3(n526), 
	.A2(n1274), 
	.A1(n1272));
   SEN_AN2_S_4 U831 (.X(n698), 
	.A2(n1647), 
	.A1(net82550));
   SEN_ND2_2 U832 (.X(n1497), 
	.A2(n1593), 
	.A1(n1592));
   SEN_ND2_T_1 U834 (.X(n874), 
	.A2(net84404), 
	.A1(n809));
   SEN_AOAI211_6 U835 (.X(n1817), 
	.C(n1806), 
	.B(n1807), 
	.A2(net82203), 
	.A1(net82202));
   SEN_ND2B_V1_6 U836 (.X(net82899), 
	.B(n402), 
	.A(net94314));
   SEN_EN2_S_4 U837 (.X(n1414), 
	.A2(net94314), 
	.A1(n376));
   SEN_INV_3 U838 (.X(n316), 
	.A(net83413));
   SEN_ND2B_V1DG_4 U839 (.X(net83413), 
	.B(net84045), 
	.A(net84046));
   SEN_EN2_8 U840 (.X(n900), 
	.A2(net86299), 
	.A1(n106));
   SEN_OR2_5 U841 (.X(net86299), 
	.A2(net84283), 
	.A1(n450));
   SEN_ND2_T_6 U842 (.X(n327), 
	.A2(net83334), 
	.A1(net87796));
   SEN_ND2_T_2 U843 (.X(n1055), 
	.A2(net83875), 
	.A1(n1034));
   SEN_INV_S_6 U844 (.X(n1034), 
	.A(n1035));
   SEN_INV_S_6 U845 (.X(net82467), 
	.A(net82462));
   SEN_INV_0P65 U846 (.X(n1547), 
	.A(n1596));
   SEN_AOI21_S_1 U848 (.X(net83630), 
	.B(n300), 
	.A2(net83513), 
	.A1(net83512));
   SEN_EO2_G_8 U849 (.X(net83721), 
	.A2(net83825), 
	.A1(n1116));
   SEN_ND2_T_5 U850 (.X(n1646), 
	.A2(n1644), 
	.A1(n1645));
   SEN_ND2B_V1DG_4 U851 (.X(n352), 
	.B(n353), 
	.A(n335));
   SEN_AN3_2 U852 (.X(n481), 
	.A3(n264), 
	.A2(n263), 
	.A1(n2046));
   SEN_EO2_0P5 U854 (.X(n741), 
	.A2(pprow3_qual[1]), 
	.A1(pprow2_qual[3]));
   SEN_EN2_S_2 U855 (.X(net82079), 
	.A2(net91024), 
	.A1(net82080));
   SEN_NR2_G_2 U856 (.X(net83303), 
	.A2(n479), 
	.A1(net83304));
   SEN_ND2_T_3 U857 (.X(net84068), 
	.A2(n513), 
	.A1(n511));
   SEN_AOI21_G_8 U859 (.X(net82404), 
	.B(n405), 
	.A2(n404), 
	.A1(n411));
   SEN_EO2_S_3 U860 (.X(n495), 
	.A2(net82206), 
	.A1(net82207));
   SEN_EO3_6 U861 (.X(net82206), 
	.A3(n1798), 
	.A2(n1797), 
	.A1(n252));
   SEN_OAI21_S_4 U862 (.X(n1138), 
	.B(n1176), 
	.A2(n1308), 
	.A1(n1084));
   SEN_OR4B_8 U864 (.X(n311), 
	.B3(n316), 
	.B2(net96981), 
	.B1(n315), 
	.A(net83412));
   SEN_EO2_G_4 U865 (.X(net84189), 
	.A2(n885), 
	.A1(n712));
   SEN_OAOI211_4 U866 (.X(n294), 
	.C(net83630), 
	.B(net83508), 
	.A2(net83168), 
	.A1(net83629));
   SEN_ND2_T_2 U867 (.X(n885), 
	.A2(n877), 
	.A1(n926));
   SEN_INV_2 U868 (.X(net82061), 
	.A(net82075));
   SEN_ND2_3 U869 (.X(n1322), 
	.A2(n604), 
	.A1(n1382));
   SEN_NR2_T_1 U870 (.X(n270), 
	.A2(n271), 
	.A1(net84394));
   SEN_OA21_4 U872 (.X(net102542), 
	.B(net82980), 
	.A2(net95559), 
	.A1(net95557));
   SEN_EO2_1 U874 (.X(net84404), 
	.A2(net84433), 
	.A1(n84));
   SEN_EN2_DG_1 U875 (.X(net84433), 
	.A2(n867), 
	.A1(n539));
   SEN_ND2_2 U876 (.X(net87827), 
	.A2(net83381), 
	.A1(net84177));
   SEN_ND3_T_2 U877 (.X(net84177), 
	.A3(n206), 
	.A2(n292), 
	.A1(net84183));
   SEN_ND2_2 U878 (.X(n1263), 
	.A2(n24), 
	.A1(net83919));
   SEN_INV_3 U879 (.X(n1351), 
	.A(n1350));
   SEN_ND2_T_2 U880 (.X(net82431), 
	.A2(net82636), 
	.A1(net91053));
   SEN_AO21B_8 U881 (.X(n1517), 
	.B(n1477), 
	.A2(n754), 
	.A1(n1476));
   SEN_AOAI211_6 U882 (.X(n1320), 
	.C(n117), 
	.B(n1310), 
	.A2(n1311), 
	.A1(n1312));
   SEN_OR2_2 U883 (.X(n1312), 
	.A2(pprow5_qual[6]), 
	.A1(pprow4_qual[8]));
   SEN_ND2_4 U884 (.X(net84029), 
	.A2(net100928), 
	.A1(net84111));
   SEN_AO21B_8 U885 (.X(net83629), 
	.B(net83848), 
	.A2(net83849), 
	.A1(n299));
   SEN_ND2_T_3 U886 (.X(net83381), 
	.A2(net84275), 
	.A1(n292));
   SEN_AOI22_T_3 U887 (.X(n1427), 
	.B2(pprow0_qual[20]), 
	.B1(C[20]), 
	.A2(n1367), 
	.A1(n1368));
   SEN_ND2_S_2 U888 (.X(n1394), 
	.A2(n1425), 
	.A1(n1427));
   SEN_EN2_S_3 U889 (.X(net82247), 
	.A2(net82251), 
	.A1(n1791));
   SEN_ND2_S_4 U890 (.X(net83064), 
	.A2(net101261), 
	.A1(n452));
   SEN_INV_S_6 U891 (.X(net88104), 
	.A(net82836));
   SEN_EN2_S_2 U892 (.X(n453), 
	.A2(net83152), 
	.A1(n454));
   SEN_NR2_T_2 U893 (.X(net84450), 
	.A2(pprow0_qual[2]), 
	.A1(net84732));
   SEN_INV_AS_10 U894 (.X(net88079), 
	.A(net82428));
   SEN_INV_8 U895 (.X(n307), 
	.A(net84187));
   SEN_ND2_T_1 U896 (.X(n1347), 
	.A2(n604), 
	.A1(n1346));
   SEN_EO2_DG_2 U898 (.X(n465), 
	.A2(net83096), 
	.A1(net83097));
   SEN_INV_AS_10 U899 (.X(n1677), 
	.A(n1676));
   SEN_EN2_5 U900 (.X(n1676), 
	.A2(n32), 
	.A1(n1609));
   SEN_INV_S_1 U901 (.X(n462), 
	.A(n1677));
   SEN_EO2_S_6 U902 (.X(net82428), 
	.A2(net82512), 
	.A1(net86466));
   SEN_EO2_G_2 U903 (.X(net86466), 
	.A2(net82513), 
	.A1(net82514));
   SEN_ND2_T_5 U904 (.X(n1663), 
	.A2(n1714), 
	.A1(net82436));
   SEN_ND2_T_5 U905 (.X(n1650), 
	.A2(net82770), 
	.A1(net82771));
   SEN_EO2_6 U906 (.X(net82771), 
	.A2(n107), 
	.A1(n1497));
   SEN_NR2_G_4 U907 (.X(net83372), 
	.A2(net83376), 
	.A1(n1269));
   SEN_INV_S_3 U909 (.X(n1253), 
	.A(n1252));
   SEN_ND2_3 U910 (.X(n1252), 
	.A2(pprow1_qual[13]), 
	.A1(pprow1_qual[15]));
   SEN_ND2_3 U911 (.X(n1743), 
	.A2(n1715), 
	.A1(n1765));
   SEN_INV_1P5 U912 (.X(n1766), 
	.A(n1765));
   SEN_NR2B_2 U913 (.X(n317), 
	.B(net86390), 
	.A(net83817));
   SEN_BUF_S_3 U914 (.X(net97377), 
	.A(net84217));
   SEN_ND2_S_3 U915 (.X(net83817), 
	.A2(n980), 
	.A1(n981));
   SEN_ND2_T_4 U916 (.X(net83890), 
	.A2(net84013), 
	.A1(net84012));
   SEN_INV_4 U917 (.X(net84013), 
	.A(pprow3_qual[4]));
   SEN_INV_2 U918 (.X(net84012), 
	.A(pprow2_qual[6]));
   SEN_ND2_T_5 U919 (.X(n1553), 
	.A2(n1650), 
	.A1(n1663));
   SEN_ND2_T_2 U920 (.X(n1358), 
	.A2(n1276), 
	.A1(n1277));
   SEN_AOAI211_8 U922 (.X(net83090), 
	.C(n1361), 
	.B(n1362), 
	.A2(n397), 
	.A1(n1363));
   SEN_AO21B_6 U923 (.X(n1362), 
	.B(n770), 
	.A2(net83189), 
	.A1(n1360));
   SEN_NR2_T_4 U925 (.X(n1307), 
	.A2(n1177), 
	.A1(n1178));
   SEN_ND2_T_8 U926 (.X(n1481), 
	.A2(n1385), 
	.A1(n1384));
   SEN_INV_6 U927 (.X(net83549), 
	.A(net83540));
   SEN_ND3_S_12 U928 (.X(net82831), 
	.A3(net82845), 
	.A2(net82846), 
	.A1(n325));
   SEN_AOAI211_8 U929 (.X(net82846), 
	.C(net86517), 
	.B(n1445), 
	.A2(n1446), 
	.A1(n1447));
   SEN_EN2_S_3 U930 (.X(net87790), 
	.A2(n1092), 
	.A1(n1093));
   SEN_ND2B_V1DG_2 U931 (.X(n1242), 
	.B(n1241), 
	.A(n1314));
   SEN_INV_S_4 U932 (.X(n604), 
	.A(n603));
   SEN_NR2B_4 U933 (.X(n1346), 
	.B(n648), 
	.A(net86321));
   SEN_ND2_T_8 U934 (.X(net82395), 
	.A2(n1673), 
	.A1(n1674));
   SEN_AOAI211_8 U935 (.X(net82100), 
	.C(net82235), 
	.B(net82234), 
	.A2(net82233), 
	.A1(n494));
   SEN_ND2B_V1DG_8 U936 (.X(net83507), 
	.B(net83846), 
	.A(net83168));
   SEN_INV_4 U937 (.X(net83846), 
	.A(net83629));
   SEN_OAI21_S_8 U938 (.X(n1626), 
	.B(n1619), 
	.A2(n2101), 
	.A1(net82595));
   SEN_OAOI211_4 U939 (.X(n1086), 
	.C(n637), 
	.B(n1085), 
	.A2(n399), 
	.A1(n1180));
   SEN_EO2_DG_8 U942 (.X(n86), 
	.A2(pprow11_qual[0]), 
	.A1(pprow10_qual[2]));
   SEN_INV_S_1 U943 (.X(net82884), 
	.A(net82768));
   SEN_AO21_4 U944 (.X(n757), 
	.B(n1308), 
	.A2(n1084), 
	.A1(n399));
   SEN_INV_4 U946 (.X(n1144), 
	.A(n1145));
   SEN_EN2_DG_8 U947 (.X(n87), 
	.A2(pprow7_qual[11]), 
	.A1(pprow6_qual[13]));
   SEN_OAI21_S_4 U949 (.X(net83786), 
	.B(net84001), 
	.A2(net95748), 
	.A1(net83999));
   SEN_AOI22_T_4 U951 (.X(n1762), 
	.B2(C[27]), 
	.B1(pprow0_qual[27]), 
	.A2(n1706), 
	.A1(n1705));
   SEN_OR2_5 U952 (.X(net83300), 
	.A2(net83461), 
	.A1(net83462));
   SEN_INV_S_3 U954 (.X(n866), 
	.A(pprow0_qual[3]));
   SEN_INV_2 U955 (.X(net83508), 
	.A(net83172));
   SEN_ND2_S_8 U957 (.X(n1679), 
	.A2(n1677), 
	.A1(net85815));
   SEN_OAI21_S_8 U958 (.X(n1473), 
	.B(n1407), 
	.A2(n1408), 
	.A1(n1409));
   SEN_OA2BB2_4 U959 (.X(net82074), 
	.B2(net82078), 
	.B1(net82077), 
	.A2(net82076), 
	.A1(net82075));
   SEN_AOAI211_8 U960 (.X(n1705), 
	.C(n1639), 
	.B(n1640), 
	.A2(n1641), 
	.A1(n1642));
   SEN_ND2_T_4 U961 (.X(net82839), 
	.A2(n1456), 
	.A1(n1457));
   SEN_ND2_3 U962 (.X(net84366), 
	.A2(n867), 
	.A1(n868));
   SEN_NR2_T_8 U963 (.X(n1625), 
	.A2(n1622), 
	.A1(n240));
   SEN_OAI21_T_3 U964 (.X(n225), 
	.B(n220), 
	.A2(n126), 
	.A1(net85351));
   SEN_EN2_5 U965 (.X(net83309), 
	.A2(n225), 
	.A1(n224));
   SEN_OAI21_T_3 U966 (.X(net82186), 
	.B(net82190), 
	.A2(net82189), 
	.A1(net82188));
   SEN_EO2_5 U967 (.X(net82636), 
	.A2(n1531), 
	.A1(n1532));
   SEN_AOI21_G_4 U968 (.X(n1531), 
	.B(n1529), 
	.A2(n1578), 
	.A1(n1530));
   SEN_EN2_S_3 U969 (.X(net83163), 
	.A2(n1288), 
	.A1(n375));
   SEN_EN2_S_6 U970 (.X(net83164), 
	.A2(n460), 
	.A1(n459));
   SEN_AO21B_4 U971 (.X(n460), 
	.B(n1293), 
	.A2(n1294), 
	.A1(net86332));
   SEN_AOAI211_6 U972 (.X(net82251), 
	.C(n1761), 
	.B(n1762), 
	.A2(n1763), 
	.A1(n1764));
   SEN_EN3_6 U973 (.X(n1647), 
	.A3(n1642), 
	.A2(n1641), 
	.A1(n1640));
   SEN_ND2B_V1_3 U974 (.X(n1158), 
	.B(net83829), 
	.A(C[14]));
   SEN_EN2_S_2 U975 (.X(net83206), 
	.A2(net83164), 
	.A1(net83163));
   SEN_ND2_T_4 U976 (.X(n1163), 
	.A2(n595), 
	.A1(n594));
   SEN_ND2_4 U977 (.X(n595), 
	.A2(n1117), 
	.A1(n592));
   SEN_AN3B_8 U978 (.X(n1447), 
	.B2(n1437), 
	.B1(n1438), 
	.A(net82970));
   SEN_EO3_3 U979 (.X(n897), 
	.A3(n901), 
	.A2(n550), 
	.A1(net84217));
   SEN_EN2_S_6 U980 (.X(net82387), 
	.A2(n1805), 
	.A1(n1738));
   SEN_EO2_5 U981 (.X(n1574), 
	.A2(net95993), 
	.A1(n1515));
   SEN_AOI21_S_4 U982 (.X(n1515), 
	.B(net82798), 
	.A2(n1565), 
	.A1(n1514));
   SEN_ND2B_S_4 U983 (.X(net82845), 
	.B(n1398), 
	.A(net83064));
   SEN_ND2_T_8 U984 (.X(net85071), 
	.A2(net83385), 
	.A1(net83387));
   SEN_AO21B_1 U985 (.X(n699), 
	.B(net84186), 
	.A2(net84193), 
	.A1(net84217));
   SEN_EO2_G_8 U987 (.X(n1129), 
	.A2(n1092), 
	.A1(n1093));
   SEN_EO2_8 U988 (.X(net82084), 
	.A2(n1810), 
	.A1(n1811));
   SEN_ND2_S_8 U989 (.X(net94287), 
	.A2(pprow0_qual[1]), 
	.A1(net84734));
   SEN_AN3_4 U990 (.X(net83689), 
	.A3(net83582), 
	.A2(net86258), 
	.A1(net86257));
   SEN_ND2_T_1 U991 (.X(n430), 
	.A2(net83572), 
	.A1(net83571));
   SEN_EO2_8 U993 (.X(net83953), 
	.A2(n753), 
	.A1(n752));
   SEN_AO31_4 U994 (.X(n753), 
	.B(net83960), 
	.A3(net83887), 
	.A2(net83998), 
	.A1(net83559));
   SEN_INV_1P25 U995 (.X(n1156), 
	.A(n778));
   SEN_ND2B_V1_4 U996 (.X(n1280), 
	.B(n1246), 
	.A(pprow1_qual[16]));
   SEN_INV_S_3 U997 (.X(n1246), 
	.A(pprow1_qual[14]));
   SEN_EO2_3 U998 (.X(net90316), 
	.A2(net86493), 
	.A1(net82063));
   SEN_EN2_DG_4 U999 (.X(n250), 
	.A2(n2101), 
	.A1(net82595));
   SEN_ND2_T_8 U1000 (.X(net84391), 
	.A2(net84350), 
	.A1(net84395));
   SEN_OA21_4 U1001 (.X(n1026), 
	.B(n1156), 
	.A2(net85334), 
	.A1(net84028));
   SEN_EO2_6 U1002 (.X(net83540), 
	.A2(n1181), 
	.A1(n1182));
   SEN_EO2_1 U1003 (.X(n389), 
	.A2(n244), 
	.A1(net83540));
   SEN_AOI21_S_1 U1004 (.X(net84405), 
	.B(net84425), 
	.A2(n84), 
	.A1(net84366));
   SEN_EO2_8 U1006 (.X(n1604), 
	.A2(n652), 
	.A1(n433));
   SEN_AO31_4 U1007 (.X(n652), 
	.B(n1551), 
	.A3(net82736), 
	.A2(n1552), 
	.A1(net82734));
   SEN_ND2_G_4 U1008 (.X(net83170), 
	.A2(net90814), 
	.A1(net83171));
   SEN_OAI21B_3 U1009 (.X(net82426), 
	.B(net86518), 
	.A2(net82634), 
	.A1(net90668));
   SEN_EO2_5 U1010 (.X(n1614), 
	.A2(n735), 
	.A1(n1608));
   SEN_ND2_S_3 U1011 (.X(n492), 
	.A2(net82197), 
	.A1(net82196));
   SEN_INV_S_3 U1012 (.X(net83684), 
	.A(net83679));
   SEN_ND2B_S_8 U1013 (.X(n563), 
	.B(net86213), 
	.A(net85173));
   SEN_INV_1P5 U1014 (.X(n1310), 
	.A(n1313));
   SEN_OR2_2P5 U1015 (.X(net82512), 
	.A2(net87101), 
	.A1(net87100));
   SEN_EN2_S_6 U1017 (.X(net84274), 
	.A2(n446), 
	.A1(n374));
   SEN_EN2_8 U1018 (.X(net82183), 
	.A2(net82055), 
	.A1(net82057));
   SEN_EO3_6 U1019 (.X(n1596), 
	.A3(n1599), 
	.A2(n561), 
	.A1(n2052));
   SEN_ND2_G_4 U1020 (.X(n1595), 
	.A2(net82745), 
	.A1(n1548));
   SEN_ND2_8 U1021 (.X(net82058), 
	.A2(net82335), 
	.A1(net82336));
   SEN_ND2_T_1 U1022 (.X(net82067), 
	.A2(net82069), 
	.A1(net82068));
   SEN_INV_S_4 U1024 (.X(net83648), 
	.A(net83527));
   SEN_INV_4 U1025 (.X(n1398), 
	.A(n1397));
   SEN_EO2_8 U1026 (.X(n1397), 
	.A2(n466), 
	.A1(n465));
   SEN_AO21B_6 U1027 (.X(n466), 
	.B(net83103), 
	.A2(net83098), 
	.A1(net83209));
   SEN_BUF_S_6 U1028 (.X(net95748), 
	.A(net84000));
   SEN_INV_S_6 U1029 (.X(net83999), 
	.A(net84002));
   SEN_INV_S_3 U1030 (.X(net87101), 
	.A(net82197));
   SEN_ND2_T_1 U1031 (.X(n594), 
	.A2(n593), 
	.A1(n1118));
   SEN_EN3_DG_8 U1032 (.X(net82462), 
	.A3(pprow0_qual[27]), 
	.A2(n1703), 
	.A1(n1705));
   SEN_EN2_S_2 U1033 (.X(n666), 
	.A2(n1604), 
	.A1(n1602));
   SEN_AO21B_8 U1034 (.X(n468), 
	.B(n469), 
	.A2(n474), 
	.A1(net86477));
   SEN_INV_4 U1036 (.X(n90), 
	.A(n1700));
   SEN_INV_5 U1037 (.X(n1700), 
	.A(n1646));
   SEN_ND2_S_6 U1038 (.X(n1699), 
	.A2(net82467), 
	.A1(net82466));
   SEN_AN2_3 U1039 (.X(n93), 
	.A2(net83582), 
	.A1(net86258));
   SEN_ND2_T_1P5 U1040 (.X(net87769), 
	.A2(n93), 
	.A1(net86257));
   SEN_ND2_G_3 U1041 (.X(net83582), 
	.A2(pprow3_qual[7]), 
	.A1(pprow2_qual[9]));
   SEN_OAI21_S_3 U1042 (.X(n1272), 
	.B(n1190), 
	.A2(n1191), 
	.A1(n1152));
   SEN_ND2_T_2 U1043 (.X(n1274), 
	.A2(n1203), 
	.A1(n1246));
   SEN_ND2_G_1 U1044 (.X(n526), 
	.A2(n1153), 
	.A1(n1223));
   SEN_ND2_2 U1046 (.X(n95), 
	.A2(n1001), 
	.A1(n925));
   SEN_ND2_3 U1047 (.X(n1003), 
	.A2(n96), 
	.A1(n926));
   SEN_INV_S_3 U1048 (.X(n96), 
	.A(n95));
   SEN_ND2_3 U1049 (.X(n925), 
	.A2(pprow1_qual[2]), 
	.A1(pprow1_qual[4]));
   SEN_AN3_4 U1051 (.X(n1005), 
	.A3(n769), 
	.A2(n1003), 
	.A1(n558));
   SEN_ND3_2 U1052 (.X(n968), 
	.A3(n999), 
	.A2(n927), 
	.A1(n1003));
   SEN_NR2_T_1 U1053 (.X(n97), 
	.A2(n1284), 
	.A1(n1357));
   SEN_NR2_T_1 U1054 (.X(n1286), 
	.A2(n98), 
	.A1(n1285));
   SEN_INV_S_2 U1055 (.X(n98), 
	.A(n97));
   SEN_ND2_1P5 U1056 (.X(net82743), 
	.A2(net82878), 
	.A1(n99));
   SEN_EO2_2 U1057 (.X(net82876), 
	.A2(n346), 
	.A1(n112));
   SEN_ND2_1 U1058 (.X(n101), 
	.A2(pprow3_qual[9]), 
	.A1(pprow2_qual[11]));
   SEN_INV_2 U1059 (.X(n102), 
	.A(n424));
   SEN_AN3_4 U1060 (.X(net85351), 
	.A3(n102), 
	.A2(n101), 
	.A1(n100));
   SEN_AOI31_3 U1062 (.X(n424), 
	.B(n428), 
	.A3(n425), 
	.A2(n426), 
	.A1(n427));
   SEN_EO2_3 U1063 (.X(net83461), 
	.A2(net85351), 
	.A1(n223));
   SEN_INV_S_4 U1065 (.X(net95559), 
	.A(net83077));
   SEN_OR3B_2 U1066 (.X(n1454), 
	.B2(n1449), 
	.B1(n1448), 
	.A(n1452));
   SEN_AN2_S_0P5 U1067 (.X(n120), 
	.A2(net82965), 
	.A1(net82967));
   SEN_INV_8 U1068 (.X(n1068), 
	.A(n1066));
   SEN_ND3_T_1P5 U1069 (.X(n1023), 
	.A3(n702), 
	.A2(n1147), 
	.A1(n1149));
   SEN_ND2_8 U1070 (.X(net83552), 
	.A2(net83954), 
	.A1(net83953));
   SEN_ND2_T_2 U1071 (.X(n1112), 
	.A2(n1149), 
	.A1(n702));
   SEN_ND2_T_1P5 U1072 (.X(net84437), 
	.A2(net84417), 
	.A1(net84392));
   SEN_AOI21_3 U1073 (.X(n1577), 
	.B(n1575), 
	.A2(n1619), 
	.A1(n1576));
   SEN_ND2_T_3 U1074 (.X(n1576), 
	.A2(n1620), 
	.A1(n781));
   SEN_EO2_S_1 U1075 (.X(n1716), 
	.A2(net86491), 
	.A1(net82323));
   SEN_INV_S_6 U1076 (.X(net83733), 
	.A(net83645));
   SEN_INV_3 U1077 (.X(net87541), 
	.A(net86494));
   SEN_ND2_T_2 U1078 (.X(net87543), 
	.A2(net86494), 
	.A1(net82062));
   SEN_EO2_4 U1080 (.X(n1328), 
	.A2(n1295), 
	.A1(net83152));
   SEN_EO2_2 U1081 (.X(n682), 
	.A2(net82717), 
	.A1(n1561));
   SEN_INV_S_6 U1082 (.X(net82285), 
	.A(net82332));
   SEN_AN2_6 U1083 (.X(net86333), 
	.A2(net83304), 
	.A1(net83301));
   SEN_ND2_3 U1084 (.X(n1772), 
	.A2(net82285), 
	.A1(net82284));
   SEN_EO2_2 U1085 (.X(n457), 
	.A2(net83455), 
	.A1(net83454));
   SEN_ND2_G_3 U1086 (.X(n1675), 
	.A2(n590), 
	.A1(n589));
   SEN_ND2_2 U1087 (.X(n590), 
	.A2(n463), 
	.A1(n587));
   SEN_ND2_4 U1088 (.X(net82195), 
	.A2(net82387), 
	.A1(net82386));
   SEN_INV_S_6 U1089 (.X(n882), 
	.A(n880));
   SEN_ND2_4 U1090 (.X(net83414), 
	.A2(n574), 
	.A1(n573));
   SEN_EO2_G_8 U1091 (.X(net83845), 
	.A2(net83933), 
	.A1(n1064));
   SEN_BUF_S_3 U1092 (.X(n467), 
	.A(net83723));
   SEN_INV_3 U1093 (.X(n1421), 
	.A(n1422));
   SEN_EN2_S_2 U1094 (.X(n1422), 
	.A2(n562), 
	.A1(n680));
   SEN_EN2_5 U1095 (.X(n1587), 
	.A2(n1576), 
	.A1(n1525));
   SEN_ND2_S_3 U1096 (.X(net82187), 
	.A2(net82189), 
	.A1(net82188));
   SEN_EO2_2 U1098 (.X(n517), 
	.A2(net82251), 
	.A1(n116));
   SEN_INV_S_3 U1099 (.X(net82420), 
	.A(n155));
   SEN_EO2_S_3 U1100 (.X(net83723), 
	.A2(n1114), 
	.A1(n1115));
   SEN_OAOI211_4 U1101 (.X(n1114), 
	.C(n1110), 
	.B(n1111), 
	.A2(n1112), 
	.A1(n1113));
   SEN_ND2B_6 U1102 (.X(net84111), 
	.B(net85173), 
	.A(net83833));
   SEN_AOI21_S_4 U1103 (.X(n197), 
	.B(n188), 
	.A2(net83965), 
	.A1(n192));
   SEN_NR2_S_2 U1104 (.X(n192), 
	.A2(net84001), 
	.A1(net83999));
   SEN_NR2_G_2 U1105 (.X(n775), 
	.A2(n1739), 
	.A1(n1740));
   SEN_ND2_S_3 U1106 (.X(net82280), 
	.A2(n1739), 
	.A1(n1740));
   SEN_ND2B_6 U1107 (.X(n1018), 
	.B(n956), 
	.A(n957));
   SEN_EO2_S_3 U1108 (.X(net82063), 
	.A2(net82061), 
	.A1(net82060));
   SEN_OAI21_S_8 U1109 (.X(n1770), 
	.B(net82280), 
	.A2(n1769), 
	.A1(n775));
   SEN_EN2_1 U1111 (.X(n1532), 
	.A2(n1587), 
	.A1(n1588));
   SEN_NR2_T_2 U1112 (.X(net88103), 
	.A2(net82831), 
	.A1(net94176));
   SEN_AO21B_4 U1113 (.X(n1550), 
	.B(n1595), 
	.A2(n1593), 
	.A1(net82743));
   SEN_INV_1P5 U1114 (.X(net82066), 
	.A(net82068));
   SEN_EO2_S_6 U1115 (.X(net86494), 
	.A2(net82068), 
	.A1(net82059));
   SEN_INV_S_2 U1116 (.X(n494), 
	.A(net82236));
   SEN_ND2_S_2 U1117 (.X(net87813), 
	.A2(n625), 
	.A1(n1530));
   SEN_INV_S_2 U1118 (.X(n624), 
	.A(n1530));
   SEN_EO2_3 U1119 (.X(n956), 
	.A2(n738), 
	.A1(n737));
   SEN_AO21B_2 U1120 (.X(n738), 
	.B(n965), 
	.A2(n558), 
	.A1(n943));
   SEN_INV_4 U1121 (.X(n323), 
	.A(net83844));
   SEN_INV_2 U1122 (.X(n1457), 
	.A(n1460));
   SEN_ND2_S_4 U1123 (.X(net82842), 
	.A2(net82934), 
	.A1(n1460));
   SEN_EO2_1 U1124 (.X(n1412), 
	.A2(n1410), 
	.A1(n740));
   SEN_OAI21_3 U1125 (.X(n1224), 
	.B(n1270), 
	.A2(n1249), 
	.A1(n1204));
   SEN_EO2_2 U1126 (.X(n1651), 
	.A2(n1643), 
	.A1(net82550));
   SEN_EN2_6 U1127 (.X(n1297), 
	.A2(n627), 
	.A1(n546));
   SEN_EN2_DG_2 U1128 (.X(n546), 
	.A2(pprow7_qual[3]), 
	.A1(pprow6_qual[5]));
   SEN_INV_1P25 U1129 (.X(n535), 
	.A(n867));
   SEN_INV_3 U1130 (.X(net84352), 
	.A(net84355));
   SEN_ND2_T_2 U1131 (.X(net84355), 
	.A2(pprow0_qual[5]), 
	.A1(C[5]));
   SEN_OAI21_3 U1132 (.X(net82587), 
	.B(n1578), 
	.A2(n1588), 
	.A1(n1587));
   SEN_INV_2 U1133 (.X(net82390), 
	.A(net82387));
   SEN_EN2_S_3 U1134 (.X(net86534), 
	.A2(net82389), 
	.A1(net82387));
   SEN_INV_3 U1136 (.X(net83964), 
	.A(net83786));
   SEN_BUF_1 U1137 (.X(n478), 
	.A(net83454));
   SEN_AOAI211_8 U1138 (.X(net91024), 
	.C(n1806), 
	.B(n1807), 
	.A2(net82203), 
	.A1(net82202));
   SEN_NR2_S_0P8 U1139 (.X(n1177), 
	.A2(pprow4_qual[6]), 
	.A1(pprow5_qual[4]));
   SEN_ND2_T_5 U1141 (.X(net82196), 
	.A2(net82514), 
	.A1(net82513));
   SEN_EO2_4 U1142 (.X(n1019), 
	.A2(n721), 
	.A1(n1023));
   SEN_AN4B_1 U1143 (.X(n1287), 
	.B3(n1359), 
	.B2(net83192), 
	.B1(n1358), 
	.A(n1286));
   SEN_ND2B_V1_1 U1144 (.X(n329), 
	.B(net83090), 
	.A(n328));
   SEN_EO2_1 U1145 (.X(n939), 
	.A2(net85984), 
	.A1(n741));
   SEN_ND2B_V1_4 U1146 (.X(net83610), 
	.B(n1188), 
	.A(n1187));
   SEN_ND2_4 U1147 (.X(net82843), 
	.A2(n1397), 
	.A1(net83064));
   SEN_ND2_T_4 U1149 (.X(net84228), 
	.A2(net84159), 
	.A1(net86078));
   SEN_AO21B_6 U1150 (.X(net82385), 
	.B(net82196), 
	.A2(net82193), 
	.A1(net82512));
   SEN_INV_S_1 U1151 (.X(net82674), 
	.A(net82587));
   SEN_EO2_8 U1152 (.X(net91053), 
	.A2(n1553), 
	.A1(n666));
   SEN_OAI21_S_3 U1153 (.X(n1141), 
	.B(n38), 
	.A2(n1138), 
	.A1(n1139));
   SEN_OAI21_S_8 U1154 (.X(n353), 
	.B(n347), 
	.A2(n345), 
	.A1(net98293));
   SEN_EN2_S_3 U1155 (.X(n664), 
	.A2(n1672), 
	.A1(net82499));
   SEN_INV_3 U1156 (.X(n1672), 
	.A(n1675));
   SEN_NR2_S_2 U1157 (.X(n1288), 
	.A2(net83197), 
	.A1(n1287));
   SEN_EO2_S_3 U1158 (.X(n522), 
	.A2(n1486), 
	.A1(n1487));
   SEN_ND2_S_1P5 U1159 (.X(n514), 
	.A2(n523), 
	.A1(n1282));
   SEN_ND2_2 U1160 (.X(n1282), 
	.A2(n1005), 
	.A1(n1006));
   SEN_INV_5 U1161 (.X(n995), 
	.A(n1004));
   SEN_INV_S_4 U1162 (.X(n1089), 
	.A(pprow2_qual[7]));
   SEN_EO2_8 U1163 (.X(n1327), 
	.A2(n1323), 
	.A1(net83214));
   SEN_ND2_6 U1164 (.X(net83214), 
	.A2(n473), 
	.A1(net86477));
   SEN_EO2_S_3 U1165 (.X(n1069), 
	.A2(n1024), 
	.A1(n1025));
   SEN_AOI21B_2 U1166 (.X(n1024), 
	.B(n1148), 
	.A2(n545), 
	.A1(n1023));
   SEN_EN2_S_2 U1167 (.X(n1100), 
	.A2(net87790), 
	.A1(net83681));
   SEN_OAI211_2 U1168 (.X(n943), 
	.B2(n966), 
	.B1(n968), 
	.A2(n963), 
	.A1(n998));
   SEN_OA21_2 U1169 (.X(n103), 
	.B(net82460), 
	.A2(n1702), 
	.A1(n1701));
   SEN_INV_4 U1170 (.X(net82523), 
	.A(net82520));
   SEN_EO2_S_3 U1171 (.X(net82520), 
	.A2(net86455), 
	.A1(net86454));
   SEN_NR3_T_6 U1172 (.X(n1363), 
	.A3(net83197), 
	.A2(n1355), 
	.A1(n1356));
   SEN_ND2_T_1P5 U1173 (.X(n1355), 
	.A2(n1283), 
	.A1(n1282));
   SEN_OAI21_5 U1175 (.X(net82075), 
	.B(net82187), 
	.A2(net82186), 
	.A1(n491));
   SEN_OAOI211_4 U1176 (.X(n491), 
	.C(net82194), 
	.B(net82193), 
	.A2(n492), 
	.A1(net87100));
   SEN_INV_4 U1177 (.X(n881), 
	.A(n246));
   SEN_EO2_2 U1178 (.X(n246), 
	.A2(n871), 
	.A1(n247));
   SEN_INV_1 U1179 (.X(n868), 
	.A(n539));
   SEN_ND2_S_4 U1180 (.X(net84378), 
	.A2(n535), 
	.A1(n539));
   SEN_EO2_2 U1181 (.X(n539), 
	.A2(n863), 
	.A1(n865));
   SEN_EO2_G_4 U1182 (.X(net83678), 
	.A2(n1140), 
	.A1(n1141));
   SEN_AN2_2 U1183 (.X(net86385), 
	.A2(net87790), 
	.A1(net83681));
   SEN_INV_4 U1184 (.X(n363), 
	.A(net82347));
   SEN_EN3_6 U1185 (.X(net82347), 
	.A3(n1764), 
	.A2(n1763), 
	.A1(n1762));
   SEN_INV_S_3 U1186 (.X(n1572), 
	.A(n1573));
   SEN_EO2_8 U1188 (.X(net82068), 
	.A2(net82241), 
	.A1(net82183));
   SEN_ND2_0P5 U1189 (.X(n1389), 
	.A2(pprow5_qual[9]), 
	.A1(pprow4_qual[11]));
   SEN_ND2_2 U1190 (.X(n1360), 
	.A2(n529), 
	.A1(n1358));
   SEN_AN2_5 U1191 (.X(n529), 
	.A2(net83192), 
	.A1(n1359));
   SEN_ND2_S_0P5 U1192 (.X(n1374), 
	.A2(pprow7_qual[5]), 
	.A1(pprow6_qual[7]));
   SEN_OR2_1 U1193 (.X(n750), 
	.A2(pprow6_qual[7]), 
	.A1(pprow7_qual[5]));
   SEN_ND2_S_4 U1194 (.X(n441), 
	.A2(net83171), 
	.A1(net82980));
   SEN_AOAI211_3 U1195 (.X(n1765), 
	.C(n1712), 
	.B(n1713), 
	.A2(n1714), 
	.A1(net82436));
   SEN_INV_3 U1197 (.X(n1353), 
	.A(n1284));
   SEN_ND2_G_0P65 U1198 (.X(n1477), 
	.A2(pprow5_qual[11]), 
	.A1(pprow4_qual[13]));
   SEN_ND2_S_0P5 U1200 (.X(n371), 
	.A2(net91392), 
	.A1(net82562));
   SEN_INV_1P25 U1201 (.X(net91392), 
	.A(pprow1_qual[24]));
   SEN_ND2_G_1 U1202 (.X(n966), 
	.A2(pprow1_qual[4]), 
	.A1(pprow1_qual[6]));
   SEN_ND2_2 U1203 (.X(net84073), 
	.A2(net84007), 
	.A1(net86076));
   SEN_ND2_S_0P65 U1204 (.X(n220), 
	.A2(pprow2_qual[12]), 
	.A1(pprow3_qual[10]));
   SEN_INV_1 U1205 (.X(n216), 
	.A(pprow3_qual[10]));
   SEN_INV_1 U1206 (.X(n215), 
	.A(pprow2_qual[12]));
   SEN_AOI32_1 U1207 (.X(n1276), 
	.B2(n557), 
	.B1(n1273), 
	.A3(n1275), 
	.A2(n1274), 
	.A1(n537));
   SEN_NR2_G_3 U1208 (.X(n1385), 
	.A2(n1380), 
	.A1(n1381));
   SEN_NR2_T_1 U1209 (.X(n1381), 
	.A2(n1387), 
	.A1(n1386));
   SEN_EO2_S_3 U1210 (.X(net82741), 
	.A2(n336), 
	.A1(n113));
   SEN_INV_S_1 U1211 (.X(n1559), 
	.A(pprow8_qual[7]));
   SEN_INV_S_1 U1212 (.X(n1558), 
	.A(pprow9_qual[5]));
   SEN_INV_S_0P5 U1213 (.X(net91390), 
	.A(pprow1_qual[26]));
   SEN_ND2_S_0P5 U1214 (.X(net91419), 
	.A2(pprow1_qual[24]), 
	.A1(pprow1_qual[26]));
   SEN_EO2_1 U1215 (.X(n106), 
	.A2(net84730), 
	.A1(n449));
   SEN_NR2_S_2 U1216 (.X(n778), 
	.A2(pprow0_qual[12]), 
	.A1(C[12]));
   SEN_ND3_T_2 U1218 (.X(n1357), 
	.A3(n1270), 
	.A2(n1247), 
	.A1(n1202));
   SEN_INV_S_3 U1219 (.X(n1689), 
	.A(n1633));
   SEN_AOAI211_3 U1220 (.X(n1633), 
	.C(n1629), 
	.B(n1630), 
	.A2(n1631), 
	.A1(n1632));
   SEN_OA2BB2_4 U1223 (.X(n1678), 
	.B2(net85815), 
	.B1(n1677), 
	.A2(n700), 
	.A1(n1679));
   SEN_EN2_S_2 U1224 (.X(n1723), 
	.A2(net82420), 
	.A1(n1685));
   SEN_EO2_S_0P5 U1225 (.X(n729), 
	.A2(n528), 
	.A1(n533));
   SEN_NR2_T_1P5 U1226 (.X(net82244), 
	.A2(net82246), 
	.A1(net82247));
   SEN_EO2_1 U1227 (.X(net82246), 
	.A2(n366), 
	.A1(net82248));
   SEN_ND2B_V1_4 U1228 (.X(n1208), 
	.B(n1164), 
	.A(n236));
   SEN_INV_S_3 U1229 (.X(n1164), 
	.A(n1163));
   SEN_INV_1P5 U1231 (.X(n188), 
	.A(net83578));
   SEN_INV_S_0P5 U1232 (.X(n335), 
	.A(pprow1_qual[21]));
   SEN_ND2_T_1P5 U1233 (.X(n1132), 
	.A2(net83581), 
	.A1(net83890));
   SEN_OR2_2 U1234 (.X(net83577), 
	.A2(pprow3_qual[7]), 
	.A1(pprow2_qual[9]));
   SEN_INV_S_3 U1235 (.X(net83573), 
	.A(net83891));
   SEN_ND2_2 U1236 (.X(n1313), 
	.A2(pprow5_qual[6]), 
	.A1(pprow4_qual[8]));
   SEN_ND2_2 U1237 (.X(n1284), 
	.A2(n1279), 
	.A1(n1278));
   SEN_ND2B_V1_2 U1238 (.X(n1428), 
	.B(n1424), 
	.A(C[22]));
   SEN_INV_S_1P5 U1239 (.X(n328), 
	.A(pprow1_qual[17]));
   SEN_ND2_T_1 U1240 (.X(n1543), 
	.A2(C[23]), 
	.A1(pprow0_qual[23]));
   SEN_INV_S_1 U1241 (.X(n138), 
	.A(pprow6_qual[11]));
   SEN_INV_S_0P5 U1242 (.X(net91386), 
	.A(pprow1_qual[25]));
   SEN_ND2_T_1P5 U1243 (.X(n1150), 
	.A2(n1107), 
	.A1(n1108));
   SEN_ND2_G_1 U1244 (.X(n1108), 
	.A2(n1022), 
	.A1(n1109));
   SEN_ND2_S_4 U1245 (.X(n1198), 
	.A2(n1008), 
	.A1(n999));
   SEN_INV_S_1 U1246 (.X(n1293), 
	.A(n1368));
   SEN_ND2_1P5 U1247 (.X(net83192), 
	.A2(net83359), 
	.A1(n328));
   SEN_ND2B_V1_2 U1248 (.X(n1429), 
	.B(n1392), 
	.A(C[21]));
   SEN_INV_1P5 U1249 (.X(n397), 
	.A(n1357));
   SEN_ND2_2 U1250 (.X(n646), 
	.A2(n1483), 
	.A1(n1482));
   SEN_OR2_1 U1251 (.X(n245), 
	.A2(n1484), 
	.A1(net82889));
   SEN_ND2_8 U1253 (.X(n1514), 
	.A2(n1479), 
	.A1(net82899));
   SEN_NR2_1 U1254 (.X(n1479), 
	.A2(net82903), 
	.A1(net82902));
   SEN_NR2B_1 U1255 (.X(net82902), 
	.B(n401), 
	.A(n109));
   SEN_EO2_S_0P5 U1256 (.X(n742), 
	.A2(pprow5_qual[15]), 
	.A1(pprow4_qual[17]));
   SEN_NR2_S_0P5 U1258 (.X(n368), 
	.A2(pprow1_qual[24]), 
	.A1(pprow1_qual[26]));
   SEN_INV_3 U1260 (.X(n549), 
	.A(n548));
   SEN_NR2_S_5 U1261 (.X(n548), 
	.A2(n1697), 
	.A1(n698));
   SEN_EN2_0P5 U1262 (.X(n743), 
	.A2(pprow13_qual[1]), 
	.A1(pprow12_qual[3]));
   SEN_OAI21_5 U1263 (.X(n566), 
	.B(net84410), 
	.A2(net94287), 
	.A1(net84450));
   SEN_EN2_S_1 U1265 (.X(n374), 
	.A2(n387), 
	.A1(net84288));
   SEN_INV_S_4 U1266 (.X(n1022), 
	.A(pprow1_qual[8]));
   SEN_ND2_T_2 U1267 (.X(n1107), 
	.A2(n1153), 
	.A1(n1058));
   SEN_ND2_T_4 U1268 (.X(n1083), 
	.A2(pprow5_qual[0]), 
	.A1(pprow4_qual[2]));
   SEN_EO2_3 U1269 (.X(net83875), 
	.A2(n1011), 
	.A1(n709));
   SEN_ND2_S_3 U1270 (.X(n1192), 
	.A2(n1148), 
	.A1(n1149));
   SEN_ND2B_V1_3 U1271 (.X(n1255), 
	.B(net83435), 
	.A(C[18]));
   SEN_ND2_T_1 U1272 (.X(n1290), 
	.A2(n1255), 
	.A1(net83434));
   SEN_INV_S_0P5 U1273 (.X(n229), 
	.A(net83114));
   SEN_ND2_0P5 U1274 (.X(n382), 
	.A2(pprow5_qual[8]), 
	.A1(pprow4_qual[10]));
   SEN_OR2_1 U1275 (.X(n381), 
	.A2(pprow4_qual[10]), 
	.A1(pprow5_qual[8]));
   SEN_ND2_S_3 U1276 (.X(net83114), 
	.A2(n213), 
	.A1(n212));
   SEN_INV_2 U1277 (.X(n212), 
	.A(pprow2_qual[14]));
   SEN_INV_S_2 U1278 (.X(n213), 
	.A(pprow3_qual[12]));
   SEN_NR2B_V1_1 U1279 (.X(n219), 
	.B(n217), 
	.A(pprow3_qual[11]));
   SEN_ND2_S_0P5 U1280 (.X(net83111), 
	.A2(pprow3_qual[12]), 
	.A1(pprow2_qual[14]));
   SEN_INV_2 U1281 (.X(n627), 
	.A(n1338));
   SEN_OR2_1 U1282 (.X(n532), 
	.A2(pprow6_qual[8]), 
	.A1(pprow7_qual[6]));
   SEN_EO2_S_0P5 U1283 (.X(n715), 
	.A2(pprow7_qual[6]), 
	.A1(pprow6_qual[8]));
   SEN_INV_1 U1284 (.X(n1416), 
	.A(n1412));
   SEN_EN2_0P5 U1285 (.X(n1631), 
	.A2(n816), 
	.A1(pprow12_qual[0]));
   SEN_OAI21_5 U1286 (.X(n1612), 
	.B(n1562), 
	.A2(n602), 
	.A1(n1563));
   SEN_AOAI211_4 U1287 (.X(n1744), 
	.C(n1688), 
	.B(n1689), 
	.A2(n261), 
	.A1(n1690));
   SEN_INV_S_1 U1288 (.X(n1687), 
	.A(n1690));
   SEN_EN2_1 U1289 (.X(net82248), 
	.A2(pprow1_qual[25]), 
	.A1(pprow1_qual[27]));
   SEN_INV_S_1 U1290 (.X(n1739), 
	.A(n1741));
   SEN_INV_2 U1291 (.X(n287), 
	.A(\bmul/neg1 ));
   SEN_ND2B_2 U1292 (.X(net84414), 
	.B(n866), 
	.A(C[3]));
   SEN_ND2_T_1 U1293 (.X(n635), 
	.A2(n725), 
	.A1(n632));
   SEN_ND2_S_1 U1295 (.X(n1061), 
	.A2(n1148), 
	.A1(n1147));
   SEN_EN2_0P5 U1296 (.X(n1218), 
	.A2(n1227), 
	.A1(n2051));
   SEN_ND3_1 U1297 (.X(n1254), 
	.A3(n1250), 
	.A2(n1251), 
	.A1(n774));
   SEN_EO2_2 U1298 (.X(n1377), 
	.A2(n1373), 
	.A1(n706));
   SEN_EO2_S_0P5 U1299 (.X(n706), 
	.A2(pprow7_qual[5]), 
	.A1(pprow6_qual[7]));
   SEN_ND2_2 U1300 (.X(n1585), 
	.A2(n1528), 
	.A1(n522));
   SEN_INV_S_1 U1301 (.X(n1627), 
	.A(n1631));
   SEN_INV_S_1 U1302 (.X(n1603), 
	.A(n1602));
   SEN_ND2_S_0P8 U1303 (.X(n1656), 
	.A2(n1660), 
	.A1(n1651));
   SEN_INV_S_1 U1304 (.X(n1575), 
	.A(n1621));
   SEN_OR2_2P5 U1305 (.X(net83815), 
	.A2(n952), 
	.A1(n951));
   SEN_AOI31_2 U1306 (.X(n978), 
	.B(net84146), 
	.A3(net84116), 
	.A2(n976), 
	.A1(n977));
   SEN_INV_3 U1307 (.X(net82077), 
	.A(net82079));
   SEN_INV_2 U1308 (.X(n282), 
	.A(n286));
   SEN_EO2_1 U1309 (.X(n286), 
	.A2(net84654), 
	.A1(n284));
   SEN_INV_S_1 U1310 (.X(n284), 
	.A(pprow1_qual[0]));
   SEN_EO2_S_0P5 U1311 (.X(n234), 
	.A2(n239), 
	.A1(net83844));
   SEN_EN2_0P5 U1312 (.X(n1262), 
	.A2(net83389), 
	.A1(net83390));
   SEN_INV_4 U1313 (.X(n326), 
	.A(net82842));
   SEN_NR2_S_2 U1314 (.X(n194), 
	.A2(net84011), 
	.A1(net83999));
   SEN_INV_S_1 U1315 (.X(n332), 
	.A(pprow1_qual[18]));
   SEN_ND2_2 U1316 (.X(n621), 
	.A2(net87822), 
	.A1(net87821));
   SEN_INV_S_1 U1317 (.X(net87822), 
	.A(n445));
   SEN_INV_2 U1318 (.X(n1203), 
	.A(pprow1_qual[12]));
   SEN_EO2_S_0P5 U1319 (.X(n726), 
	.A2(pprow3_qual[8]), 
	.A1(pprow2_qual[10]));
   SEN_ND2_2 U1320 (.X(n1136), 
	.A2(pprow5_qual[2]), 
	.A1(pprow4_qual[4]));
   SEN_OR2_5 U1321 (.X(n1051), 
	.A2(pprow5_qual[1]), 
	.A1(pprow4_qual[3]));
   SEN_OR2_2 U1322 (.X(net83566), 
	.A2(pprow3_qual[9]), 
	.A1(pprow2_qual[11]));
   SEN_ND2_2 U1323 (.X(n426), 
	.A2(n431), 
	.A1(n136));
   SEN_OAI21B_2 U1324 (.X(n427), 
	.B(net83570), 
	.A2(n430), 
	.A1(n429));
   SEN_ND2_G_1 U1325 (.X(net87797), 
	.A2(n187), 
	.A1(net83574));
   SEN_INV_S_1 U1326 (.X(n187), 
	.A(n189));
   SEN_NR2B_1 U1327 (.X(n344), 
	.B(n121), 
	.A(pprow1_qual[19]));
   SEN_NR2B_1 U1328 (.X(n341), 
	.B(n121), 
	.A(pprow1_qual[17]));
   SEN_NR2_1 U1329 (.X(n342), 
	.A2(n343), 
	.A1(n121));
   SEN_ND2_G_1 U1330 (.X(n343), 
	.A2(pprow1_qual[19]), 
	.A1(pprow1_qual[17]));
   SEN_NR2B_1 U1331 (.X(n334), 
	.B(n332), 
	.A(pprow1_qual[20]));
   SEN_ND2_G_1 U1332 (.X(n1283), 
	.A2(n1201), 
	.A1(n1200));
   SEN_ND2_G_1 U1333 (.X(n1356), 
	.A2(n1353), 
	.A1(n1354));
   SEN_INV_S_1 U1334 (.X(n333), 
	.A(pprow1_qual[20]));
   SEN_INV_S_1 U1335 (.X(n340), 
	.A(net82758));
   SEN_INV_S_1 U1336 (.X(n401), 
	.A(net82701));
   SEN_NR2B_1 U1337 (.X(n402), 
	.B(n401), 
	.A(net82901));
   SEN_INV_S_1 U1338 (.X(net82903), 
	.A(net82705));
   SEN_INV_S_1 U1339 (.X(n337), 
	.A(n355));
   SEN_ND2B_1 U1340 (.X(n355), 
	.B(pprow1_qual[21]), 
	.A(n330));
   SEN_INV_2 U1341 (.X(n339), 
	.A(n354));
   SEN_ND2B_1 U1342 (.X(n1752), 
	.B(pprow12_qual[1]), 
	.A(n1637));
   SEN_ND2_G_1 U1343 (.X(n1504), 
	.A2(n1501), 
	.A1(n1502));
   SEN_ND2B_1 U1344 (.X(n141), 
	.B(n129), 
	.A(n145));
   SEN_INV_S_1 U1345 (.X(n145), 
	.A(n158));
   SEN_ND2_G_1 U1346 (.X(n418), 
	.A2(net82705), 
	.A1(net82706));
   SEN_INV_S_1 U1347 (.X(n153), 
	.A(n141));
   SEN_INV_S_1 U1348 (.X(n157), 
	.A(pprow6_qual[13]));
   SEN_INV_S_1 U1349 (.X(n156), 
	.A(pprow7_qual[11]));
   SEN_NR2_1 U1350 (.X(n147), 
	.A2(n146), 
	.A1(n127));
   SEN_NR2_1 U1351 (.X(n150), 
	.A2(n149), 
	.A1(net82721));
   SEN_NR2B_1 U1352 (.X(n149), 
	.B(n138), 
	.A(pprow7_qual[9]));
   SEN_OAI21B_4 U1353 (.X(net91408), 
	.B(n110), 
	.A2(n115), 
	.A1(net82455));
   SEN_AN2_S_1 U1354 (.X(n447), 
	.A2(n445), 
	.A1(n442));
   SEN_INV_S_1 U1355 (.X(net84288), 
	.A(pprow0_qual[8]));
   SEN_ND2_G_1 U1356 (.X(net84233), 
	.A2(net84153), 
	.A1(n443));
   SEN_ND2_2 U1357 (.X(net84150), 
	.A2(pprow0_qual[9]), 
	.A1(C[9]));
   SEN_INV_2 U1358 (.X(n942), 
	.A(pprow1_qual[5]));
   SEN_INV_3 U1359 (.X(n997), 
	.A(pprow1_qual[7]));
   SEN_BUF_S_1 U1360 (.X(n616), 
	.A(n1001));
   SEN_INV_S_1 U1361 (.X(n924), 
	.A(n906));
   SEN_INV_3 U1362 (.X(n1058), 
	.A(pprow1_qual[9]));
   SEN_INV_3 U1363 (.X(net83580), 
	.A(net83890));
   SEN_OAI21_S_2 U1364 (.X(net83960), 
	.B(net83574), 
	.A2(net83578), 
	.A1(net83580));
   SEN_ND2_2 U1366 (.X(net83570), 
	.A2(net83577), 
	.A1(net83581));
   SEN_NR2B_2 U1367 (.X(n185), 
	.B(net83578), 
	.A(net83890));
   SEN_INV_S_1 U1368 (.X(n638), 
	.A(n726));
   SEN_NR2_2 U1369 (.X(net83790), 
	.A2(n2045), 
	.A1(net86385));
   SEN_INV_S_1 U1370 (.X(n264), 
	.A(n483));
   SEN_ND2_G_3 U1371 (.X(n1196), 
	.A2(n996), 
	.A1(n1007));
   SEN_INV_S_1 U1372 (.X(n1223), 
	.A(pprow1_qual[13]));
   SEN_INV_S_1 U1373 (.X(n217), 
	.A(pprow2_qual[13]));
   SEN_INV_S_1 U1374 (.X(n222), 
	.A(n233));
   SEN_ND2_G_1 U1375 (.X(n233), 
	.A2(n217), 
	.A1(n218));
   SEN_INV_S_1 U1376 (.X(n218), 
	.A(pprow3_qual[11]));
   SEN_NR2_1 U1377 (.X(n221), 
	.A2(n220), 
	.A1(n222));
   SEN_ND2_G_1 U1378 (.X(n1314), 
	.A2(n1239), 
	.A1(n1240));
   SEN_EN2_0P5 U1379 (.X(n223), 
	.A2(pprow2_qual[12]), 
	.A1(pprow3_qual[10]));
   SEN_INV_S_1 U1380 (.X(n1301), 
	.A(pprow7_qual[3]));
   SEN_ND2_G_1 U1381 (.X(n1337), 
	.A2(pprow7_qual[3]), 
	.A1(pprow6_qual[5]));
   SEN_NR2_4 U1382 (.X(n644), 
	.A2(net83036), 
	.A1(n1478));
   SEN_ND2_G_1 U1383 (.X(n1411), 
	.A2(pprow5_qual[10]), 
	.A1(pprow4_qual[12]));
   SEN_EO2_S_0P5 U1384 (.X(n740), 
	.A2(pprow5_qual[10]), 
	.A1(pprow4_qual[12]));
   SEN_OR2_2P5 U1385 (.X(net82878), 
	.A2(net82982), 
	.A1(net82981));
   SEN_NR2_1 U1386 (.X(n347), 
	.A2(n342), 
	.A1(n334));
   SEN_NR2_1 U1387 (.X(n345), 
	.A2(n344), 
	.A1(n341));
   SEN_INV_S_1 U1388 (.X(n1424), 
	.A(pprow0_qual[22]));
   SEN_INV_S_1 U1389 (.X(n330), 
	.A(pprow1_qual[19]));
   SEN_NR2_1 U1390 (.X(n1544), 
	.A2(n1543), 
	.A1(n1546));
   SEN_INV_S_1 U1391 (.X(n1546), 
	.A(n1542));
   SEN_INV_S_1 U1392 (.X(net82798), 
	.A(net82706));
   SEN_INV_S_1 U1393 (.X(n406), 
	.A(pprow3_qual[17]));
   SEN_INV_S_1 U1394 (.X(n407), 
	.A(pprow2_qual[19]));
   SEN_EO2_3 U1395 (.X(n1508), 
	.A2(n1470), 
	.A1(n1471));
   SEN_INV_S_6 U1396 (.X(n1548), 
	.A(n1549));
   SEN_EN2_0P5 U1397 (.X(n372), 
	.A2(pprow1_qual[23]), 
	.A1(pprow1_qual[25]));
   SEN_EN2_S_2 U1398 (.X(net82550), 
	.A2(net82565), 
	.A1(net94383));
   SEN_EN2_0P5 U1399 (.X(net94383), 
	.A2(pprow1_qual[22]), 
	.A1(pprow1_qual[24]));
   SEN_INV_S_1 U1400 (.X(n1691), 
	.A(n1752));
   SEN_AO21B_6 U1401 (.X(n1522), 
	.B(n1519), 
	.A2(n1518), 
	.A1(n266));
   SEN_INV_S_1 U1402 (.X(n139), 
	.A(pprow7_qual[9]));
   SEN_ND2_G_1 U1403 (.X(n158), 
	.A2(n139), 
	.A1(n138));
   SEN_AN2_S_1 U1404 (.X(n1607), 
	.A2(pprow9_qual[6]), 
	.A1(pprow8_qual[8]));
   SEN_ND2_G_1 U1405 (.X(n146), 
	.A2(pprow6_qual[12]), 
	.A1(pprow7_qual[10]));
   SEN_NR2B_1 U1406 (.X(n148), 
	.B(n138), 
	.A(pprow7_qual[9]));
   SEN_ND2_G_1 U1407 (.X(n420), 
	.A2(pprow2_qual[20]), 
	.A1(net82508));
   SEN_ND2_G_1 U1408 (.X(n421), 
	.A2(pprow3_qual[18]), 
	.A1(net82508));
   SEN_ND2_G_1 U1409 (.X(n405), 
	.A2(n410), 
	.A1(n409));
   SEN_ND2_G_1 U1410 (.X(n410), 
	.A2(pprow2_qual[21]), 
	.A1(pprow3_qual[19]));
   SEN_ND2_G_1 U1411 (.X(n409), 
	.A2(net82508), 
	.A1(n124));
   SEN_INV_1 U1412 (.X(n419), 
	.A(n404));
   SEN_OAI21_S_2 U1413 (.X(n155), 
	.B(n154), 
	.A2(n152), 
	.A1(n150));
   SEN_NR2_1 U1414 (.X(n154), 
	.A2(n147), 
	.A1(net82486));
   SEN_ND2B_1 U1415 (.X(n152), 
	.B(n153), 
	.A(n127));
   SEN_ND2B_1 U1416 (.X(net88113), 
	.B(n363), 
	.A(net82348));
   SEN_INV_S_3 U1417 (.X(net84361), 
	.A(pprow0_qual[6]));
   SEN_EO2_S_0P5 U1418 (.X(n737), 
	.A2(n527), 
	.A1(pprow1_qual[8]));
   SEN_INV_S_1 U1419 (.X(net84160), 
	.A(pprow0_qual[10]));
   SEN_ND2_4 U1420 (.X(n1004), 
	.A2(n942), 
	.A1(n997));
   SEN_INV_S_1 U1421 (.X(n1195), 
	.A(n999));
   SEN_AO21B_4 U1422 (.X(n996), 
	.B(n1197), 
	.A2(pprow1_qual[0]), 
	.A1(pprow1_qual[1]));
   SEN_INV_S_1 U1423 (.X(net84200), 
	.A(net84001));
   SEN_EN2_1 U1425 (.X(net84057), 
	.A2(pprow3_qual[2]), 
	.A1(pprow2_qual[4]));
   SEN_INV_2 U1426 (.X(net83991), 
	.A(net83875));
   SEN_EN2_0P5 U1427 (.X(n1093), 
	.A2(pprow3_qual[7]), 
	.A1(pprow2_qual[9]));
   SEN_ND2_G_1 U1428 (.X(net83520), 
	.A2(pprow0_qual[16]), 
	.A1(C[16]));
   SEN_ND2_G_1 U1429 (.X(net83646), 
	.A2(pprow0_qual[15]), 
	.A1(C[15]));
   SEN_ND2_2 U1430 (.X(net83583), 
	.A2(pprow3_qual[8]), 
	.A1(pprow2_qual[10]));
   SEN_ND2_G_1 U1432 (.X(n1270), 
	.A2(pprow1_qual[12]), 
	.A1(pprow1_qual[14]));
   SEN_BUF_S_1 U1433 (.X(n434), 
	.A(n1354));
   SEN_EO2_S_0P5 U1434 (.X(n1244), 
	.A2(pprow5_qual[7]), 
	.A1(pprow4_qual[9]));
   SEN_EN2_0P5 U1435 (.X(n224), 
	.A2(pprow2_qual[13]), 
	.A1(pprow3_qual[11]));
   SEN_EO2_S_0P5 U1436 (.X(n459), 
	.A2(C[20]), 
	.A1(n1364));
   SEN_EO2_S_0P5 U1437 (.X(n375), 
	.A2(n525), 
	.A1(pprow1_qual[18]));
   SEN_EN2_0P5 U1438 (.X(net98319), 
	.A2(pprow1_qual[17]), 
	.A1(pprow1_qual[19]));
   SEN_INV_S_1 U1439 (.X(n1392), 
	.A(pprow0_qual[21]));
   SEN_EO2_S_0P5 U1442 (.X(n376), 
	.A2(pprow3_qual[14]), 
	.A1(pprow2_qual[16]));
   SEN_INV_S_1 U1443 (.X(net82977), 
	.A(net82878));
   SEN_ND2B_2 U1444 (.X(n1539), 
	.B(n815), 
	.A(n1488));
   SEN_ND2B_1 U1446 (.X(net95993), 
	.B(n400), 
	.A(n131));
   SEN_ND2_G_1 U1447 (.X(n400), 
	.A2(pprow3_qual[17]), 
	.A1(pprow2_qual[19]));
   SEN_EN2_0P5 U1448 (.X(n160), 
	.A2(pprow7_qual[9]), 
	.A1(pprow6_qual[11]));
   SEN_INV_6 U1449 (.X(net82773), 
	.A(net82771));
   SEN_ND2_2 U1450 (.X(n1713), 
	.A2(n1649), 
	.A1(n1650));
   SEN_INV_2 U1451 (.X(net82466), 
	.A(n370));
   SEN_INV_2 U1452 (.X(n254), 
	.A(n253));
   SEN_ND2_G_1 U1453 (.X(n253), 
	.A2(n1593), 
	.A1(n1594));
   SEN_INV_S_4 U1454 (.X(n1697), 
	.A(n1598));
   SEN_EN2_0P5 U1455 (.X(n413), 
	.A2(pprow3_qual[18]), 
	.A1(pprow2_qual[20]));
   SEN_ND2_T_1 U1457 (.X(n1611), 
	.A2(n1610), 
	.A1(n161));
   SEN_ND2_G_1 U1458 (.X(n411), 
	.A2(n420), 
	.A1(n421));
   SEN_INV_2 U1459 (.X(net82203), 
	.A(net82207));
   SEN_INV_3 U1460 (.X(net82202), 
	.A(net82206));
   SEN_EO2_2 U1461 (.X(n1808), 
	.A2(n717), 
	.A1(net82098));
   SEN_ND2B_1 U1462 (.X(n518), 
	.B(net85748), 
	.A(net91406));
   SEN_INV_1 U1463 (.X(net82165), 
	.A(net82167));
   SEN_NR2_T_1 U1464 (.X(net91363), 
	.A2(net91405), 
	.A1(net91397));
   SEN_ND2B_1 U1465 (.X(net91405), 
	.B(net85748), 
	.A(net91398));
   SEN_EN2_0P5 U1466 (.X(n183), 
	.A2(n182), 
	.A1(pprow9_qual[11]));
   SEN_INV_S_1 U1467 (.X(net91399), 
	.A(net91406));
   SEN_NR2_1 U1468 (.X(net91396), 
	.A2(net91398), 
	.A1(net91397));
   SEN_NR2_1 U1469 (.X(n359), 
	.A2(n361), 
	.A1(net91397));
   SEN_ND2_G_1 U1470 (.X(n361), 
	.A2(net90737), 
	.A1(net91410));
   SEN_INV_1 U1471 (.X(net82233), 
	.A(net82237));
   SEN_EO2_G_2 U1472 (.X(net85897), 
	.A2(n1816), 
	.A1(n758));
   SEN_AOI21_S_2 U1473 (.X(n366), 
	.B(net91413), 
	.A2(n367), 
	.A1(n369));
   SEN_INV_S_1 U1474 (.X(n367), 
	.A(n368));
   SEN_INV_S_1 U1475 (.X(net91413), 
	.A(net91419));
   SEN_OAI21B_4 U1476 (.X(net97350), 
	.B(n110), 
	.A2(n115), 
	.A1(net82455));
   SEN_ND2_G_1 U1477 (.X(n490), 
	.A2(net91406), 
	.A1(net91419));
   SEN_INV_S_1 U1478 (.X(net91407), 
	.A(net91415));
   SEN_NR2_1 U1479 (.X(net91415), 
	.A2(pprow1_qual[24]), 
	.A1(pprow1_qual[26]));
   SEN_ND2_G_1 U1480 (.X(net91406), 
	.A2(pprow1_qual[25]), 
	.A1(pprow1_qual[27]));
   SEN_INV_S_1 U1481 (.X(net91398), 
	.A(net91410));
   SEN_ND2_2 U1483 (.X(net84410), 
	.A2(pprow0_qual[2]), 
	.A1(net84732));
   SEN_EO2_S_0P5 U1484 (.X(n247), 
	.A2(n377), 
	.A1(n528));
   SEN_EO2_S_0P5 U1485 (.X(n915), 
	.A2(n913), 
	.A1(n933));
   SEN_ND2B_V1_2 U1486 (.X(net84116), 
	.B(net84160), 
	.A(C[10]));
   SEN_AN2_3 U1487 (.X(n704), 
	.A2(n969), 
	.A1(n1022));
   SEN_INV_2 U1488 (.X(n969), 
	.A(pprow1_qual[6]));
   SEN_INV_2 U1489 (.X(n1009), 
	.A(n994));
   SEN_ND2_T_1 U1490 (.X(n971), 
	.A2(n967), 
	.A1(n968));
   SEN_EN2_0P5 U1491 (.X(n538), 
	.A2(net97397), 
	.A1(net83936));
   SEN_EN2_0P5 U1492 (.X(n1025), 
	.A2(pprow1_qual[9]), 
	.A1(pprow1_qual[11]));
   SEN_ND2_6 U1493 (.X(n1103), 
	.A2(net84042), 
	.A1(n1018));
   SEN_ND2_2 U1494 (.X(n383), 
	.A2(net83875), 
	.A1(n1034));
   SEN_INV_S_1 U1496 (.X(net83516), 
	.A(pprow0_qual[17]));
   SEN_EO2_1 U1497 (.X(net86022), 
	.A2(pprow3_qual[9]), 
	.A1(pprow2_qual[11]));
   SEN_INV_S_1 U1498 (.X(net83614), 
	.A(net83612));
   SEN_EN2_0P5 U1499 (.X(n1238), 
	.A2(n1298), 
	.A1(n1297));
   SEN_MUXI2_S_2 U1500 (.X(net83223), 
	.S(n228), 
	.D1(n227), 
	.D0(n226));
   SEN_EO2_S_0P5 U1501 (.X(n227), 
	.A2(pprow3_qual[12]), 
	.A1(pprow2_qual[14]));
   SEN_ND2B_1 U1502 (.X(n226), 
	.B(net83111), 
	.A(n229));
   SEN_ND2B_1 U1503 (.X(net83127), 
	.B(net83220), 
	.A(net83223));
   SEN_EO2_DG_1 U1504 (.X(n1386), 
	.A2(n708), 
	.A1(n1388));
   SEN_EO2_S_0P5 U1505 (.X(n713), 
	.A2(pprow7_qual[7]), 
	.A1(pprow6_qual[9]));
   SEN_EO2_1 U1506 (.X(n667), 
	.A2(n522), 
	.A1(n1528));
   SEN_OAI21_5 U1507 (.X(n1657), 
	.B(n1645), 
	.A2(n1697), 
	.A1(n1698));
   SEN_INV_2 U1508 (.X(n1658), 
	.A(n1651));
   SEN_ND2_2 U1509 (.X(net82858), 
	.A2(net85257), 
	.A1(net82859));
   SEN_INV_1 U1510 (.X(n1665), 
	.A(n1713));
   SEN_INV_4 U1511 (.X(n1736), 
	.A(n1734));
   SEN_INV_2 U1512 (.X(n1737), 
	.A(n1735));
   SEN_ND2_2 U1513 (.X(net82394), 
	.A2(n1675), 
	.A1(net82499));
   SEN_AOAI211_2 U1514 (.X(n252), 
	.C(n1731), 
	.B(net82404), 
	.A2(n1732), 
	.A1(n1733));
   SEN_ND2_G_3 U1515 (.X(n584), 
	.A2(n248), 
	.A1(n1743));
   SEN_EO2_S_0P5 U1516 (.X(n1696), 
	.A2(n1749), 
	.A1(n1746));
   SEN_INV_S_3 U1517 (.X(net82194), 
	.A(net82195));
   SEN_EN2_S_4 U1518 (.X(net85931), 
	.A2(net82167), 
	.A1(n357));
   SEN_NR2_1 U1519 (.X(net90740), 
	.A2(n360), 
	.A1(n359));
   SEN_NR2_1 U1520 (.X(n360), 
	.A2(net91406), 
	.A1(net82179));
   SEN_INV_S_1 U1521 (.X(n1708), 
	.A(n1707));
   SEN_INV_2 U1522 (.X(n1769), 
	.A(n1768));
   SEN_EO2_S_0P5 U1523 (.X(n690), 
	.A2(n20), 
	.A1(n1780));
   SEN_INV_4 U1524 (.X(net84732), 
	.A(n290));
   SEN_EO2_S_0P5 U1525 (.X(n712), 
	.A2(n530), 
	.A1(pprow1_qual[2]));
   SEN_INV_2 U1526 (.X(n541), 
	.A(n540));
   SEN_INV_8 U1527 (.X(n1080), 
	.A(n1076));
   SEN_EO2_S_0P5 U1528 (.X(n1064), 
	.A2(C[14]), 
	.A1(net83829));
   SEN_OAOI211_3 U1529 (.X(n1062), 
	.C(n1059), 
	.B(n1060), 
	.A2(n1061), 
	.A1(n1112));
   SEN_ND2_G_1 U1530 (.X(n1041), 
	.A2(n1013), 
	.A1(n811));
   SEN_ND2B_4 U1531 (.X(n574), 
	.B(n457), 
	.A(net83453));
   SEN_EO2_S_0P5 U1532 (.X(n695), 
	.A2(net101248), 
	.A1(net83424));
   SEN_ND2_G_1 U1533 (.X(net83436), 
	.A2(n132), 
	.A1(net83189));
   SEN_EN2_0P5 U1534 (.X(n1295), 
	.A2(net83206), 
	.A1(net84636));
   SEN_INV_S_1 U1535 (.X(n454), 
	.A(net83206));
   SEN_EO2_G_2 U1536 (.X(n1462), 
	.A2(n560), 
	.A1(n689));
   SEN_EO2_S_0P5 U1537 (.X(n689), 
	.A2(n1474), 
	.A1(n1475));
   SEN_INV_2 U1538 (.X(net83095), 
	.A(net83098));
   SEN_ND2_3 U1540 (.X(net82190), 
	.A2(net82390), 
	.A1(net82389));
   SEN_BUF_2 U1541 (.X(n816), 
	.A(\bmul/neg13 ));
   SEN_BUF_S_4 U1542 (.X(n814), 
	.A(\bmul/neg9 ));
   SEN_EO2_S_0P5 U1543 (.X(n763), 
	.A2(net84654), 
	.A1(A[2]));
   SEN_ND2_G_1 U1544 (.X(n619), 
	.A2(net87845), 
	.A1(net87844));
   SEN_INV_S_1 U1545 (.X(net87844), 
	.A(pprow0_qual[0]));
   SEN_BUF_S_1 U1546 (.X(n808), 
	.A(\dp_cluster_0/N32 ));
   SEN_INV_2 U1547 (.X(net94322), 
	.A(net94321));
   SEN_INV_S_1 U1548 (.X(net94321), 
	.A(net84441));
   SEN_EO2_2 U1550 (.X(n952), 
	.A2(n931), 
	.A1(n932));
   SEN_INV_5 U1551 (.X(net84047), 
	.A(net84045));
   SEN_EN2_0P5 U1553 (.X(n1554), 
	.A2(net82641), 
	.A1(net82636));
   SEN_INV_S_1 U1554 (.X(n596), 
	.A(n1555));
   SEN_ND2_G_1 U1555 (.X(net82182), 
	.A2(net82056), 
	.A1(net82183));
   SEN_EO2_1 U1556 (.X(\bmul/one8 ), 
	.A2(n437), 
	.A1(A[16]));
   SEN_EO2_1 U1557 (.X(\bmul/one9 ), 
	.A2(n813), 
	.A1(A[18]));
   SEN_EO2_S_0P5 U1558 (.X(\bmul/one6 ), 
	.A2(n399), 
	.A1(A[12]));
   SEN_EO2_S_0P5 U1559 (.X(\bmul/one5 ), 
	.A2(\bmul/neg4 ), 
	.A1(A[10]));
   SEN_EO2_S_0P5 U1560 (.X(\dp_cluster_0/N290 ), 
	.A2(n280), 
	.A1(net89933));
   SEN_EN2_0P5 U1561 (.X(n280), 
	.A2(n283), 
	.A1(n282));
   SEN_EO2_S_0P5 U1562 (.X(Z[10]), 
	.A2(n984), 
	.A1(n655));
   SEN_OR2_1 U1563 (.X(n1119), 
	.A2(net83919), 
	.A1(n24));
   SEN_EO2_S_0P5 U1564 (.X(n672), 
	.A2(n569), 
	.A1(n1211));
   SEN_EO2_S_0P5 U1565 (.X(Z[19]), 
	.A2(n1325), 
	.A1(n676));
   SEN_EO2_S_0P5 U1566 (.X(Z[23]), 
	.A2(net82931), 
	.A1(net82930));
   SEN_EO2_S_0P5 U1567 (.X(Z[24]), 
	.A2(net82819), 
	.A1(n653));
   SEN_EO2_S_0P5 U1568 (.X(Z[26]), 
	.A2(n1666), 
	.A1(n654));
   SEN_EO2_S_0P5 U1569 (.X(n654), 
	.A2(net82523), 
	.A1(n19));
   SEN_EN2_0P5 U1570 (.X(Z[28]), 
	.A2(net82322), 
	.A1(n1716));
   SEN_EN2_1 U1571 (.X(net82320), 
	.A2(net86498), 
	.A1(net86381));
   SEN_ND2B_6 U1572 (.X(n1299), 
	.B(n1296), 
	.A(n1297));
   SEN_ND2_G_3 U1573 (.X(net87800), 
	.A2(net87797), 
	.A1(n186));
   SEN_AOI31_4 U1574 (.X(net82527), 
	.B(n1662), 
	.A3(n1664), 
	.A2(n1665), 
	.A1(n1663));
   SEN_ND2B_S_8 U1576 (.X(n443), 
	.B(n449), 
	.A(net84730));
   SEN_EO2_4 U1577 (.X(n1597), 
	.A2(net82659), 
	.A1(n759));
   SEN_INV_4 U1578 (.X(net82659), 
	.A(n350));
   SEN_AN2_S_8 U1579 (.X(net86517), 
	.A2(n1443), 
	.A1(n1444));
   SEN_AN2_6 U1580 (.X(n502), 
	.A2(n398), 
	.A1(net83329));
   SEN_INV_S_1 U1581 (.X(n1529), 
	.A(n1585));
   SEN_ND2_0P5 U1582 (.X(n1012), 
	.A2(net83550), 
	.A1(net83951));
   SEN_ND2_3 U1583 (.X(net84385), 
	.A2(n878), 
	.A1(n879));
   SEN_INV_2 U1584 (.X(n497), 
	.A(net82209));
   SEN_ND2_G_4 U1585 (.X(net82209), 
	.A2(n1736), 
	.A1(n1737));
   SEN_AOI211_G_2 U1586 (.X(net84230), 
	.B2(net84232), 
	.B1(net84119), 
	.A2(net84152), 
	.A1(net84231));
   SEN_AOAI211_6 U1588 (.X(net83521), 
	.C(net83646), 
	.B(net83731), 
	.A2(net83730), 
	.A1(net83729));
   SEN_EN2_DG_1 U1589 (.X(net82284), 
	.A2(n690), 
	.A1(n35));
   SEN_INV_S_1 U1590 (.X(n346), 
	.A(n353));
   SEN_AOI21_G_0P75 U1591 (.X(n489), 
	.B(n490), 
	.A2(net97350), 
	.A1(net91407));
   SEN_INV_4 U1592 (.X(net91426), 
	.A(net97350));
   SEN_EN2_DG_1 U1593 (.X(net82641), 
	.A2(n666), 
	.A1(n1553));
   SEN_BUF_1 U1594 (.X(net90993), 
	.A(net83413));
   SEN_ND2_T_2 U1595 (.X(n1440), 
	.A2(n1210), 
	.A1(n1211));
   SEN_EN2_S_3 U1597 (.X(n1210), 
	.A2(n1162), 
	.A1(net86306));
   SEN_ND2B_3 U1598 (.X(n1442), 
	.B(net82965), 
	.A(n1440));
   SEN_EO2_8 U1599 (.X(n583), 
	.A2(net82354), 
	.A1(n105));
   SEN_BUF_1 U1600 (.X(n104), 
	.A(n957));
   SEN_INV_32 U1601 (.X(n105), 
	.A(n1836));
   SEN_AN4B_2 U1602 (.X(n1204), 
	.B3(n1202), 
	.B2(n1247), 
	.B1(n434), 
	.A(n514));
   SEN_INV_S_2 U1603 (.X(n1050), 
	.A(n1048));
   SEN_ND2_G_1 U1604 (.X(n1225), 
	.A2(net83626), 
	.A1(n1264));
   SEN_INV_S_3 U1606 (.X(n288), 
	.A(C[1]));
   SEN_ND3_S_4 U1607 (.X(net83437), 
	.A3(n1279), 
	.A2(n1278), 
	.A1(n1254));
   SEN_ND2_3 U1608 (.X(n1278), 
	.A2(n1253), 
	.A1(n1280));
   SEN_ND3_T_4 U1609 (.X(net84359), 
	.A3(net84350), 
	.A2(net84385), 
	.A1(net84384));
   SEN_NR2_6 U1610 (.X(net83371), 
	.A2(net83380), 
	.A1(n591));
   SEN_OR3B_2 U1611 (.X(n945), 
	.B2(net84232), 
	.B1(net84237), 
	.A(net84147));
   SEN_AOI31_3 U1613 (.X(net84226), 
	.B(net84230), 
	.A3(net84228), 
	.A2(net84229), 
	.A1(net84227));
   SEN_EN2_0P5 U1616 (.X(net82938), 
	.A2(net86273), 
	.A1(net82939));
   SEN_EO2_2 U1617 (.X(net86273), 
	.A2(net82981), 
	.A1(net82982));
   SEN_ND2B_6 U1618 (.X(n1209), 
	.B(n1122), 
	.A(n1120));
   SEN_BUF_2 U1619 (.X(n107), 
	.A(n1496));
   SEN_EN2_0P5 U1621 (.X(n108), 
	.A2(pprow1_qual[24]), 
	.A1(pprow1_qual[26]));
   SEN_AN2_S_1 U1622 (.X(n109), 
	.A2(pprow3_qual[14]), 
	.A1(pprow2_qual[16]));
   SEN_AN2_S_1 U1623 (.X(n110), 
	.A2(pprow1_qual[23]), 
	.A1(pprow1_qual[25]));
   SEN_BUF_S_2 U1624 (.X(n558), 
	.A(n1004));
   SEN_AN2_S_1 U1625 (.X(n111), 
	.A2(n335), 
	.A1(net82454));
   SEN_INV_S_1 U1626 (.X(n561), 
	.A(C[25]));
   SEN_BUF_S_1 U1627 (.X(n815), 
	.A(\bmul/neg12 ));
   SEN_INV_3 U1628 (.X(n1153), 
	.A(pprow1_qual[11]));
   SEN_EN2_0P5 U1629 (.X(n112), 
	.A2(pprow1_qual[19]), 
	.A1(pprow1_qual[21]));
   SEN_EN2_0P5 U1630 (.X(n113), 
	.A2(pprow1_qual[20]), 
	.A1(pprow1_qual[22]));
   SEN_ND2_G_1 U1631 (.X(net83189), 
	.A2(pprow1_qual[15]), 
	.A1(pprow1_qual[17]));
   SEN_INV_2 U1632 (.X(n1632), 
	.A(n1628));
   SEN_INV_2 U1633 (.X(n1002), 
	.A(n902));
   SEN_ND2_G_3 U1634 (.X(n902), 
	.A2(n884), 
	.A1(n922));
   SEN_ND2_G_1 U1635 (.X(n1048), 
	.A2(pprow4_qual[0]), 
	.A1(pprow4_qual[1]));
   SEN_AN2_S_1 U1636 (.X(n115), 
	.A2(net82454), 
	.A1(net91386));
   SEN_EN2_0P5 U1637 (.X(n116), 
	.A2(n1791), 
	.A1(net82248));
   SEN_INV_2 U1638 (.X(n904), 
	.A(pprow1_qual[3]));
   SEN_INV_3 U1639 (.X(net83510), 
	.A(net83506));
   SEN_EN2_0P5 U1640 (.X(net82179), 
	.A2(pprow1_qual[26]), 
	.A1(pprow1_qual[28]));
   SEN_OR2_1 U1641 (.X(n117), 
	.A2(pprow4_qual[9]), 
	.A1(pprow5_qual[7]));
   SEN_BUF_S_1 U1642 (.X(n813), 
	.A(\bmul/neg8 ));
   SEN_OR2_1 U1643 (.X(n118), 
	.A2(pprow8_qual[12]), 
	.A1(pprow9_qual[10]));
   SEN_OR2_1 U1644 (.X(n119), 
	.A2(pprow10_qual[8]), 
	.A1(pprow11_qual[6]));
   SEN_AN2_S_1 U1645 (.X(n121), 
	.A2(n332), 
	.A1(n333));
   SEN_INV_2 U1646 (.X(n922), 
	.A(pprow1_qual[4]));
   SEN_EO2_S_0P5 U1647 (.X(n122), 
	.A2(pprow5_qual[6]), 
	.A1(pprow4_qual[8]));
   SEN_OR2_1 U1648 (.X(n123), 
	.A2(pprow12_qual[4]), 
	.A1(pprow13_qual[2]));
   SEN_AN2_S_1 U1649 (.X(n124), 
	.A2(pprow2_qual[20]), 
	.A1(pprow3_qual[18]));
   SEN_INV_4 U1650 (.X(n1201), 
	.A(n1196));
   SEN_EO2_S_0P5 U1651 (.X(n125), 
	.A2(pprow3_qual[15]), 
	.A1(pprow2_qual[17]));
   SEN_AN2_S_1 U1652 (.X(n126), 
	.A2(n215), 
	.A1(n216));
   SEN_INV_2 U1653 (.X(n476), 
	.A(net83455));
   SEN_EO2_DG_2 U1654 (.X(net83455), 
	.A2(n1218), 
	.A1(n1230));
   SEN_AN2_S_1 U1655 (.X(n127), 
	.A2(n156), 
	.A1(n157));
   SEN_OA21_2 U1656 (.X(n128), 
	.B(net95748), 
	.A2(net84006), 
	.A1(net84251));
   SEN_EN2_3 U1658 (.X(n161), 
	.A2(n159), 
	.A1(n162));
   SEN_OR2_1 U1659 (.X(n129), 
	.A2(pprow7_qual[10]), 
	.A1(pprow6_qual[12]));
   SEN_AN2_S_1 U1660 (.X(n130), 
	.A2(net91406), 
	.A1(net91398));
   SEN_INV_S_3 U1661 (.X(n1211), 
	.A(n1207));
   SEN_AN2_S_1 U1662 (.X(n131), 
	.A2(n407), 
	.A1(n406));
   SEN_OR2_1 U1663 (.X(n132), 
	.A2(pprow1_qual[15]), 
	.A1(pprow1_qual[17]));
   SEN_OR2_1 U1664 (.X(n133), 
	.A2(net91390), 
	.A1(net82171));
   SEN_OR2_1 U1665 (.X(n135), 
	.A2(n126), 
	.A1(n222));
   SEN_AN2_1 U1666 (.X(n136), 
	.A2(n188), 
	.A1(net83577));
   SEN_AN2_S_1 U1667 (.X(n137), 
	.A2(n1390), 
	.A1(net83114));
   SEN_EN2_0P5 U1668 (.X(n531), 
	.A2(C[10]), 
	.A1(net84160));
   SEN_ND2_T_1 U1669 (.X(n1383), 
	.A2(net83309), 
	.A1(n1304));
   SEN_INV_2 U1670 (.X(net83295), 
	.A(net83309));
   SEN_AOI211_G_2 U1671 (.X(n1655), 
	.B2(n1697), 
	.B1(n1653), 
	.A2(n1654), 
	.A1(n1698));
   SEN_NR2B_4 U1672 (.X(n151), 
	.B(n139), 
	.A(pprow6_qual[11]));
   SEN_OAI21_S_8 U1673 (.X(n159), 
	.B(n158), 
	.A2(n151), 
	.A1(net82721));
   SEN_INV_S_4 U1674 (.X(n144), 
	.A(n146));
   SEN_EN2_5 U1675 (.X(n162), 
	.A2(pprow6_qual[12]), 
	.A1(pprow7_qual[10]));
   SEN_AOI22_T_0P5 U1697 (.X(net82123), 
	.B2(pprow12_qual[4]), 
	.B1(pprow13_qual[2]), 
	.A2(n123), 
	.A1(net82130));
   SEN_OA2BB2_4 U1698 (.X(n179), 
	.B2(n181), 
	.B1(net85926), 
	.A2(n180), 
	.A1(net82137));
   SEN_INV_2 U1699 (.X(n181), 
	.A(net82141));
   SEN_ND2_T_2 U1700 (.X(n180), 
	.A2(net85926), 
	.A1(n181));
   SEN_EN2_0P5 U1701 (.X(n182), 
	.A2(pprow8_qual[13]), 
	.A1(pprow7_qual[15]));
   SEN_ND2_6 U1702 (.X(net83787), 
	.A2(net84005), 
	.A1(n650));
   SEN_OR2_DG_2 U1703 (.X(n184), 
	.A2(C[23]), 
	.A1(pprow0_qual[23]));
   SEN_INV_AS_10 U1704 (.X(n1137), 
	.A(n1175));
   SEN_INV_4 U1706 (.X(net87990), 
	.A(n206));
   SEN_ND2_G_1 U1707 (.X(n445), 
	.A2(pprow0_qual[7]), 
	.A1(net84730));
   SEN_INV_S_1 U1710 (.X(net84237), 
	.A(n442));
   SEN_INV_3 U1711 (.X(net82201), 
	.A(net82080));
   SEN_EN2_S_6 U1712 (.X(net82080), 
	.A2(n701), 
	.A1(n1808));
   SEN_INV_8 U1713 (.X(n292), 
	.A(n298));
   SEN_INV_S_1 U1714 (.X(net84425), 
	.A(net84378));
   SEN_INV_S_3 U1715 (.X(n206), 
	.A(n2054));
   SEN_EN2_S_3 U1717 (.X(net82934), 
	.A2(net82935), 
	.A1(net82936));
   SEN_ND2_2 U1718 (.X(net83513), 
	.A2(n567), 
	.A1(net83632));
   SEN_ND2_4 U1719 (.X(n195), 
	.A2(n194), 
	.A1(n196));
   SEN_INV_S_4 U1722 (.X(n191), 
	.A(net87797));
   SEN_OAI21_G_8 U1724 (.X(n186), 
	.B(n197), 
	.A2(n200), 
	.A1(n195));
   SEN_ND3B_2 U1725 (.X(net84005), 
	.B2(net84002), 
	.B1(net84007), 
	.A(net84006));
   SEN_ND2_S_3 U1726 (.X(n203), 
	.A2(net83891), 
	.A1(net83965));
   SEN_ND2_G_1 U1727 (.X(net83782), 
	.A2(net83891), 
	.A1(net83965));
   SEN_INV_S_6 U1728 (.X(net83962), 
	.A(n198));
   SEN_BUF_1 U1729 (.X(n202), 
	.A(net83961));
   SEN_INV_3 U1730 (.X(n201), 
	.A(\bmul/neg3 ));
   SEN_EO2_3 U1731 (.X(net84445), 
	.A2(net84448), 
	.A1(n862));
   SEN_NR2_T_2 U1732 (.X(net84448), 
	.A2(n204), 
	.A1(net84449));
   SEN_EO2_8 U1735 (.X(net86446), 
	.A2(net82773), 
	.A1(net82770));
   SEN_EN2_5 U1737 (.X(n1350), 
	.A2(n1322), 
	.A1(n205));
   SEN_ND2_G_1 U1739 (.X(n555), 
	.A2(n1201), 
	.A1(n1200));
   SEN_INV_3 U1740 (.X(n1126), 
	.A(n1123));
   SEN_NR2_T_1P5 U1742 (.X(net84281), 
	.A2(n444), 
	.A1(net84283));
   SEN_EN2_6 U1744 (.X(net82981), 
	.A2(n1396), 
	.A1(n208));
   SEN_EN2_DG_8 U1745 (.X(n208), 
	.A2(C[22]), 
	.A1(n1424));
   SEN_ND3_T_1P5 U1748 (.X(n1266), 
	.A3(n1439), 
	.A2(net82965), 
	.A1(n1263));
   SEN_EN2_S_3 U1749 (.X(n1709), 
	.A2(n1648), 
	.A1(n665));
   SEN_AOAI211_8 U1750 (.X(n1799), 
	.C(n1731), 
	.B(net82404), 
	.A2(n1732), 
	.A1(n1733));
   SEN_ND2B_V1DG_2 U1751 (.X(n322), 
	.B(net84445), 
	.A(net84441));
   SEN_NR2_1 U1752 (.X(n911), 
	.A2(n909), 
	.A1(n910));
   SEN_ND2_G_3 U1753 (.X(net84364), 
	.A2(n308), 
	.A1(n307));
   SEN_ND2_1P5 U1754 (.X(n573), 
	.A2(net88089), 
	.A1(net83453));
   SEN_ND2_3 U1755 (.X(n1806), 
	.A2(net82207), 
	.A1(net82206));
   SEN_EO3_1 U1756 (.X(n236), 
	.A3(n1127), 
	.A2(n1123), 
	.A1(n1102));
   SEN_EN2_3 U1757 (.X(n1423), 
	.A2(n692), 
	.A1(n1413));
   SEN_INV_1 U1758 (.X(net82516), 
	.A(net82514));
   SEN_AOI22_0P5 U1759 (.X(n209), 
	.B2(n1297), 
	.B1(n1298), 
	.A2(n1300), 
	.A1(n1299));
   SEN_EO2_6 U1761 (.X(net82323), 
	.A2(net86534), 
	.A1(net82385));
   SEN_NR2_1 U1762 (.X(n871), 
	.A2(n960), 
	.A1(n870));
   SEN_NR2_1 U1763 (.X(n870), 
	.A2(n876), 
	.A1(n869));
   SEN_ND2B_V1_2 U1764 (.X(n362), 
	.B(n363), 
	.A(net82348));
   SEN_INV_S_0P5 U1766 (.X(n1302), 
	.A(n1330));
   SEN_AO21B_1 U1767 (.X(n1296), 
	.B(n1330), 
	.A2(n1233), 
	.A1(n1234));
   SEN_ND2_0P5 U1770 (.X(n306), 
	.A2(net84364), 
	.A1(n305));
   SEN_ND2_T_4 U1771 (.X(net87549), 
	.A2(net84000), 
	.A1(net84006));
   SEN_AN2_3 U1772 (.X(n1375), 
	.A2(n1378), 
	.A1(n1377));
   SEN_AO21_1 U1773 (.X(net84441), 
	.B(n864), 
	.A2(n869), 
	.A1(n876));
   SEN_OA21_4 U1774 (.X(n303), 
	.B(net84191), 
	.A2(n308), 
	.A1(net84372));
   SEN_AN2_6 U1775 (.X(n1662), 
	.A2(n1711), 
	.A1(n384));
   SEN_ND2_0P8 U1776 (.X(n523), 
	.A2(n1201), 
	.A1(n1200));
   SEN_AO21B_4 U1778 (.X(n235), 
	.B(n1072), 
	.A2(net83862), 
	.A1(n1073));
   SEN_EO2_0P5 U1780 (.X(net84370), 
	.A2(n307), 
	.A1(net84189));
   SEN_INV_2 U1781 (.X(n1128), 
	.A(n1055));
   SEN_EO2_S_3 U1782 (.X(n1686), 
	.A2(n731), 
	.A1(n1694));
   SEN_AOAI211_6 U1783 (.X(n1694), 
	.C(n1634), 
	.B(n520), 
	.A2(n1635), 
	.A1(n1636));
   SEN_INV_4 U1784 (.X(net90746), 
	.A(net82162));
   SEN_INV_S_1 U1785 (.X(net91065), 
	.A(net83223));
   SEN_EO2_G_2 U1787 (.X(n1343), 
	.A2(n1302), 
	.A1(n1303));
   SEN_INV_2P5 U1788 (.X(n261), 
	.A(n1686));
   SEN_EN2_DG_1 U1790 (.X(net82069), 
	.A2(n697), 
	.A1(n34));
   SEN_EO2_0P5 U1792 (.X(n239), 
	.A2(n1064), 
	.A1(net83933));
   SEN_INV_S_6 U1793 (.X(n240), 
	.A(n781));
   SEN_INV_1P25 U1794 (.X(net82180), 
	.A(net82183));
   SEN_EN2_S_2 U1795 (.X(n1528), 
	.A2(n628), 
	.A1(n681));
   SEN_BUF_2 U1796 (.X(n241), 
	.A(net83610));
   SEN_AN3_4 U1797 (.X(n242), 
	.A3(n472), 
	.A2(net83331), 
	.A1(n327));
   SEN_INV_S_2 U1798 (.X(n1380), 
	.A(n1379));
   SEN_EO2_3 U1799 (.X(n243), 
	.A2(net86023), 
	.A1(net86022));
   SEN_EO2_1 U1800 (.X(n244), 
	.A2(net86023), 
	.A1(net86022));
   SEN_NR2_T_4 U1801 (.X(n1178), 
	.A2(n553), 
	.A1(n626));
   SEN_BUF_2 U1804 (.X(n248), 
	.A(n1768));
   SEN_ND2B_2 U1805 (.X(n1768), 
	.B(n1707), 
	.A(n1709));
   SEN_INV_2 U1806 (.X(net84411), 
	.A(net84413));
   SEN_INV_S_0P5 U1807 (.X(net82946), 
	.A(net82845));
   SEN_EN2_S_6 U1808 (.X(net82499), 
	.A2(n415), 
	.A1(n414));
   SEN_ND2B_V1_3 U1809 (.X(n1340), 
	.B(n1339), 
	.A(n1343));
   SEN_ND3_S_2 U1810 (.X(n1325), 
	.A3(n1267), 
	.A2(net83395), 
	.A1(n1441));
   SEN_BUF_S_4 U1811 (.X(net100928), 
	.A(net86213));
   SEN_INV_2 U1812 (.X(n1480), 
	.A(n1524));
   SEN_INV_2 U1813 (.X(n1527), 
	.A(n522));
   SEN_EO2_G_2 U1814 (.X(n1378), 
	.A2(n714), 
	.A1(n1370));
   SEN_ND2_G_3 U1815 (.X(n1509), 
	.A2(n1507), 
	.A1(n1508));
   SEN_ND3_8 U1816 (.X(n1584), 
	.A3(n1583), 
	.A2(n1582), 
	.A1(n1463));
   SEN_EO2_0P5 U1817 (.X(\dp_cluster_0/N289 ), 
	.A2(n2047), 
	.A1(net91110));
   SEN_AN2_S_3 U1818 (.X(n702), 
	.A2(n1247), 
	.A1(n556));
   SEN_ND2_2 U1819 (.X(n642), 
	.A2(net87762), 
	.A1(net86459));
   SEN_ND2_6 U1820 (.X(net83830), 
	.A2(n563), 
	.A1(net87761));
   SEN_INV_1 U1821 (.X(net82515), 
	.A(net82513));
   SEN_ND2B_6 U1822 (.X(n1330), 
	.B(pprow8_qual[1]), 
	.A(n1233));
   SEN_AOI22_4 U1823 (.X(net83025), 
	.B2(net83097), 
	.B1(net83096), 
	.A2(net83095), 
	.A1(net83094));
   SEN_INV_3 U1824 (.X(net83329), 
	.A(net83334));
   SEN_OR4B_4 U1825 (.X(n1432), 
	.B3(net82997), 
	.B2(n1430), 
	.B1(n1431), 
	.A(net82998));
   SEN_ND2_S_4 U1826 (.X(n1644), 
	.A2(net82555), 
	.A1(n1643));
   SEN_EN2_0P5 U1827 (.X(n933), 
	.A2(pprow2_qual[2]), 
	.A1(pprow3_qual[0]));
   SEN_AOAI211_6 U1828 (.X(n1785), 
	.C(n1755), 
	.B(n1756), 
	.A2(n1757), 
	.A1(n1758));
   SEN_ND2_4 U1829 (.X(net84006), 
	.A2(pprow3_qual[0]), 
	.A1(pprow2_qual[2]));
   SEN_EO2_DG_1 U1830 (.X(net83220), 
	.A2(n707), 
	.A1(n1344));
   SEN_OR2_1 U1831 (.X(n694), 
	.A2(n700), 
	.A1(n1680));
   SEN_BUF_1 U1832 (.X(n437), 
	.A(n812));
   SEN_AO21B_6 U1833 (.X(n581), 
	.B(n2038), 
	.A2(n1260), 
	.A1(net83418));
   SEN_EO3_6 U1835 (.X(n267), 
	.A3(pprow3_qual[16]), 
	.A2(pprow2_qual[18]), 
	.A1(n1514));
   SEN_ND2_T_8 U1836 (.X(n1698), 
	.A2(n254), 
	.A1(n1592));
   SEN_BUF_1 U1838 (.X(n255), 
	.A(pprow5_qual[3]));
   SEN_INV_1P25 U1839 (.X(net84351), 
	.A(net84357));
   SEN_ND2_G_1 U1840 (.X(n263), 
	.A2(net83552), 
	.A1(n488));
   SEN_INV_6 U1841 (.X(n408), 
	.A(net82703));
   SEN_ND2_T_2 U1842 (.X(n1767), 
	.A2(n1708), 
	.A1(n1709));
   SEN_ND2_3 U1843 (.X(net83098), 
	.A2(n1350), 
	.A1(n1349));
   SEN_OR2_DG_8 U1845 (.X(n257), 
	.A2(pprow6_qual[4]), 
	.A1(pprow7_qual[2]));
   SEN_INV_4 U1847 (.X(n1680), 
	.A(n1613));
   SEN_INV_2P5 U1848 (.X(n1298), 
	.A(n1296));
   SEN_EN2_1 U1849 (.X(n693), 
	.A2(net85815), 
	.A1(n462));
   SEN_INV_8 U1850 (.X(n1097), 
	.A(n1094));
   SEN_INV_S_0P5 U1851 (.X(n660), 
	.A(n1103));
   SEN_OA2BB2_4 U1852 (.X(net82975), 
	.B2(net82977), 
	.B1(net102542), 
	.A2(net82976), 
	.A1(net82734));
   SEN_BUF_1 U1853 (.X(n258), 
	.A(n541));
   SEN_INV_4 U1854 (.X(n916), 
	.A(n920));
   SEN_OR3B_4 U1855 (.X(n1306), 
	.B2(n1180), 
	.B1(n810), 
	.A(n1179));
   SEN_ND2_T_3 U1856 (.X(net83965), 
	.A2(n504), 
	.A1(n503));
   SEN_ND2_T_6 U1857 (.X(net83891), 
	.A2(n1088), 
	.A1(n1089));
   SEN_NR2_S_1 U1858 (.X(net83958), 
	.A2(net83580), 
	.A1(net83782));
   SEN_INV_S_0P5 U1859 (.X(n259), 
	.A(net84241));
   SEN_INV_S_0P5 U1860 (.X(n260), 
	.A(n1079));
   SEN_NR2_G_0P65 U1861 (.X(n910), 
	.A2(n905), 
	.A1(n963));
   SEN_ND2_T_0P5 U1862 (.X(n909), 
	.A2(n908), 
	.A1(n616));
   SEN_ND2_S_4 U1863 (.X(net97222), 
	.A2(net84196), 
	.A1(net89993));
   SEN_AO21B_2 U1864 (.X(net95846), 
	.B(net83849), 
	.A2(net83372), 
	.A1(net83371));
   SEN_NR2B_V1DG_3 U1865 (.X(n979), 
	.B(n975), 
	.A(net86124));
   SEN_INV_3 U1866 (.X(net87763), 
	.A(net86459));
   SEN_OA22_1 U1867 (.X(n488), 
	.B2(n485), 
	.B1(net86274), 
	.A2(n484), 
	.A1(n2043));
   SEN_OAI21_G_8 U1868 (.X(n1674), 
	.B(n1624), 
	.A2(n1626), 
	.A1(n1625));
   SEN_INV_4 U1869 (.X(net95561), 
	.A(net82879));
   SEN_ND2_2 U1870 (.X(net94058), 
	.A2(n265), 
	.A1(n379));
   SEN_ND2_T_1 U1871 (.X(n977), 
	.A2(net84148), 
	.A1(net84147));
   SEN_INV_1P5 U1872 (.X(n1415), 
	.A(n1414));
   SEN_EN3_6 U1873 (.X(n1188), 
	.A3(net83678), 
	.A2(net90884), 
	.A1(n1142));
   SEN_OR2_2P5 U1874 (.X(n1049), 
	.A2(pprow5_qual[0]), 
	.A1(pprow4_qual[2]));
   SEN_AOI21B_3 U1875 (.X(n1032), 
	.B(n1083), 
	.A2(n1049), 
	.A1(n1031));
   SEN_EO2_2 U1877 (.X(net82237), 
	.A2(n1796), 
	.A1(n728));
   SEN_INV_2 U1878 (.X(n961), 
	.A(n1199));
   SEN_OR4B_4 U1879 (.X(n1354), 
	.B3(n1195), 
	.B2(n1199), 
	.B1(n1196), 
	.A(n1194));
   SEN_OAOI211_4 U1880 (.X(n973), 
	.C(n1009), 
	.B(n970), 
	.A2(n971), 
	.A1(n972));
   SEN_INV_4 U1881 (.X(net94359), 
	.A(net85046));
   SEN_INV_1P25 U1882 (.X(n1535), 
	.A(pprow10_qual[2]));
   SEN_AOAI211_G_1 U1883 (.X(n1782), 
	.C(n1751), 
	.B(n1752), 
	.A2(n1753), 
	.A1(n1754));
   SEN_INV_1 U1884 (.X(n1485), 
	.A(n1519));
   SEN_INV_1P25 U1885 (.X(n309), 
	.A(n307));
   SEN_NR2_T_6 U1886 (.X(net85173), 
	.A2(net84358), 
	.A1(net86078));
   SEN_AO21B_4 U1887 (.X(net86655), 
	.B(n1258), 
	.A2(n1365), 
	.A1(net86332));
   SEN_AOI21_T_3 U1888 (.X(n422), 
	.B(n405), 
	.A2(n404), 
	.A1(n403));
   SEN_INV_S_0P5 U1889 (.X(n268), 
	.A(net83298));
   SEN_INV_S_4 U1890 (.X(n269), 
	.A(pprow0_qual[2]));
   SEN_ND2B_4 U1891 (.X(n275), 
	.B(n283), 
	.A(n282));
   SEN_ND2_S_0P5 U1892 (.X(n281), 
	.A2(pprow0_qual[2]), 
	.A1(net84732));
   SEN_ND2_T_3 U1893 (.X(net84392), 
	.A2(n269), 
	.A1(n290));
   SEN_INV_4 U1894 (.X(n291), 
	.A(n287));
   SEN_ND2_G_1 U1895 (.X(n285), 
	.A2(pprow0_qual[1]), 
	.A1(net84734));
   SEN_INV_1 U1896 (.X(net84654), 
	.A(n287));
   SEN_EO2_G_4 U1897 (.X(net83499), 
	.A2(n294), 
	.A1(net83627));
   SEN_INV_4 U1898 (.X(net83498), 
	.A(net83499));
   SEN_OAI21_S_8 U1899 (.X(net83370), 
	.B(net83513), 
	.A2(net83512), 
	.A1(n293));
   SEN_AOA211_DG_8 U1901 (.X(n299), 
	.C(n292), 
	.B(net84275), 
	.A2(n297), 
	.A1(net84183));
   SEN_INV_2P5 U1902 (.X(net82427), 
	.A(net82313));
   SEN_ND2_S_2 U1903 (.X(net82634), 
	.A2(net82317), 
	.A1(net82315));
   SEN_INV_1 U1904 (.X(net82833), 
	.A(net82829));
   SEN_INV_S_6 U1905 (.X(n302), 
	.A(net82839));
   SEN_EO2_0P5 U1906 (.X(net82930), 
	.A2(net82827), 
	.A1(net82829));
   SEN_INV_4 U1907 (.X(net90258), 
	.A(net84183));
   SEN_INV_S_0P5 U1908 (.X(net89992), 
	.A(net84273));
   SEN_AOI31_1 U1910 (.X(net84371), 
	.B(n305), 
	.A3(net84365), 
	.A2(net84366), 
	.A1(net83383));
   SEN_INV_2 U1911 (.X(n308), 
	.A(net84189));
   SEN_AOI211_0P5 U1912 (.X(net83495), 
	.B2(n315), 
	.B1(net83496), 
	.A2(net82965), 
	.A1(net83397));
   SEN_ND4B_1 U1913 (.X(net83626), 
	.B3(net90993), 
	.B2(net83412), 
	.B1(net83408), 
	.A(net96981));
   SEN_NR2_G_2 U1914 (.X(net96981), 
	.A2(net83919), 
	.A1(net83918));
   SEN_ND2B_V1_2 U1915 (.X(net83412), 
	.B(net83813), 
	.A(net83820));
   SEN_MUX2_4 U1916 (.X(net83497), 
	.S(net94064), 
	.D1(net94058), 
	.D0(net94057));
   SEN_AO21B_4 U1917 (.X(net86382), 
	.B(net82195), 
	.A2(net82190), 
	.A1(net82385));
   SEN_EO2_2 U1918 (.X(net82383), 
	.A2(net82188), 
	.A1(net82189));
   SEN_AOI21B_3 U1919 (.X(net82321), 
	.B(net82308), 
	.A2(net82302), 
	.A1(net82322));
   SEN_ND2B_6 U1920 (.X(net83383), 
	.B(net84378), 
	.A(n321));
   SEN_EN3_0P5 U1921 (.X(\dp_cluster_0/N291 ), 
	.A3(net84443), 
	.A2(net84442), 
	.A1(net94322));
   SEN_INV_4 U1922 (.X(net83384), 
	.A(net83168));
   SEN_AN3_8 U1923 (.X(net94176), 
	.A3(net86517), 
	.A2(n41), 
	.A1(net82850));
   SEN_ND2_T_0P5 U1924 (.X(net83395), 
	.A2(net82850), 
	.A1(n41));
   SEN_ND3_S_0P5 U1925 (.X(net82941), 
	.A3(net82850), 
	.A2(n41), 
	.A1(net86517));
   SEN_NR2_S_0P5 U1926 (.X(net82931), 
	.A2(n326), 
	.A1(net82932));
   SEN_AN2_3 U1927 (.X(net86483), 
	.A2(net82842), 
	.A1(n324));
   SEN_INV_S_3 U1928 (.X(n324), 
	.A(net82843));
   SEN_AOI21B_3 U1929 (.X(n1162), 
	.B(net83512), 
	.A2(n436), 
	.A1(net83507));
   SEN_EO2_2 U1930 (.X(Z[27]), 
	.A2(n1667), 
	.A1(n1668));
   SEN_AOI21B_2 U1931 (.X(n1667), 
	.B(net82432), 
	.A2(net82430), 
	.A1(n1666));
   SEN_INV_8 U1932 (.X(net82503), 
	.A(net82499));
   SEN_AO21B_2 U1933 (.X(n1399), 
	.B(n1455), 
	.A2(n1326), 
	.A1(n1443));
   SEN_ND3_T_2 U1934 (.X(net83789), 
	.A3(net83685), 
	.A2(n482), 
	.A1(net83550));
   SEN_EO3_6 U1935 (.X(n1524), 
	.A3(n1513), 
	.A2(n1512), 
	.A1(n1514));
   SEN_EN2_DG_8 U1936 (.X(n1323), 
	.A2(n1350), 
	.A1(n1349));
   SEN_ND2_6 U1937 (.X(n1384), 
	.A2(n601), 
	.A1(n1382));
   SEN_EO2_4 U1938 (.X(net82188), 
	.A2(n496), 
	.A1(n495));
   SEN_AOI31_3 U1939 (.X(n496), 
	.B(n497), 
	.A3(net82394), 
	.A2(net82210), 
	.A1(net82395));
   SEN_NR2_T_4 U1940 (.X(n348), 
	.A2(n337), 
	.A1(n340));
   SEN_AN2_6 U1941 (.X(n349), 
	.A2(n333), 
	.A1(net82562));
   SEN_ND3_T_4 U1942 (.X(n351), 
	.A3(n348), 
	.A2(n352), 
	.A1(n354));
   SEN_INV_S_0P5 U1943 (.X(net90737), 
	.A(net82179));
   SEN_EN2_0P5 U1944 (.X(n357), 
	.A2(C[30]), 
	.A1(n356));
   SEN_INV_S_1 U1945 (.X(n356), 
	.A(pprow0_qual[30]));
   SEN_AOAI211_3 U1946 (.X(net82162), 
	.C(net82166), 
	.B(net82165), 
	.A2(n356), 
	.A1(net82163));
   SEN_OAI21B_2 U1947 (.X(n369), 
	.B(n110), 
	.A2(n115), 
	.A1(net82455));
   SEN_NR2_T_4 U1948 (.X(n365), 
	.A2(n110), 
	.A1(n108));
   SEN_OAI21_5 U1949 (.X(net87786), 
	.B(n365), 
	.A2(n115), 
	.A1(net82455));
   SEN_INV_0P8 U1950 (.X(net82454), 
	.A(pprow1_qual[23]));
   SEN_INV_S_2 U1951 (.X(net82078), 
	.A(net82082));
   SEN_ND2_2 U1952 (.X(net82076), 
	.A2(net82077), 
	.A1(net82078));
   SEN_ND2_S_0P5 U1953 (.X(net82564), 
	.A2(pprow1_qual[22]), 
	.A1(pprow1_qual[24]));
   SEN_INV_S_0P5 U1954 (.X(net82562), 
	.A(pprow1_qual[22]));
   SEN_INV_S_0P5 U1955 (.X(n1654), 
	.A(n1652));
   SEN_EN2_DG_4 U1956 (.X(n433), 
	.A2(n1547), 
	.A1(n1597));
   SEN_BUF_1 U1957 (.X(net97397), 
	.A(C[13]));
   SEN_AO21B_2 U1958 (.X(n730), 
	.B(n925), 
	.A2(n902), 
	.A1(n885));
   SEN_EN2_1 U1959 (.X(n498), 
	.A2(net82236), 
	.A1(net82237));
   SEN_OA2BB2_8 U1960 (.X(n1810), 
	.B2(n1808), 
	.B1(n701), 
	.A2(n1809), 
	.A1(n1817));
   SEN_BUF_1 U1961 (.X(n386), 
	.A(n1376));
   SEN_INV_2 U1962 (.X(n1349), 
	.A(n1352));
   SEN_BUF_1 U1963 (.X(n373), 
	.A(n1440));
   SEN_ND2_T_4 U1964 (.X(n1185), 
	.A2(n1184), 
	.A1(n1187));
   SEN_BUF_1 U1965 (.X(n377), 
	.A(pprow1_qual[1]));
   SEN_INV_S_2 U1966 (.X(n1781), 
	.A(n1777));
   SEN_INV_S_1P5 U1968 (.X(n380), 
	.A(n484));
   SEN_EO2_2 U1969 (.X(n987), 
	.A2(n686), 
	.A1(net84121));
   SEN_NR2B_V1_8 U1970 (.X(net86078), 
	.B(net84391), 
	.A(n566));
   SEN_NR2_6 U1971 (.X(n1200), 
	.A2(n623), 
	.A1(n1199));
   SEN_EN2_3 U1972 (.X(n671), 
	.A2(n1742), 
	.A1(n1741));
   SEN_EO2_S_3 U1973 (.X(net83844), 
	.A2(n1062), 
	.A1(n1063));
   SEN_EN2_DG_1 U1974 (.X(n1660), 
	.A2(n683), 
	.A1(n1630));
   SEN_ND2_T_1 U1975 (.X(n1056), 
	.A2(net83798), 
	.A1(n383));
   SEN_EO2_DG_8 U1976 (.X(n385), 
	.A2(n636), 
	.A1(net83295));
   SEN_BUF_1 U1977 (.X(n387), 
	.A(C[8]));
   SEN_EN2_5 U1978 (.X(net82429), 
	.A2(net82527), 
	.A1(n388));
   SEN_EO2_DG_8 U1979 (.X(n388), 
	.A2(n1709), 
	.A1(n1707));
   SEN_AN2_S_1P5 U1980 (.X(n700), 
	.A2(n1614), 
	.A1(net82616));
   SEN_NR2_G_1 U1981 (.X(n429), 
	.A2(net83574), 
	.A1(net83573));
   SEN_EO2_G_1 U1982 (.X(n692), 
	.A2(n1414), 
	.A1(n1416));
   SEN_NR2_T_0P5 U1983 (.X(n1000), 
	.A2(pprow1_qual[8]), 
	.A1(pprow1_qual[6]));
   SEN_INV_2 U1984 (.X(n391), 
	.A(n1605));
   SEN_AN2_S_1 U1985 (.X(n392), 
	.A2(pprow0_qual[7]), 
	.A1(pprow0_qual[8]));
   SEN_OAOI211_4 U1986 (.X(net83743), 
	.C(n1273), 
	.B(n669), 
	.A2(n1154), 
	.A1(n1155));
   SEN_EO2_2 U1987 (.X(n1042), 
	.A2(n1034), 
	.A1(net83875));
   SEN_OAI21_S_4 U1989 (.X(net84413), 
	.B(n878), 
	.A2(n879), 
	.A1(net84415));
   SEN_ND2B_V1_8 U1990 (.X(net82721), 
	.B(n1506), 
	.A(n768));
   SEN_INV_1 U1991 (.X(n1193), 
	.A(n1008));
   SEN_ND2_S_0P5 U1992 (.X(n394), 
	.A2(net83844), 
	.A1(net83843));
   SEN_EO2_1 U1993 (.X(net94057), 
	.A2(net83612), 
	.A1(net83611));
   SEN_ND3_T_3 U1994 (.X(n877), 
	.A3(n996), 
	.A2(n779), 
	.A1(n923));
   SEN_ND2_2 U1995 (.X(n1688), 
	.A2(n1686), 
	.A1(n1687));
   SEN_OAI21_G_16 U1996 (.X(n404), 
	.B(n417), 
	.A2(n416), 
	.A1(n408));
   SEN_ND2_8 U1997 (.X(net82348), 
	.A2(net87786), 
	.A1(net87787));
   SEN_ND3_S_2 U1998 (.X(n1113), 
	.A3(n1148), 
	.A2(n620), 
	.A1(n1147));
   SEN_EO2_8 U1999 (.X(net83153), 
	.A2(n456), 
	.A1(n455));
   SEN_BUF_6 U2000 (.X(n810), 
	.A(\bmul/neg5 ));
   SEN_INV_1 U2001 (.X(net88056), 
	.A(net84734));
   SEN_OAOI211_4 U2002 (.X(n1648), 
	.C(n698), 
	.B(n1700), 
	.A2(n1697), 
	.A1(n1698));
   SEN_ND2_4 U2003 (.X(n1233), 
	.A2(pprow8_qual[0]), 
	.A1(n814));
   SEN_OAOI211_8 U2004 (.X(n1796), 
	.C(n1717), 
	.B(n1718), 
	.A2(pprow8_qual[10]), 
	.A1(pprow9_qual[8]));
   SEN_AOI21B_4 U2005 (.X(net83530), 
	.B(n1252), 
	.A2(n1281), 
	.A1(n1224));
   SEN_EO3_DG_1 U2006 (.X(n1352), 
	.A3(n1343), 
	.A2(n1342), 
	.A1(n209));
   SEN_EN2_DG_8 U2007 (.X(n396), 
	.A2(C[16]), 
	.A1(net83640));
   SEN_AOAI211_6 U2008 (.X(n1186), 
	.C(n1124), 
	.B(n1125), 
	.A2(n1126), 
	.A1(n1127));
   SEN_ND3_T_4 U2009 (.X(net84115), 
	.A3(n443), 
	.A2(net84153), 
	.A1(net84152));
   SEN_ND2_4 U2010 (.X(net83798), 
	.A2(n485), 
	.A1(n484));
   SEN_OAOI211_G_8 U2011 (.X(n1682), 
	.C(n1607), 
	.B(n1608), 
	.A2(pprow8_qual[8]), 
	.A1(pprow9_qual[6]));
   SEN_ND2_T_4 U2012 (.X(net87787), 
	.A2(n108), 
	.A1(net91408));
   SEN_EO2_4 U2013 (.X(n665), 
	.A2(net82467), 
	.A1(net82466));
   SEN_EN2_8 U2014 (.X(n1094), 
	.A2(n1054), 
	.A1(n618));
   SEN_EN2_1 U2015 (.X(n1040), 
	.A2(n380), 
	.A1(net83954));
   SEN_INV_4 U2016 (.X(net82521), 
	.A(net82522));
   SEN_NR2_0P8 U2017 (.X(n510), 
	.A2(net84057), 
	.A1(net84063));
   SEN_NR2_T_4 U2018 (.X(n412), 
	.A2(pprow3_qual[18]), 
	.A1(pprow2_qual[20]));
   SEN_ND2_4 U2019 (.X(n416), 
	.A2(net82701), 
	.A1(net82702));
   SEN_AOI22_T_4 U2020 (.X(n417), 
	.B2(pprow3_qual[17]), 
	.B1(pprow2_qual[19]), 
	.A2(n418), 
	.A1(net82702));
   SEN_OAI21B_4 U2021 (.X(n415), 
	.B(n124), 
	.A2(n412), 
	.A1(n419));
   SEN_ND2_4 U2022 (.X(n403), 
	.A2(n421), 
	.A1(n420));
   SEN_EN2_5 U2023 (.X(n414), 
	.A2(net82510), 
	.A1(net82511));
   SEN_ND2_2 U2024 (.X(n428), 
	.A2(net83566), 
	.A1(net83565));
   SEN_AN2_S_1P5 U2025 (.X(n425), 
	.A2(net83583), 
	.A1(net83582));
   SEN_AN3B_2 U2026 (.X(n431), 
	.B2(net83891), 
	.B1(net83581), 
	.A(net83580));
   SEN_INV_S_6 U2027 (.X(n432), 
	.A(net83787));
   SEN_OR2_2 U2028 (.X(net83565), 
	.A2(pprow3_qual[8]), 
	.A1(pprow2_qual[10]));
   SEN_NR2_T_3 U2029 (.X(net85252), 
	.A2(n130), 
	.A1(n489));
   SEN_ND2B_V1_1 U2030 (.X(n891), 
	.B(pprow2_qual[1]), 
	.A(n934));
   SEN_ND2_6 U2031 (.X(n1624), 
	.A2(n1623), 
	.A1(net82595));
   SEN_INV_4 U2032 (.X(net82555), 
	.A(net82550));
   SEN_ND2_2 U2033 (.X(net87542), 
	.A2(net103418), 
	.A1(net87541));
   SEN_NR2_6 U2034 (.X(net82161), 
	.A2(n516), 
	.A1(net91363));
   SEN_INV_4 U2035 (.X(n1109), 
	.A(pprow1_qual[10]));
   SEN_ND2_T_2 U2036 (.X(n1190), 
	.A2(pprow1_qual[10]), 
	.A1(pprow1_qual[12]));
   SEN_AOAI211_8 U2037 (.X(n1590), 
	.C(n1533), 
	.B(net82768), 
	.A2(n1534), 
	.A1(n1535));
   SEN_OAI21_S_4 U2038 (.X(net82850), 
	.B(net95817), 
	.A2(n1266), 
	.A1(n1265));
   SEN_AOI21_S_4 U2039 (.X(n1160), 
	.B(n1159), 
	.A2(net83735), 
	.A1(n778));
   SEN_ND2B_6 U2040 (.X(n1592), 
	.B(net82875), 
	.A(net87627));
   SEN_AN3_4 U2041 (.X(n651), 
	.A3(net95774), 
	.A2(net84056), 
	.A1(net84063));
   SEN_ND2B_V1_4 U2042 (.X(net87799), 
	.B(net87798), 
	.A(net87797));
   SEN_INV_2 U2043 (.X(n1133), 
	.A(n1132));
   SEN_INV_2 U2044 (.X(net83781), 
	.A(n203));
   SEN_INV_S_3 U2045 (.X(n1712), 
	.A(n1711));
   SEN_ND2_G_4 U2046 (.X(net84001), 
	.A2(pprow3_qual[2]), 
	.A1(pprow2_qual[4]));
   SEN_EO2_G_8 U2047 (.X(n1581), 
	.A2(n1419), 
	.A1(n1420));
   SEN_INV_3 U2048 (.X(n884), 
	.A(pprow1_qual[2]));
   SEN_ND2_G_4 U2049 (.X(n1197), 
	.A2(pprow1_qual[0]), 
	.A1(pprow1_qual[2]));
   SEN_BUF_1 U2051 (.X(n560), 
	.A(n1473));
   SEN_INV_0P5 U2052 (.X(n438), 
	.A(n511));
   SEN_INV_S_8 U2053 (.X(n1052), 
	.A(n1051));
   SEN_ND2_4 U2054 (.X(n1008), 
	.A2(n997), 
	.A1(n1058));
   SEN_OAI21_G_1 U2055 (.X(n1017), 
	.B(net83820), 
	.A2(n989), 
	.A1(net86390));
   SEN_INV_S_2 U2056 (.X(n989), 
	.A(n986));
   SEN_ND2_T_1 U2057 (.X(n934), 
	.A2(pprow2_qual[0]), 
	.A1(net84650));
   SEN_ND2_2 U2059 (.X(net84058), 
	.A2(net84056), 
	.A1(net84063));
   SEN_ND2_0P8 U2060 (.X(n1213), 
	.A2(pprow7_qual[0]), 
	.A1(pprow6_qual[2]));
   SEN_NR2_G_4 U2061 (.X(n1510), 
	.A2(n1508), 
	.A1(n1507));
   SEN_EO2_1 U2062 (.X(n681), 
	.A2(n1508), 
	.A1(n1507));
   SEN_AN3_S_4 U2064 (.X(n617), 
	.A3(net83958), 
	.A2(n36), 
	.A1(net83559));
   SEN_INV_S_2 U2066 (.X(net83209), 
	.A(net83214));
   SEN_EN3_6 U2067 (.X(net84045), 
	.A3(n1019), 
	.A2(n534), 
	.A1(net84081));
   SEN_AN5_4 U2068 (.X(n456), 
	.A5(net84636), 
	.A4(net83205), 
	.A3(net83203), 
	.A2(net83166), 
	.A1(n22));
   SEN_ND2_2 U2070 (.X(net83571), 
	.A2(pprow3_qual[5]), 
	.A1(pprow2_qual[7]));
   SEN_ND2_T_1 U2071 (.X(n1533), 
	.A2(pprow11_qual[0]), 
	.A1(pprow10_qual[2]));
   SEN_ND2_G_1 U2072 (.X(n589), 
	.A2(n588), 
	.A1(n742));
   SEN_INV_2 U2073 (.X(n463), 
	.A(n588));
   SEN_INV_S_0P5 U2074 (.X(net95774), 
	.A(net83999));
   SEN_INV_0P65 U2075 (.X(n1331), 
	.A(pprow9_qual[0]));
   SEN_INV_S_6 U2077 (.X(n623), 
	.A(n622));
   SEN_AOI21_S_4 U2078 (.X(net83156), 
	.B(n439), 
	.A2(net82983), 
	.A1(net94217));
   SEN_ND2B_4 U2079 (.X(net83608), 
	.B(n379), 
	.A(net83609));
   SEN_EO3_DG_4 U2080 (.X(n1207), 
	.A3(n251), 
	.A2(n1187), 
	.A1(n1186));
   SEN_EO2_0P5 U2081 (.X(n721), 
	.A2(pprow1_qual[8]), 
	.A1(pprow1_qual[10]));
   SEN_ND2_T_3 U2082 (.X(n903), 
	.A2(n876), 
	.A1(n904));
   SEN_NR2_G_4 U2083 (.X(n622), 
	.A2(n1197), 
	.A1(n1198));
   SEN_INV_S_0P5 U2084 (.X(n550), 
	.A(n898));
   SEN_INV_S_6 U2085 (.X(net84395), 
	.A(net84357));
   SEN_INV_S_2 U2086 (.X(net82389), 
	.A(net82386));
   SEN_AOI21B_1 U2087 (.X(n1167), 
	.B(n1213), 
	.A2(n766), 
	.A1(n812));
   SEN_BUF_1P5 U2088 (.X(n774), 
	.A(n1280));
   SEN_ND2_4 U2089 (.X(n1645), 
	.A2(n1598), 
	.A1(n1652));
   SEN_ND2B_V1DG_8 U2090 (.X(net83951), 
	.B(n1033), 
	.A(net83993));
   SEN_AO2BB2_DG_4 U2091 (.X(n1174), 
	.B2(pprow4_qual[5]), 
	.B1(pprow5_qual[3]), 
	.A2(n1136), 
	.A1(n1137));
   SEN_AO2BB2_DG_4 U2092 (.X(n553), 
	.B2(pprow4_qual[5]), 
	.B1(pprow5_qual[3]), 
	.A2(n1136), 
	.A1(n1137));
   SEN_INV_S_0P5 U2093 (.X(n967), 
	.A(n1010));
   SEN_ND3_T_0P5 U2094 (.X(n1285), 
	.A3(n1354), 
	.A2(n523), 
	.A1(n556));
   SEN_INV_S_6 U2095 (.X(net84202), 
	.A(pprow3_qual[2]));
   SEN_ND2_T_2 U2096 (.X(n1622), 
	.A2(n1620), 
	.A1(n1621));
   SEN_NR2_S_2 U2097 (.X(net82702), 
	.A2(n1566), 
	.A1(n131));
   SEN_INV_2 U2098 (.X(n1566), 
	.A(n1565));
   SEN_OAOI211_2 U2100 (.X(n628), 
	.C(n1472), 
	.B(n560), 
	.A2(n1474), 
	.A1(n1475));
   SEN_INV_S_4 U2102 (.X(n1202), 
	.A(n1248));
   SEN_ND2_1P5 U2103 (.X(n1149), 
	.A2(pprow1_qual[7]), 
	.A1(pprow1_qual[9]));
   SEN_OAOI211_8 U2104 (.X(n1813), 
	.C(n1792), 
	.B(n1793), 
	.A2(pprow6_qual[15]), 
	.A1(pprow7_qual[13]));
   SEN_AOAI211_8 U2105 (.X(n1608), 
	.C(n1556), 
	.B(n1557), 
	.A2(n1558), 
	.A1(n1559));
   SEN_EN2_1 U2106 (.X(n1561), 
	.A2(n1557), 
	.A1(n732));
   SEN_NR2_S_2 U2107 (.X(n509), 
	.A2(n511), 
	.A1(n510));
   SEN_NR2_T_4 U2108 (.X(n439), 
	.A2(net83157), 
	.A1(net83071));
   SEN_INV_S_0P5 U2109 (.X(n448), 
	.A(n443));
   SEN_INV_S_1 U2110 (.X(n449), 
	.A(pprow0_qual[7]));
   SEN_BUF_6 U2111 (.X(net84730), 
	.A(C[7]));
   SEN_ND2_2 U2112 (.X(n442), 
	.A2(pprow0_qual[6]), 
	.A1(C[6]));
   SEN_ND2_2 U2113 (.X(net84118), 
	.A2(net84150), 
	.A1(n442));
   SEN_OAI211_4 U2114 (.X(net84354), 
	.B2(net84393), 
	.B1(net84392), 
	.A2(net84734), 
	.A1(pprow0_qual[1]));
   SEN_OA2BB2_2 U2115 (.X(net84409), 
	.B2(net94287), 
	.B1(net84418), 
	.A2(net84417), 
	.A1(net84392));
   SEN_INV_S_1 U2116 (.X(n451), 
	.A(pprow0_qual[5]));
   SEN_EO2_S_0P5 U2117 (.X(net84407), 
	.A2(C[5]), 
	.A1(n451));
   SEN_ND2_4 U2118 (.X(net84357), 
	.A2(net84414), 
	.A1(net84384));
   SEN_BUF_S_1 U2119 (.X(net84636), 
	.A(\bmul/neg10 ));
   SEN_NR2_S_4 U2120 (.X(n455), 
	.A2(net2268), 
	.A1(n454));
   SEN_ND2_T_2 U2121 (.X(net87761), 
	.A2(net86213), 
	.A1(net83833));
   SEN_INV_0P65 U2122 (.X(net84232), 
	.A(net84150));
   SEN_AOI21B_4 U2123 (.X(net83459), 
	.B(net83299), 
	.A2(n268), 
	.A1(n1245));
   SEN_ND2B_3 U2124 (.X(n641), 
	.B(net87763), 
	.A(net87762));
   SEN_AOI31_3 U2125 (.X(net84408), 
	.B(net84412), 
	.A3(net84411), 
	.A2(net84410), 
	.A1(net84409));
   SEN_AN2_3 U2126 (.X(n663), 
	.A2(n248), 
	.A1(n1743));
   SEN_OAI21_S_1 U2127 (.X(net83919), 
	.B(n260), 
	.A2(n1046), 
	.A1(n521));
   SEN_ND2_2 U2128 (.X(net82193), 
	.A2(net82516), 
	.A1(net82515));
   SEN_EO2_2 U2129 (.X(n937), 
	.A2(n935), 
	.A1(n936));
   SEN_ND3B_2 U2130 (.X(n935), 
	.B2(\bmul/neg4 ), 
	.B1(pprow2_qual[1]), 
	.A(n934));
   SEN_OAOI211_0P5 U2131 (.X(n464), 
	.C(n894), 
	.B(n895), 
	.A2(n896), 
	.A1(n258));
   SEN_EN2_DG_4 U2132 (.X(net83534), 
	.A2(n461), 
	.A1(net83461));
   SEN_ND2_S_3 U2133 (.X(n1010), 
	.A2(n965), 
	.A1(n966));
   SEN_AO21B_1 U2134 (.X(n986), 
	.B(net83814), 
	.A2(net83817), 
	.A1(n984));
   SEN_NR3_G_1 U2135 (.X(net83496), 
	.A3(n1225), 
	.A2(net82970), 
	.A1(n1226));
   SEN_ND2B_S_4 U2136 (.X(n1311), 
	.B(n1219), 
	.A(pprow4_qual[7]));
   SEN_ND2_S_0P5 U2137 (.X(n907), 
	.A2(n926), 
	.A1(n925));
   SEN_AOI22_T_6 U2138 (.X(net82098), 
	.B2(pprow2_qual[23]), 
	.B1(pprow3_qual[21]), 
	.A2(n1800), 
	.A1(n1799));
   SEN_EO2_3 U2139 (.X(net82982), 
	.A2(net90917), 
	.A1(n710));
   SEN_INV_2 U2140 (.X(n975), 
	.A(n976));
   SEN_OR2_10 U2141 (.X(n1175), 
	.A2(pprow5_qual[3]), 
	.A1(pprow4_qual[5]));
   SEN_EO2_2 U2142 (.X(Z[29]), 
	.A2(net82321), 
	.A1(net82320));
   SEN_AO31_2 U2143 (.X(net86258), 
	.B(net83570), 
	.A3(net83572), 
	.A2(net83777), 
	.A1(n1135));
   SEN_ND2B_6 U2144 (.X(net82768), 
	.B(pprow10_qual[1]), 
	.A(net82973));
   SEN_INV_2 U2145 (.X(n982), 
	.A(n980));
   SEN_EO2_2 U2146 (.X(n980), 
	.A2(n948), 
	.A1(n949));
   SEN_AOAI211_6 U2147 (.X(n1730), 
	.C(n1726), 
	.B(n1727), 
	.A2(n1728), 
	.A1(n1729));
   SEN_NR2_6 U2148 (.X(n1396), 
	.A2(n578), 
	.A1(n577));
   SEN_INV_S_3 U2149 (.X(net84201), 
	.A(pprow2_qual[4]));
   SEN_AO21B_1 U2150 (.X(net85984), 
	.B(net84006), 
	.A2(net86076), 
	.A1(net84650));
   SEN_INV_8 U2151 (.X(n485), 
	.A(net83954));
   SEN_NR2_S_4 U2152 (.X(n501), 
	.A2(net82582), 
	.A1(net82581));
   SEN_OAI21_S_8 U2153 (.X(n493), 
	.B(n500), 
	.A2(n499), 
	.A1(net82583));
   SEN_INV_S_6 U2154 (.X(n499), 
	.A(net82586));
   SEN_ND2_4 U2155 (.X(net83578), 
	.A2(pprow3_qual[3]), 
	.A1(pprow2_qual[5]));
   SEN_INV_1P5 U2156 (.X(n504), 
	.A(pprow3_qual[3]));
   SEN_INV_1 U2157 (.X(n503), 
	.A(pprow2_qual[5]));
   SEN_EO2_S_0P5 U2158 (.X(net85880), 
	.A2(pprow3_qual[3]), 
	.A1(pprow2_qual[5]));
   SEN_AO21B_1 U2159 (.X(net86455), 
	.B(net82586), 
	.A2(net82674), 
	.A1(net82583));
   SEN_EO2_0P5 U2160 (.X(net84246), 
	.A2(n513), 
	.A1(n511));
   SEN_ND2B_4 U2162 (.X(net84384), 
	.B(n872), 
	.A(C[4]));
   SEN_INV_0P8 U2163 (.X(net83829), 
	.A(pprow0_qual[14]));
   SEN_AOAI211_8 U2164 (.X(n1376), 
	.C(n1340), 
	.B(n1341), 
	.A2(n1342), 
	.A1(n1343));
   SEN_EN2_DG_1 U2165 (.X(n1231), 
	.A2(n814), 
	.A1(pprow8_qual[0]));
   SEN_EO2_1 U2166 (.X(n709), 
	.A2(pprow5_qual[0]), 
	.A1(pprow4_qual[2]));
   SEN_AOAI211_6 U2167 (.X(net82137), 
	.C(n1778), 
	.B(n1779), 
	.A2(n1780), 
	.A1(n1781));
   SEN_INV_1 U2168 (.X(net83796), 
	.A(net83798));
   SEN_EN2_DG_1 U2169 (.X(n949), 
	.A2(n956), 
	.A1(n104));
   SEN_ND2_4 U2170 (.X(n516), 
	.A2(n133), 
	.A1(n518));
   SEN_EO2_0P5 U2171 (.X(n862), 
	.A2(n866), 
	.A1(C[3]));
   SEN_ND2_T_2 U2172 (.X(n879), 
	.A2(pprow0_qual[3]), 
	.A1(C[3]));
   SEN_ND2_G_1 U2173 (.X(n965), 
	.A2(pprow1_qual[7]), 
	.A1(pprow1_qual[5]));
   SEN_BUF_1 U2174 (.X(n521), 
	.A(n1047));
   SEN_EO2_DG_1 U2175 (.X(n725), 
	.A2(n533), 
	.A1(pprow1_qual[7]));
   SEN_BUF_1 U2176 (.X(n524), 
	.A(C[4]));
   SEN_ND3_T_4 U2177 (.X(n1199), 
	.A3(n906), 
	.A2(n903), 
	.A1(n902));
   SEN_BUF_1 U2178 (.X(n525), 
	.A(pprow1_qual[16]));
   SEN_ND2_T_1P5 U2179 (.X(n1275), 
	.A2(n1153), 
	.A1(n1223));
   SEN_INV_0P8 U2180 (.X(net84449), 
	.A(net84437));
   SEN_INV_3 U2181 (.X(n876), 
	.A(pprow1_qual[1]));
   SEN_BUF_1 U2182 (.X(n527), 
	.A(pprow1_qual[6]));
   SEN_ND2B_V1_2 U2183 (.X(n1154), 
	.B(n702), 
	.A(n1192));
   SEN_INV_S_0P5 U2185 (.X(n528), 
	.A(n904));
   SEN_ND2_0P5 U2186 (.X(n1329), 
	.A2(pprow9_qual[0]), 
	.A1(pprow8_qual[2]));
   SEN_INV_S_0P5 U2187 (.X(n530), 
	.A(n922));
   SEN_ND2_G_1 U2188 (.X(n1237), 
	.A2(pprow7_qual[2]), 
	.A1(pprow6_qual[4]));
   SEN_INV_3 U2189 (.X(n1059), 
	.A(n1191));
   SEN_ND2_G_2 U2190 (.X(n1191), 
	.A2(pprow1_qual[9]), 
	.A1(pprow1_qual[11]));
   SEN_AO21B_8 U2191 (.X(n1469), 
	.B(n1404), 
	.A2(n532), 
	.A1(n1403));
   SEN_INV_S_0P5 U2192 (.X(n533), 
	.A(n942));
   SEN_INV_S_0P5 U2193 (.X(n534), 
	.A(n1021));
   SEN_INV_0P65 U2194 (.X(n960), 
	.A(n1197));
   SEN_ND2B_4 U2195 (.X(n923), 
	.B(n1197), 
	.A(n291));
   SEN_AOI21_G_1 U2196 (.X(n1111), 
	.B(n1152), 
	.A2(n780), 
	.A1(n620));
   SEN_INV_S_6 U2197 (.X(n1152), 
	.A(n1151));
   SEN_INV_4 U2198 (.X(n1461), 
	.A(n1581));
   SEN_AOAI211_3 U2199 (.X(net82071), 
	.C(net82182), 
	.B(net90615), 
	.A2(net82181), 
	.A1(net82180));
   SEN_EO2_DG_1 U2200 (.X(net86279), 
	.A2(n1436), 
	.A1(net82876));
   SEN_INV_S_1 U2201 (.X(net90884), 
	.A(net83684));
   SEN_INV_S_0P5 U2202 (.X(net90880), 
	.A(net84047));
   SEN_EO2_DG_1 U2203 (.X(net86010), 
	.A2(pprow1_qual[14]), 
	.A1(n525));
   SEN_INV_0P8 U2204 (.X(net84271), 
	.A(net84220));
   SEN_INV_S_0P5 U2205 (.X(n542), 
	.A(n946));
   SEN_EN2_S_1 U2206 (.X(n543), 
	.A2(n738), 
	.A1(n737));
   SEN_EN2_DG_1 U2207 (.X(n727), 
	.A2(n944), 
	.A1(C[9]));
   SEN_EN2_S_2 U2208 (.X(n955), 
	.A2(n953), 
	.A1(n954));
   SEN_OA21_2 U2209 (.X(net86698), 
	.B(net84150), 
	.A2(net84157), 
	.A1(net84156));
   SEN_AO21B_4 U2210 (.X(n544), 
	.B(n978), 
	.A2(n979), 
	.A1(net84111));
   SEN_ND2_S_0P5 U2211 (.X(n545), 
	.A2(n1022), 
	.A1(n1109));
   SEN_ND2_S_0P8 U2212 (.X(n780), 
	.A2(n551), 
	.A1(n545));
   SEN_AN2_S_0P5 U2213 (.X(n1060), 
	.A2(n545), 
	.A1(n551));
   SEN_AOI21B_1 U2214 (.X(n1250), 
	.B(n1281), 
	.A2(n1249), 
	.A1(n1270));
   SEN_AO21B_4 U2215 (.X(net84147), 
	.B(net84152), 
	.A2(net84239), 
	.A1(net84238));
   SEN_ND3_T_4 U2216 (.X(n1216), 
	.A3(n766), 
	.A2(n812), 
	.A1(n1215));
   SEN_ND2_S_0P5 U2218 (.X(n777), 
	.A2(n542), 
	.A1(net84221));
   SEN_INV_S_0P5 U2219 (.X(net90815), 
	.A(n202));
   SEN_INV_4 U2220 (.X(n1088), 
	.A(pprow3_qual[5]));
   SEN_EO2_DG_1 U2221 (.X(n752), 
	.A2(pprow3_qual[5]), 
	.A1(pprow2_qual[7]));
   SEN_ND2_G_1 U2222 (.X(net84046), 
	.A2(n1016), 
	.A1(n1041));
   SEN_EN2_S_1 U2223 (.X(n1014), 
	.A2(n1012), 
	.A1(n1042));
   SEN_INV_1 U2224 (.X(net83197), 
	.A(net83189));
   SEN_AOI31_0P5 U2225 (.X(net82932), 
	.B(n1458), 
	.A3(n1459), 
	.A2(net82941), 
	.A1(n2040));
   SEN_INV_2 U2226 (.X(net90705), 
	.A(net90704));
   SEN_EO2_8 U2227 (.X(n1811), 
	.A2(net90746), 
	.A1(net82161));
   SEN_OR2_2P5 U2228 (.X(n586), 
	.A2(n1724), 
	.A1(n1723));
   SEN_OR4B_4 U2229 (.X(n559), 
	.B3(n1433), 
	.B2(n1434), 
	.B1(n1435), 
	.A(n1432));
   SEN_AN2_DG_3 U2230 (.X(n570), 
	.A2(net84233), 
	.A1(n929));
   SEN_INV_0P65 U2231 (.X(n929), 
	.A(n928));
   SEN_INV_S_1 U2232 (.X(n1070), 
	.A(n1105));
   SEN_BUF_1 U2233 (.X(net90615), 
	.A(net95872));
   SEN_ND3_S_8 U2234 (.X(n1075), 
	.A3(n811), 
	.A2(n1045), 
	.A1(n1047));
   SEN_ND2_3 U2235 (.X(n1240), 
	.A2(pprow5_qual[4]), 
	.A1(pprow4_qual[6]));
   SEN_OR2_5 U2236 (.X(n650), 
	.A2(net84004), 
	.A1(net84003));
   SEN_OR2_5 U2237 (.X(net84008), 
	.A2(pprow2_qual[2]), 
	.A1(pprow3_qual[0]));
   SEN_INV_2 U2238 (.X(n647), 
	.A(n646));
   SEN_BUF_1 U2239 (.X(n551), 
	.A(n1107));
   SEN_NR2B_V1DG_3 U2240 (.X(n1099), 
	.B(net83677), 
	.A(net83685));
   SEN_NR2B_4 U2241 (.X(n1194), 
	.B(n1193), 
	.A(n291));
   SEN_ND2_2 U2242 (.X(n963), 
	.A2(n961), 
	.A1(n996));
   SEN_OAI21_G_4 U2243 (.X(n1292), 
	.B(n1256), 
	.A2(net83431), 
	.A1(n1257));
   SEN_INV_4 U2244 (.X(n1257), 
	.A(n1255));
   SEN_ND2_G_0P65 U2245 (.X(n1256), 
	.A2(pprow0_qual[18]), 
	.A1(C[18]));
   SEN_ND2_T_2 U2247 (.X(n1182), 
	.A2(n1240), 
	.A1(n1241));
   SEN_OA21_1 U2248 (.X(n669), 
	.B(n526), 
	.A2(n537), 
	.A1(n1272));
   SEN_INV_S_3 U2249 (.X(n1232), 
	.A(n2051));
   SEN_ND2_2 U2250 (.X(n1229), 
	.A2(n1227), 
	.A1(n2051));
   SEN_NR2B_4 U2251 (.X(net86076), 
	.B(net84009), 
	.A(net84008));
   SEN_AO21B_4 U2252 (.X(n1359), 
	.B(n1353), 
	.A2(n774), 
	.A1(n1281));
   SEN_OAI21_S_8 U2253 (.X(n1560), 
	.B(n1509), 
	.A2(n1510), 
	.A1(n1511));
   SEN_ND4_2 U2254 (.X(net83152), 
	.A4(net83166), 
	.A3(net83203), 
	.A2(net83204), 
	.A1(net83205));
   SEN_OAI21_S_3 U2256 (.X(n1605), 
	.B(n1649), 
	.A2(n1650), 
	.A1(n18));
   SEN_AOAI211_6 U2257 (.X(net82070), 
	.C(n1772), 
	.B(n1773), 
	.A2(net91564), 
	.A1(n1774));
   SEN_OR2_1 U2258 (.X(n769), 
	.A2(pprow1_qual[3]), 
	.A1(pprow1_qual[5]));
   SEN_OR2_5 U2259 (.X(n1382), 
	.A2(n1346), 
	.A1(n1345));
   SEN_EO2_DG_2 U2261 (.X(n1507), 
	.A2(n1499), 
	.A1(n718));
   SEN_EO2_0P5 U2262 (.X(n653), 
	.A2(net82824), 
	.A1(net82823));
   SEN_EN2_0P5 U2263 (.X(n873), 
	.A2(n44), 
	.A1(n881));
   SEN_AOI311_4 U2264 (.X(n1039), 
	.B2(net83989), 
	.B1(n1036), 
	.A3(n383), 
	.A2(n1037), 
	.A1(n1038));
   SEN_ND2_2 U2265 (.X(n928), 
	.A2(n259), 
	.A1(n621));
   SEN_AN2_2 U2267 (.X(n662), 
	.A2(n1438), 
	.A1(n1439));
   SEN_ND2B_6 U2268 (.X(net83094), 
	.B(net83105), 
	.A(net83096));
   SEN_EO2_2 U2269 (.X(n1406), 
	.A2(n715), 
	.A1(n1403));
   SEN_INV_S_1P5 U2270 (.X(n1610), 
	.A(n1614));
   SEN_EO2_2 U2271 (.X(n684), 
	.A2(n1387), 
	.A1(n1386));
   SEN_EN2_DG_1 U2272 (.X(Z[5]), 
	.A2(n874), 
	.A1(n875));
   SEN_INV_S_2 U2273 (.X(n603), 
	.A(n1383));
   SEN_INV_2 U2274 (.X(n1365), 
	.A(n1290));
   SEN_NR2_1 U2275 (.X(n1294), 
	.A2(n1290), 
	.A1(n1291));
   SEN_NR2_S_0P65 U2276 (.X(n1395), 
	.A2(n1430), 
	.A1(n1393));
   SEN_INV_S_6 U2277 (.X(n1079), 
	.A(n1075));
   SEN_ND2_S_1 U2278 (.X(n1267), 
	.A2(n120), 
	.A1(net83397));
   SEN_EO2_0P5 U2279 (.X(n657), 
	.A2(n1456), 
	.A1(n1457));
   SEN_ND2_S_0P5 U2280 (.X(n1458), 
	.A2(net82839), 
	.A1(net82843));
   SEN_EN2_DG_1 U2281 (.X(n1121), 
	.A2(n668), 
	.A1(n260));
   SEN_EO2_S_1 U2283 (.X(n1664), 
	.A2(n1655), 
	.A1(n1656));
   SEN_OR2_10 U2284 (.X(net82703), 
	.A2(n109), 
	.A1(n644));
   SEN_AO21B_4 U2285 (.X(net83816), 
	.B(n950), 
	.A2(n952), 
	.A1(n951));
   SEN_INV_S_3 U2286 (.X(n944), 
	.A(pprow0_qual[9]));
   SEN_ND2_G_4 U2287 (.X(n1101), 
	.A2(pprow6_qual[0]), 
	.A1(pprow6_qual[1]));
   SEN_AO21B_2 U2289 (.X(n1053), 
	.B(net83571), 
	.A2(net83891), 
	.A1(net83960));
   SEN_EO2_3 U2290 (.X(n1474), 
	.A2(n1469), 
	.A1(n713));
   SEN_ND2_6 U2291 (.X(net84009), 
	.A2(pprow2_qual[0]), 
	.A1(pprow2_qual[1]));
   SEN_ND2_S_4 U2292 (.X(n1673), 
	.A2(n1672), 
	.A1(net82503));
   SEN_OA21_2 U2293 (.X(n629), 
	.B(net83552), 
	.A2(n1128), 
	.A1(net83796));
   SEN_EO2_S_3 U2294 (.X(n1047), 
	.A2(n1039), 
	.A1(n1040));
   SEN_OA2BB2_8 U2295 (.X(n1640), 
	.B2(n561), 
	.B1(n1599), 
	.A2(n1601), 
	.A1(n1600));
   SEN_ND4B_4 U2296 (.X(n1248), 
	.B3(n1189), 
	.B2(n1190), 
	.B1(n620), 
	.A(n1192));
   SEN_INV_S_3 U2297 (.X(n1273), 
	.A(n1189));
   SEN_ND2_G_1 U2298 (.X(n1189), 
	.A2(pprow1_qual[11]), 
	.A1(pprow1_qual[13]));
   SEN_AOI21B_8 U2299 (.X(n1807), 
	.B(net82210), 
	.A2(net82209), 
	.A1(n1805));
   SEN_EN2_S_6 U2300 (.X(net83954), 
	.A2(n1032), 
	.A1(n724));
   SEN_INV_1P5 U2301 (.X(n1046), 
	.A(n1041));
   SEN_EN2_0P5 U2302 (.X(n691), 
	.A2(n161), 
	.A1(n1614));
   SEN_INV_S_0P5 U2304 (.X(net89933), 
	.A(n85));
   SEN_EN3_6 U2306 (.X(n1735), 
	.A3(n1733), 
	.A2(n1732), 
	.A1(n422));
   SEN_AOI21B_1 U2307 (.X(n931), 
	.B(net84271), 
	.A2(net84218), 
	.A1(net97377));
   SEN_OA21_2 U2308 (.X(net86699), 
	.B(net84414), 
	.A2(n204), 
	.A1(net84435));
   SEN_INV_S_0P5 U2309 (.X(net83640), 
	.A(pprow0_qual[16]));
   SEN_INV_S_1 U2310 (.X(net82855), 
	.A(net82859));
   SEN_INV_S_6 U2311 (.X(net82856), 
	.A(net85257));
   SEN_ND2_T_2 U2312 (.X(net82821), 
	.A2(net87814), 
	.A1(net87813));
   SEN_INV_S_0P5 U2313 (.X(net82820), 
	.A(net82640));
   SEN_ND2_T_8 U2314 (.X(n1463), 
	.A2(net83025), 
	.A1(n468));
   SEN_INV_S_0P5 U2315 (.X(n569), 
	.A(n1206));
   SEN_EO2_2 U2316 (.X(n1523), 
	.A2(n256), 
	.A1(n747));
   SEN_ND2_S_3 U2317 (.X(net82125), 
	.A2(n1787), 
	.A1(n1786));
   SEN_OR2_5 U2318 (.X(n999), 
	.A2(pprow1_qual[4]), 
	.A1(pprow1_qual[6]));
   SEN_EO2_2 U2319 (.X(n1525), 
	.A2(n1572), 
	.A1(n1574));
   SEN_EO3_DG_1 U2320 (.X(n985), 
	.A3(n30), 
	.A2(n33), 
	.A1(n1038));
   SEN_AOI21B_2 U2321 (.X(net83176), 
	.B(n1427), 
	.A2(n1369), 
	.A1(net86332));
   SEN_ND2B_V1DG_2 U2322 (.X(n1124), 
	.B(n1123), 
	.A(n1127));
   SEN_INV_0P8 U2323 (.X(n1044), 
	.A(n1042));
   SEN_ND4B_8 U2324 (.X(net82583), 
	.B3(n536), 
	.B2(n1585), 
	.B1(n1584), 
	.A(n1586));
   SEN_ND2_3 U2325 (.X(n1518), 
	.A2(n1415), 
	.A1(n1416));
   SEN_INV_2 U2326 (.X(n1417), 
	.A(n1518));
   SEN_EN3_6 U2327 (.X(net82207), 
	.A3(n1804), 
	.A2(n1803), 
	.A1(n1802));
   SEN_EO3_DG_1 U2328 (.X(Z[9]), 
	.A3(n950), 
	.A2(n952), 
	.A1(n951));
   SEN_AOAI211_8 U2329 (.X(net82167), 
	.C(n1788), 
	.B(net82260), 
	.A2(n1789), 
	.A1(n1790));
   SEN_EO2_0P5 U2330 (.X(n676), 
	.A2(n1450), 
	.A1(n1452));
   SEN_OAI21_S_8 U2331 (.X(net82349), 
	.B(net82460), 
	.A2(n1702), 
	.A1(n1701));
   SEN_OA21_4 U2332 (.X(n703), 
	.B(n1307), 
	.A2(n1308), 
	.A1(n211));
   SEN_INV_1 U2333 (.X(n1526), 
	.A(n1528));
   SEN_ND2_2 U2334 (.X(n1281), 
	.A2(n1223), 
	.A1(net83359));
   SEN_AOI31_3 U2335 (.X(n1243), 
	.B(n1310), 
	.A3(n1311), 
	.A2(n1242), 
	.A1(n1312));
   SEN_OAI221_2 U2336 (.X(n1090), 
	.C(net83571), 
	.B2(n1088), 
	.B1(net83574), 
	.A2(n1089), 
	.A1(net83574));
   SEN_ND2_3 U2337 (.X(n1151), 
	.A2(n1109), 
	.A1(n1203));
   SEN_AOAI211_2 U2338 (.X(n1551), 
	.C(n1594), 
	.B(n1550), 
	.A2(n1593), 
	.A1(net102542));
   SEN_OAI211_2 U2339 (.X(n1247), 
	.B2(n1008), 
	.B1(n1007), 
	.A2(n1009), 
	.A1(n1010));
   SEN_ND2_S_4 U2340 (.X(n1180), 
	.A2(n1082), 
	.A1(n1083));
   SEN_EO2_2 U2341 (.X(Z[22]), 
	.A2(n658), 
	.A1(n657));
   SEN_AO21B_2 U2342 (.X(n658), 
	.B(net82845), 
	.A2(net82843), 
	.A1(n1399));
   SEN_OR2_2P5 U2343 (.X(net83581), 
	.A2(pprow3_qual[6]), 
	.A1(pprow2_qual[8]));
   SEN_INV_0P65 U2344 (.X(net84148), 
	.A(net84118));
   SEN_AOI21B_1 U2345 (.X(net83019), 
	.B(n1579), 
	.A2(n1583), 
	.A1(n1463));
   SEN_AOAI211_8 U2346 (.X(net82091), 
	.C(n1801), 
	.B(n1802), 
	.A2(n1803), 
	.A1(n1804));
   SEN_AN2_DG_1 U2347 (.X(n578), 
	.A2(n1394), 
	.A1(n1429));
   SEN_INV_0P8 U2348 (.X(net84471), 
	.A(pprow0_qual[1]));
   SEN_INV_S_0P5 U2349 (.X(n587), 
	.A(n742));
   SEN_INV_0P5 U2350 (.X(n593), 
	.A(n1117));
   SEN_ND2_S_1 U2351 (.X(n598), 
	.A2(n1554), 
	.A1(n1555));
   SEN_ND2_T_2 U2352 (.X(n599), 
	.A2(n597), 
	.A1(n596));
   SEN_ND2_T_1 U2353 (.X(Z[25]), 
	.A2(n599), 
	.A1(n598));
   SEN_INV_2 U2354 (.X(n597), 
	.A(n1554));
   SEN_INV_2 U2355 (.X(n601), 
	.A(n600));
   SEN_NR2B_V1_1 U2356 (.X(n1071), 
	.B(n1106), 
	.A(net83862));
   SEN_BUF_S_1 U2357 (.X(n605), 
	.A(n790));
   SEN_BUF_S_1 U2358 (.X(n606), 
	.A(\bmul/two6 ));
   SEN_BUF_S_1 U2359 (.X(n607), 
	.A(\bmul/two5 ));
   SEN_BUF_6 U2360 (.X(n812), 
	.A(\bmul/neg7 ));
   SEN_BUF_S_1 U2361 (.X(n608), 
	.A(n819));
   SEN_BUF_S_1 U2362 (.X(n609), 
	.A(n791));
   SEN_BUF_S_1 U2363 (.X(n610), 
	.A(n789));
   SEN_BUF_S_1 U2364 (.X(n611), 
	.A(\bmul/one7 ));
   SEN_EO2_S_0P5 U2365 (.X(\bmul/one7 ), 
	.A2(n811), 
	.A1(A[14]));
   SEN_BUF_S_1 U2366 (.X(n811), 
	.A(\bmul/neg6 ));
   SEN_BUF_S_1 U2367 (.X(n612), 
	.A(\bmul/one6 ));
   SEN_BUF_S_1 U2368 (.X(n613), 
	.A(\bmul/one5 ));
   SEN_INV_S_0P5 U2369 (.X(n614), 
	.A(\bmul/neg4 ));
   SEN_INV_S_1 U2370 (.X(n615), 
	.A(n782));
   SEN_EO2_DG_8 U2371 (.X(n618), 
	.A2(pprow3_qual[6]), 
	.A1(pprow2_qual[8]));
   SEN_INV_S_2 U2372 (.X(n620), 
	.A(n1059));
   SEN_ND2_2 U2373 (.X(net83572), 
	.A2(pprow3_qual[6]), 
	.A1(pprow2_qual[8]));
   SEN_INV_2 U2374 (.X(net87821), 
	.A(net84286));
   SEN_NR2_S_2 U2375 (.X(net84284), 
	.A2(net84237), 
	.A1(n928));
   SEN_ND2_2 U2376 (.X(net87814), 
	.A2(n667), 
	.A1(n624));
   SEN_INV_1 U2377 (.X(n625), 
	.A(n667));
   SEN_INV_S_2 U2378 (.X(net82823), 
	.A(net82821));
   SEN_ND2_2 U2379 (.X(n1305), 
	.A2(n636), 
	.A1(net83295));
   SEN_EO2_2 U2380 (.X(n636), 
	.A2(n1243), 
	.A1(n1244));
   SEN_ND2_S_0P8 U2382 (.X(n634), 
	.A2(n633), 
	.A1(n943));
   SEN_ND2_2 U2383 (.X(net84221), 
	.A2(n635), 
	.A1(n634));
   SEN_INV_0P8 U2384 (.X(n632), 
	.A(n943));
   SEN_INV_0P5 U2385 (.X(n633), 
	.A(n725));
   SEN_INV_2 U2386 (.X(net84223), 
	.A(net84221));
   SEN_AN2_S_0P5 U2387 (.X(n637), 
	.A2(pprow5_qual[2]), 
	.A1(pprow4_qual[4]));
   SEN_INV_S_1 U2388 (.X(net83036), 
	.A(net82901));
   SEN_ND2_G_1 U2389 (.X(net83820), 
	.A2(n987), 
	.A1(n988));
   SEN_INV_1 U2390 (.X(n983), 
	.A(n981));
   SEN_OAI21_G_1 U2391 (.X(n927), 
	.B(n616), 
	.A2(n1002), 
	.A1(n924));
   SEN_ND2_S_0P5 U2392 (.X(net82705), 
	.A2(pprow3_qual[15]), 
	.A1(pprow2_qual[17]));
   SEN_ND2_G_1 U2393 (.X(n1239), 
	.A2(pprow5_qual[5]), 
	.A1(pprow4_qual[7]));
   SEN_ND2_T_0P5 U2394 (.X(n1404), 
	.A2(pprow7_qual[6]), 
	.A1(pprow6_qual[8]));
   SEN_INV_S_1 U2395 (.X(net83359), 
	.A(pprow1_qual[15]));
   SEN_INV_S_0P5 U2397 (.X(net83729), 
	.A(C[15]));
   SEN_INV_S_0P5 U2398 (.X(net83730), 
	.A(pprow0_qual[15]));
   SEN_NR2B_V1_1 U2399 (.X(n1221), 
	.B(n1240), 
	.A(n1311));
   SEN_NR2_S_0P5 U2400 (.X(n1467), 
	.A2(pprow8_qual[5]), 
	.A1(pprow9_qual[3]));
   SEN_INV_1 U2401 (.X(n1641), 
	.A(C[26]));
   SEN_INV_1 U2402 (.X(n1512), 
	.A(pprow2_qual[18]));
   SEN_ND2B_S_0P5 U2403 (.X(net83522), 
	.B(net83640), 
	.A(C[16]));
   SEN_INV_1 U2404 (.X(n1513), 
	.A(pprow3_qual[16]));
   SEN_ND2_S_0P5 U2405 (.X(net83612), 
	.A2(n1172), 
	.A1(n1230));
   SEN_ND2_S_0P5 U2406 (.X(n1172), 
	.A2(n1170), 
	.A1(n1171));
   SEN_INV_S_0P5 U2407 (.X(n1170), 
	.A(n1169));
   SEN_INV_S_1 U2408 (.X(n1642), 
	.A(pprow0_qual[26]));
   SEN_ND2_S_0P5 U2409 (.X(n1755), 
	.A2(pprow11_qual[4]), 
	.A1(pprow10_qual[6]));
   SEN_ND2_G_1 U2410 (.X(n1778), 
	.A2(n1776), 
	.A1(n1777));
   SEN_INV_1 U2411 (.X(n886), 
	.A(n888));
   SEN_INV_S_1 U2412 (.X(n1703), 
	.A(C[27]));
   SEN_AN2_S_0P5 U2413 (.X(n1400), 
	.A2(pprow9_qual[2]), 
	.A1(pprow8_qual[4]));
   SEN_EO2_S_0P5 U2414 (.X(n649), 
	.A2(pprow3_qual[13]), 
	.A1(pprow2_qual[15]));
   SEN_ND2_S_0P5 U2415 (.X(n1500), 
	.A2(pprow7_qual[7]), 
	.A1(pprow6_qual[9]));
   SEN_ND2_S_0P5 U2416 (.X(n984), 
	.A2(net83815), 
	.A1(net83816));
   SEN_INV_S_1 U2417 (.X(n917), 
	.A(n921));
   SEN_ND2_S_0P65 U2418 (.X(n1016), 
	.A2(n1014), 
	.A1(n1015));
   SEN_AOAI211_0P5 U2419 (.X(n1127), 
	.C(n1143), 
	.B(pprow6_qual[1]), 
	.A2(pprow6_qual[0]), 
	.A1(n437));
   SEN_INV_S_0P5 U2420 (.X(n1683), 
	.A(pprow9_qual[7]));
   SEN_EO2_2 U2421 (.X(net82141), 
	.A2(n734), 
	.A1(net82125));
   SEN_INV_S_1 U2422 (.X(n1502), 
	.A(pprow6_qual[10]));
   SEN_EN2_S_1 U2423 (.X(n1304), 
	.A2(n1243), 
	.A1(n1244));
   SEN_ND2_G_1 U2424 (.X(net82508), 
	.A2(net82511), 
	.A1(net82510));
   SEN_NR2_S_0P5 U2425 (.X(n1434), 
	.A2(n1425), 
	.A1(n1426));
   SEN_INV_S_1 U2427 (.X(n913), 
	.A(n891));
   SEN_ND2_S_1 U2428 (.X(n1565), 
	.A2(n1512), 
	.A1(n1513));
   SEN_EO2_S_0P5 U2429 (.X(\bmul/one10 ), 
	.A2(n814), 
	.A1(A[20]));
   SEN_EO2_2 U2430 (.X(net83506), 
	.A2(n722), 
	.A1(n1224));
   SEN_INV_0P65 U2431 (.X(n1369), 
	.A(n1430));
   SEN_INV_S_0P5 U2432 (.X(n1757), 
	.A(pprow11_qual[4]));
   SEN_INV_S_0P5 U2433 (.X(net82525), 
	.A(n23));
   SEN_EO2_DG_1 U2434 (.X(n1741), 
	.A2(n1696), 
	.A1(n1744));
   SEN_EN2_0P5 U2435 (.X(n932), 
	.A2(n542), 
	.A1(net84223));
   SEN_NR2_S_1 U2436 (.X(n1072), 
	.A2(n1070), 
	.A1(n1071));
   SEN_INV_S_0P5 U2437 (.X(net84146), 
	.A(net84108));
   SEN_INV_1 U2438 (.X(n1503), 
	.A(n1500));
   SEN_OR3B_0P5 U2439 (.X(n908), 
	.B2(n1002), 
	.B1(n924), 
	.A(n907));
   SEN_ND2_G_1 U2440 (.X(net82706), 
	.A2(pprow2_qual[18]), 
	.A1(pprow3_qual[16]));
   SEN_EO2_S_0P5 U2441 (.X(n708), 
	.A2(pprow5_qual[9]), 
	.A1(pprow4_qual[11]));
   SEN_EO2_S_0P5 U2442 (.X(n1140), 
	.A2(pprow5_qual[4]), 
	.A1(pprow4_qual[6]));
   SEN_EO2_S_0P5 U2443 (.X(n716), 
	.A2(pprow7_qual[2]), 
	.A1(pprow6_qual[4]));
   SEN_EO2_S_0P5 U2444 (.X(n1116), 
	.A2(C[15]), 
	.A1(net83730));
   SEN_INV_S_1 U2445 (.X(n1501), 
	.A(pprow7_qual[8]));
   SEN_EO2_S_0P5 U2446 (.X(n1495), 
	.A2(C[24]), 
	.A1(n1541));
   SEN_INV_S_0P5 U2447 (.X(n1492), 
	.A(n1543));
   SEN_ND2_0P5 U2448 (.X(n1335), 
	.A2(pprow7_qual[4]), 
	.A1(pprow6_qual[6]));
   SEN_OAI21_G_1 U2449 (.X(n1336), 
	.B(n1334), 
	.A2(pprow6_qual[6]), 
	.A1(pprow7_qual[4]));
   SEN_EO2_S_0P5 U2450 (.X(net83175), 
	.A2(C[21]), 
	.A1(n1392));
   SEN_ND2_S_0P5 U2451 (.X(n1372), 
	.A2(pprow9_qual[1]), 
	.A1(pprow8_qual[3]));
   SEN_NR2B_V1DG_1 U2452 (.X(n1435), 
	.B(n1424), 
	.A(C[22]));
   SEN_OR2_1 U2453 (.X(net82901), 
	.A2(pprow3_qual[14]), 
	.A1(pprow2_qual[16]));
   SEN_EO2_S_0P5 U2454 (.X(n744), 
	.A2(pprow7_qual[4]), 
	.A1(pprow6_qual[6]));
   SEN_ND2B_V1_2 U2455 (.X(n1542), 
	.B(n1541), 
	.A(C[24]));
   SEN_ND2_S_0P5 U2456 (.X(n1226), 
	.A2(n662), 
	.A1(n1263));
   SEN_EO3_DG_1 U2457 (.X(Z[21]), 
	.A3(net83064), 
	.A2(n1397), 
	.A1(n1399));
   SEN_EN2_0P5 U2458 (.X(n668), 
	.A2(n1080), 
	.A1(n1081));
   SEN_INV_S_0P5 U2459 (.X(n1653), 
	.A(n1660));
   SEN_INV_1 U2460 (.X(net84231), 
	.A(net84233));
   SEN_EN3_0P5 U2461 (.X(Z[12]), 
	.A3(net84046), 
	.A2(net90880), 
	.A1(n1017));
   SEN_EO2_1 U2462 (.X(n1027), 
	.A2(n1068), 
	.A1(n1067));
   SEN_ND2B_S_0P5 U2463 (.X(n964), 
	.B(n960), 
	.A(n1195));
   SEN_INV_S_0P5 U2464 (.X(net83889), 
	.A(net83581));
   SEN_INV_S_1 U2465 (.X(n840), 
	.A(n760));
   SEN_INV_S_1 U2466 (.X(n845), 
	.A(n761));
   SEN_INV_S_1 U2467 (.X(n835), 
	.A(n755));
   SEN_INV_S_0P5 U2468 (.X(n1838), 
	.A(n814));
   SEN_INV_S_1 U2469 (.X(n772), 
	.A(n771));
   SEN_INV_S_1 U2470 (.X(n841), 
	.A(n760));
   SEN_ND2_S_0P5 U2471 (.X(n1602), 
	.A2(n1540), 
	.A1(n1630));
   SEN_INV_S_0P5 U2472 (.X(n1538), 
	.A(n1537));
   SEN_INV_S_1 U2473 (.X(n844), 
	.A(n761));
   SEN_BUF_S_1 U2474 (.X(n820), 
	.A(n614));
   SEN_INV_S_1 U2475 (.X(n846), 
	.A(n847));
   SEN_INV_S_1 U2476 (.X(n842), 
	.A(n764));
   SEN_INV_S_1 U2477 (.X(n856), 
	.A(n857));
   SEN_INV_S_1 U2478 (.X(n848), 
	.A(n849));
   SEN_INV_S_1 U2479 (.X(n850), 
	.A(n851));
   SEN_INV_S_1 U2480 (.X(n852), 
	.A(n853));
   SEN_INV_S_1 U2481 (.X(n854), 
	.A(n855));
   SEN_INV_1 U2482 (.X(n1081), 
	.A(n1077));
   SEN_INV_S_1 U2483 (.X(n838), 
	.A(n762));
   SEN_INV_S_1 U2484 (.X(n839), 
	.A(n762));
   SEN_BUF_S_1 U2485 (.X(n818), 
	.A(n1840));
   SEN_INV_S_0P5 U2486 (.X(n1489), 
	.A(n815));
   SEN_BUF_S_1 U2487 (.X(n817), 
	.A(n1839));
   SEN_INV_S_1 U2488 (.X(net84592), 
	.A(net2259));
   SEN_INV_S_0P5 U2489 (.X(n1291), 
	.A(n1366));
   SEN_INV_S_0P5 U2490 (.X(n1841), 
	.A(n811));
   SEN_INV_S_0P5 U2491 (.X(n1393), 
	.A(n1429));
   SEN_ND2B_S_0P5 U2492 (.X(n914), 
	.B(\bmul/neg4 ), 
	.A(n915));
   SEN_INV_S_0P5 U2493 (.X(n1426), 
	.A(n1428));
   SEN_INV_S_0P5 U2494 (.X(n1837), 
	.A(n816));
   SEN_EO2_1 U2495 (.X(net85926), 
	.A2(net82130), 
	.A1(n751));
   SEN_EO2_S_0P5 U2496 (.X(\bmul/one13 ), 
	.A2(n815), 
	.A1(A[26]));
   SEN_NR2_1 U2497 (.X(\bmul/two8 ), 
	.A2(n2029), 
	.A1(\bmul/one8 ));
   SEN_NR2_1 U2498 (.X(\bmul/two5 ), 
	.A2(n2026), 
	.A1(\bmul/one5 ));
   SEN_NR2_1 U2499 (.X(\bmul/two9 ), 
	.A2(n2030), 
	.A1(\bmul/one9 ));
   SEN_NR2_1 U2500 (.X(\bmul/two11 ), 
	.A2(n2032), 
	.A1(\bmul/one11 ));
   SEN_NR2_1 U2501 (.X(\bmul/two6 ), 
	.A2(n2027), 
	.A1(\bmul/one6 ));
   SEN_NR2_1 U2502 (.X(\bmul/two10 ), 
	.A2(n2031), 
	.A1(\bmul/one10 ));
   SEN_NR2_1 U2503 (.X(\bmul/two7 ), 
	.A2(n2028), 
	.A1(\bmul/one7 ));
   SEN_EO2_S_0P5 U2504 (.X(\bmul/one11 ), 
	.A2(net84636), 
	.A1(A[22]));
   SEN_EO2_1 U2505 (.X(n714), 
	.A2(pprow9_qual[1]), 
	.A1(pprow8_qual[3]));
   SEN_INV_S_0P5 U2506 (.X(n1332), 
	.A(pprow8_qual[2]));
   SEN_EN2_0P5 U2507 (.X(n1776), 
	.A2(n1782), 
	.A1(n743));
   SEN_EO2_S_0P5 U2508 (.X(n736), 
	.A2(pprow11_qual[1]), 
	.A1(pprow10_qual[3]));
   SEN_INV_S_1 U2509 (.X(n786), 
	.A(n785));
   SEN_EO2_S_0P5 U2510 (.X(\bmul/one12 ), 
	.A2(net84634), 
	.A1(A[24]));
   SEN_INV_S_0P5 U2511 (.X(n1758), 
	.A(pprow10_qual[6]));
   SEN_ND2_S_0P5 U2512 (.X(n1751), 
	.A2(pprow13_qual[0]), 
	.A1(pprow12_qual[2]));
   SEN_INV_S_0P5 U2513 (.X(n1754), 
	.A(pprow12_qual[2]));
   SEN_INV_S_0P5 U2514 (.X(n1753), 
	.A(pprow13_qual[0]));
   SEN_INV_1 U2515 (.X(net85334), 
	.A(net84025));
   SEN_BUF_S_1 U2516 (.X(n789), 
	.A(B[11]));
   SEN_EO2_S_0P5 U2517 (.X(n756), 
	.A2(pprow5_qual[2]), 
	.A1(pprow4_qual[4]));
   SEN_BUF_S_1 U2518 (.X(n790), 
	.A(B[12]));
   SEN_INV_S_0P5 U2519 (.X(n1316), 
	.A(pprow5_qual[7]));
   SEN_BUF_S_1 U2520 (.X(n791), 
	.A(B[13]));
   SEN_EO2_S_0P5 U2521 (.X(n746), 
	.A2(pprow7_qual[0]), 
	.A1(pprow6_qual[2]));
   SEN_ND2_S_0P5 U2522 (.X(n1634), 
	.A2(pprow11_qual[2]), 
	.A1(pprow10_qual[4]));
   SEN_INV_S_0P5 U2523 (.X(n1636), 
	.A(pprow10_qual[4]));
   SEN_INV_S_0P5 U2524 (.X(n1635), 
	.A(pprow11_qual[2]));
   SEN_ND2B_1 U2525 (.X(n936), 
	.B(\bmul/neg4 ), 
	.A(n933));
   SEN_INV_S_0P5 U2526 (.X(net82972), 
	.A(pprow10_qual[1]));
   SEN_ND2B_2 U2527 (.X(n1366), 
	.B(n1289), 
	.A(C[19]));
   SEN_ND2_S_0P5 U2528 (.X(net82658), 
	.A2(pprow1_qual[21]), 
	.A1(pprow1_qual[23]));
   SEN_INV_S_0P5 U2529 (.X(n892), 
	.A(pprow2_qual[1]));
   SEN_EN2_0P5 U2530 (.X(n2025), 
	.A2(\bmul/neg4 ), 
	.A1(A[8]));
   SEN_ND2_S_0P5 U2531 (.X(n1784), 
	.A2(pprow13_qual[1]), 
	.A1(pprow12_qual[3]));
   SEN_ND2_S_0P5 U2532 (.X(n1425), 
	.A2(pprow0_qual[21]), 
	.A1(C[21]));
   SEN_ND2_S_0P5 U2533 (.X(n1787), 
	.A2(pprow11_qual[5]), 
	.A1(pprow10_qual[7]));
   SEN_ND2_S_0P5 U2534 (.X(n1466), 
	.A2(pprow9_qual[3]), 
	.A1(pprow8_qual[5]));
   SEN_ND2_T_0P5 U2535 (.X(n1637), 
	.A2(pprow12_qual[0]), 
	.A1(n816));
   SEN_INV_S_0P5 U2536 (.X(net84026), 
	.A(pprow0_qual[12]));
   SEN_ND2B_S_2 U2537 (.X(n1367), 
	.B(n1364), 
	.A(C[20]));
   SEN_INV_S_3 U2538 (.X(n1289), 
	.A(pprow0_qual[19]));
   SEN_INV_S_2 U2539 (.X(n1364), 
	.A(pprow0_qual[20]));
   SEN_NR2_S_0P5 U2540 (.X(n767), 
	.A2(pprow6_qual[9]), 
	.A1(pprow7_qual[7]));
   SEN_INV_S_0P5 U2541 (.X(n1234), 
	.A(pprow8_qual[1]));
   SEN_INV_S_1 U2542 (.X(n784), 
	.A(n783));
   SEN_AO22_1 U2543 (.X(n1368), 
	.B2(pprow0_qual[19]), 
	.B1(C[19]), 
	.A2(n1366), 
	.A1(n1292));
   SEN_INV_S_0P5 U2544 (.X(n1315), 
	.A(pprow4_qual[9]));
   SEN_OR2_DG_1 U2545 (.X(n749), 
	.A2(pprow4_qual[11]), 
	.A1(pprow5_qual[9]));
   SEN_ND2_S_0P5 U2547 (.X(net82758), 
	.A2(pprow1_qual[20]), 
	.A1(pprow1_qual[22]));
   SEN_AO22_DG_1 U2548 (.X(n768), 
	.B2(pprow7_qual[8]), 
	.B1(pprow6_qual[10]), 
	.A2(n1504), 
	.A1(n1503));
   SEN_INV_S_1 U2549 (.X(n988), 
	.A(n985));
   SEN_EO3_1 U2550 (.X(Z[13]), 
	.A3(net83919), 
	.A2(n24), 
	.A1(n1074));
   SEN_EO2_S_0P5 U2551 (.X(n655), 
	.A2(n982), 
	.A1(n983));
   SEN_EO2_S_0P5 U2552 (.X(Z[20]), 
	.A2(n1326), 
	.A1(n656));
   SEN_EO2_S_0P5 U2553 (.X(Z[18]), 
	.A2(net83495), 
	.A1(net83494));
   SEN_EN2_S_2 U2554 (.X(n1668), 
	.A2(net82525), 
	.A1(net88079));
   SEN_AO21B_1 U2555 (.X(n1165), 
	.B(n1209), 
	.A2(n659), 
	.A1(net83626));
   SEN_AN2_S_0P5 U2556 (.X(n659), 
	.A2(n1264), 
	.A1(n1263));
   SEN_AO21B_1 U2557 (.X(net83397), 
	.B(n373), 
	.A2(n1437), 
	.A1(n662));
   SEN_AO21B_1 U2558 (.X(n1074), 
	.B(net90993), 
	.A2(net83813), 
	.A1(n1017));
   SEN_ND2_G_1 U2559 (.X(net83814), 
	.A2(n982), 
	.A1(n983));
   SEN_NR2_S_0P5 U2560 (.X(n1459), 
	.A2(net82946), 
	.A1(net82847));
   SEN_INV_S_1 U2561 (.X(n1552), 
	.A(n1550));
   SEN_EO2_S_0P5 U2562 (.X(Z[6]), 
	.A2(n883), 
	.A1(n889));
   SEN_EO2_S_0P5 U2563 (.X(Z[16]), 
	.A2(n673), 
	.A1(n672));
   SEN_AO21B_1 U2564 (.X(n673), 
	.B(n2049), 
	.A2(n1439), 
	.A1(n1165));
   SEN_EN2_0P5 U2565 (.X(Z[17]), 
	.A2(n1212), 
	.A1(net83615));
   SEN_OAI21_G_1 U2566 (.X(n1212), 
	.B(net83617), 
	.A2(n1226), 
	.A1(n1225));
   SEN_INV_S_0P5 U2567 (.X(net83617), 
	.A(net83397));
   SEN_EO2_S_0P5 U2568 (.X(pprow4[5]), 
	.A2(n1898), 
	.A1(n820));
   SEN_AOI22_1 U2569 (.X(n1898), 
	.B2(n773), 
	.B1(n854), 
	.A2(n824), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2570 (.X(pprow4[0]), 
	.A2(n1915), 
	.A1(n820));
   SEN_ND2_G_1 U2571 (.X(n1915), 
	.A2(n773), 
	.A1(n829));
   SEN_EO2_S_0P5 U2572 (.X(pprow4[1]), 
	.A2(n1904), 
	.A1(n820));
   SEN_AOI22_1 U2573 (.X(n1904), 
	.B2(n772), 
	.B1(n846), 
	.A2(n824), 
	.A1(n830));
   SEN_EO2_S_0P5 U2574 (.X(pprow4[2]), 
	.A2(n1901), 
	.A1(n820));
   SEN_AOI22_1 U2575 (.X(n1901), 
	.B2(n772), 
	.B1(n848), 
	.A2(\bmul/two4 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2576 (.X(pprow4[3]), 
	.A2(n1900), 
	.A1(n820));
   SEN_AOI22_1 U2577 (.X(n1900), 
	.B2(n773), 
	.B1(n850), 
	.A2(n824), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2578 (.X(pprow4[4]), 
	.A2(n1899), 
	.A1(n820));
   SEN_AOI22_1 U2579 (.X(n1899), 
	.B2(n773), 
	.B1(n852), 
	.A2(\bmul/two4 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2580 (.X(pprow4[6]), 
	.A2(n1897), 
	.A1(n820));
   SEN_AOI22_1 U2581 (.X(n1897), 
	.B2(n773), 
	.B1(n856), 
	.A2(\bmul/two4 ), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2582 (.X(Z[11]), 
	.A2(n986), 
	.A1(n674));
   SEN_EO2_S_0P5 U2583 (.X(n674), 
	.A2(n987), 
	.A1(n988));
   SEN_EO2_S_0P5 U2584 (.X(Z[15]), 
	.A2(n1165), 
	.A1(n675));
   SEN_EO2_S_0P5 U2585 (.X(pprow1[5]), 
	.A2(\bmul/ppgen1/n6 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U2586 (.X(\bmul/ppgen1/n6 ), 
	.B2(n836), 
	.B1(n854), 
	.A2(n839), 
	.A1(n852));
   SEN_EO2_S_0P5 U2587 (.X(pprow1[6]), 
	.A2(\bmul/ppgen1/n5 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U2588 (.X(\bmul/ppgen1/n5 ), 
	.B2(n836), 
	.B1(n856), 
	.A2(n839), 
	.A1(n854));
   SEN_EO2_S_0P5 U2589 (.X(pprow1[0]), 
	.A2(\bmul/ppgen1/n35 ), 
	.A1(net84586));
   SEN_ND2_G_1 U2590 (.X(\bmul/ppgen1/n35 ), 
	.A2(n837), 
	.A1(n829));
   SEN_EO2_S_0P5 U2591 (.X(pprow1[4]), 
	.A2(\bmul/ppgen1/n7 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U2592 (.X(\bmul/ppgen1/n7 ), 
	.B2(n836), 
	.B1(n852), 
	.A2(n839), 
	.A1(n850));
   SEN_EO2_S_0P5 U2593 (.X(pprow0[0]), 
	.A2(\bmul/ppgen0/n35 ), 
	.A1(n827));
   SEN_ND2_G_1 U2594 (.X(\bmul/ppgen0/n35 ), 
	.A2(n858), 
	.A1(n829));
   SEN_EO2_S_0P5 U2595 (.X(pprow0[2]), 
	.A2(\bmul/ppgen0/n13 ), 
	.A1(n828));
   SEN_AOI22_1 U2596 (.X(\bmul/ppgen0/n13 ), 
	.B2(n807), 
	.B1(n848), 
	.A2(n833), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2597 (.X(pprow0[3]), 
	.A2(\bmul/ppgen0/n9 ), 
	.A1(n828));
   SEN_AOI22_1 U2598 (.X(\bmul/ppgen0/n9 ), 
	.B2(n807), 
	.B1(n850), 
	.A2(n833), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2599 (.X(pprow0[4]), 
	.A2(\bmul/ppgen0/n8 ), 
	.A1(n828));
   SEN_AOI22_1 U2600 (.X(\bmul/ppgen0/n8 ), 
	.B2(n858), 
	.B1(n852), 
	.A2(n833), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2601 (.X(pprow0[5]), 
	.A2(\bmul/ppgen0/n7 ), 
	.A1(n828));
   SEN_AOI22_1 U2602 (.X(\bmul/ppgen0/n7 ), 
	.B2(n807), 
	.B1(n854), 
	.A2(n833), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2603 (.X(pprow3[0]), 
	.A2(n1893), 
	.A1(net84600));
   SEN_ND2_G_1 U2604 (.X(n1893), 
	.A2(n845), 
	.A1(n829));
   SEN_EO2_S_0P5 U2605 (.X(pprow2[0]), 
	.A2(n1869), 
	.A1(n825));
   SEN_ND2_G_1 U2606 (.X(n1869), 
	.A2(n841), 
	.A1(n830));
   SEN_EO2_S_0P5 U2607 (.X(pprow2[1]), 
	.A2(n1858), 
	.A1(n825));
   SEN_AOI22_1 U2608 (.X(n1858), 
	.B2(n840), 
	.B1(n846), 
	.A2(n842), 
	.A1(n830));
   SEN_EO2_S_0P5 U2609 (.X(pprow2[4]), 
	.A2(n1849), 
	.A1(n826));
   SEN_AOI22_1 U2610 (.X(n1849), 
	.B2(n841), 
	.B1(n852), 
	.A2(n843), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2611 (.X(pprow2[5]), 
	.A2(n1848), 
	.A1(n826));
   SEN_AOI22_1 U2612 (.X(n1848), 
	.B2(n841), 
	.B1(n854), 
	.A2(n843), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2613 (.X(pprow2[6]), 
	.A2(n1847), 
	.A1(n826));
   SEN_AOI22_1 U2614 (.X(n1847), 
	.B2(n841), 
	.B1(n856), 
	.A2(n843), 
	.A1(n854));
   SEN_EO2_S_0P5 U2615 (.X(pprow3[2]), 
	.A2(n1877), 
	.A1(net84600));
   SEN_AOI22_T_0P5 U2616 (.X(n1877), 
	.B2(n845), 
	.B1(n848), 
	.A2(n823), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2617 (.X(pprow3[3]), 
	.A2(n1876), 
	.A1(n202));
   SEN_AOI22_T_0P5 U2618 (.X(n1876), 
	.B2(n845), 
	.B1(n850), 
	.A2(n823), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2619 (.X(pprow3[6]), 
	.A2(n1873), 
	.A1(n202));
   SEN_AOI22_1 U2620 (.X(n1873), 
	.B2(n845), 
	.B1(n856), 
	.A2(n823), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2621 (.X(pprow0[6]), 
	.A2(\bmul/ppgen0/n6 ), 
	.A1(n827));
   SEN_AOI22_1 U2622 (.X(\bmul/ppgen0/n6 ), 
	.B2(n807), 
	.B1(n856), 
	.A2(n833), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2623 (.X(Z[14]), 
	.A2(n678), 
	.A1(n677));
   SEN_AO21B_1 U2624 (.X(n678), 
	.B(n1119), 
	.A2(n1263), 
	.A1(n1074));
   SEN_EO2_S_0P5 U2625 (.X(pprow3[4]), 
	.A2(n1875), 
	.A1(n202));
   SEN_AOI22_T_0P5 U2626 (.X(n1875), 
	.B2(n845), 
	.B1(n852), 
	.A2(n822), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2627 (.X(pprow3[1]), 
	.A2(n1882), 
	.A1(net84600));
   SEN_AOI22_T_0P5 U2628 (.X(n1882), 
	.B2(n844), 
	.B1(n846), 
	.A2(n822), 
	.A1(n830));
   SEN_EO2_S_0P5 U2629 (.X(pprow3[5]), 
	.A2(n1874), 
	.A1(n202));
   SEN_AOI22_T_0P5 U2630 (.X(n1874), 
	.B2(n845), 
	.B1(n854), 
	.A2(n822), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2631 (.X(pprow1[1]), 
	.A2(\bmul/ppgen1/n24 ), 
	.A1(net84586));
   SEN_AOI22_T_0P5 U2632 (.X(\bmul/ppgen1/n24 ), 
	.B2(n835), 
	.B1(n846), 
	.A2(n838), 
	.A1(n829));
   SEN_EO2_S_0P5 U2633 (.X(pprow1[2]), 
	.A2(\bmul/ppgen1/n13 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U2634 (.X(\bmul/ppgen1/n13 ), 
	.B2(n836), 
	.B1(n848), 
	.A2(n839), 
	.A1(n846));
   SEN_EO2_S_0P5 U2635 (.X(pprow1[3]), 
	.A2(\bmul/ppgen1/n8 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U2636 (.X(\bmul/ppgen1/n8 ), 
	.B2(n836), 
	.B1(n850), 
	.A2(n839), 
	.A1(n848));
   SEN_EO2_S_0P5 U2637 (.X(pprow0[1]), 
	.A2(\bmul/ppgen0/n24 ), 
	.A1(n827));
   SEN_AOI22_1 U2638 (.X(\bmul/ppgen0/n24 ), 
	.B2(n807), 
	.B1(n846), 
	.A2(n832), 
	.A1(n830));
   SEN_EO2_S_0P5 U2639 (.X(pprow2[2]), 
	.A2(n1851), 
	.A1(n826));
   SEN_AOI22_1 U2640 (.X(n1851), 
	.B2(n841), 
	.B1(n848), 
	.A2(n843), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2641 (.X(pprow2[3]), 
	.A2(n1850), 
	.A1(n826));
   SEN_AOI22_1 U2642 (.X(n1850), 
	.B2(n841), 
	.B1(n850), 
	.A2(n843), 
	.A1(B[2]));
   SEN_AO21_1 U2643 (.X(n1326), 
	.B(n679), 
	.A2(n1325), 
	.A1(n1444));
   SEN_AN2_S_0P5 U2644 (.X(n679), 
	.A2(n1452), 
	.A1(n1450));
   SEN_INV_S_1 U2645 (.X(net82770), 
	.A(net82772));
   SEN_INV_S_1 U2646 (.X(n1536), 
	.A(n1539));
   SEN_INV_S_0P5 U2647 (.X(n905), 
	.A(n923));
   SEN_INV_S_1 U2648 (.X(n832), 
	.A(n687));
   SEN_INV_S_1 U2649 (.X(n833), 
	.A(n687));
   SEN_INV_S_1 U2650 (.X(net84586), 
	.A(net84592));
   SEN_INV_S_1 U2651 (.X(net84588), 
	.A(net84592));
   SEN_INV_S_1 U2652 (.X(n827), 
	.A(n808));
   SEN_INV_S_1 U2653 (.X(n828), 
	.A(n808));
   SEN_INV_S_1 U2654 (.X(net84600), 
	.A(net90815));
   SEN_INV_S_1 U2655 (.X(n825), 
	.A(n809));
   SEN_INV_S_1 U2656 (.X(n826), 
	.A(\bmul/neg2 ));
   SEN_INV_S_1 U2657 (.X(n830), 
	.A(n831));
   SEN_INV_S_1 U2658 (.X(n858), 
	.A(n859));
   SEN_INV_S_1 U2659 (.X(n834), 
	.A(n687));
   SEN_INV_S_0P5 U2660 (.X(n1130), 
	.A(n1183));
   SEN_EN3_1 U2661 (.X(n1707), 
	.A3(n1690), 
	.A2(n1686), 
	.A1(n1689));
   SEN_INV_S_1 U2662 (.X(net83828), 
	.A(net83735));
   SEN_INV_S_1 U2663 (.X(net2269), 
	.A(net84634));
   SEN_ND2B_1 U2664 (.X(n687), 
	.B(n688), 
	.A(n858));
   SEN_EO2_S_0P5 U2665 (.X(n688), 
	.A2(n808), 
	.A1(n858));
   SEN_EO2_2 U2666 (.X(net82514), 
	.A2(n694), 
	.A1(n693));
   SEN_EO2_S_0P5 U2667 (.X(n981), 
	.A2(net84246), 
	.A1(net84067));
   SEN_EO2_S_0P5 U2668 (.X(pprow6[9]), 
	.A2(n1936), 
	.A1(n1841));
   SEN_AOI22_1 U2669 (.X(n1936), 
	.B2(n786), 
	.B1(\bmul/one6 ), 
	.A2(n784), 
	.A1(\bmul/two6 ));
   SEN_EO2_S_0P5 U2670 (.X(pprow11[0]), 
	.A2(n2013), 
	.A1(net2269));
   SEN_ND2_G_1 U2671 (.X(n2013), 
	.A2(\bmul/one11 ), 
	.A1(n829));
   SEN_EO2_S_0P5 U2672 (.X(pprow11[1]), 
	.A2(n2012), 
	.A1(net2269));
   SEN_AOI22_1 U2673 (.X(n2012), 
	.B2(\bmul/one11 ), 
	.B1(n846), 
	.A2(\bmul/two11 ), 
	.A1(n830));
   SEN_EO2_S_0P5 U2674 (.X(pprow11[2]), 
	.A2(n2011), 
	.A1(net2269));
   SEN_AOI22_1 U2675 (.X(n2011), 
	.B2(\bmul/one11 ), 
	.B1(n848), 
	.A2(\bmul/two11 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2676 (.X(pprow11[3]), 
	.A2(n2010), 
	.A1(net2269));
   SEN_AOI22_1 U2677 (.X(n2010), 
	.B2(\bmul/one11 ), 
	.B1(n850), 
	.A2(\bmul/two11 ), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2678 (.X(pprow11[4]), 
	.A2(n2009), 
	.A1(net2269));
   SEN_AOI22_1 U2679 (.X(n2009), 
	.B2(\bmul/one11 ), 
	.B1(n852), 
	.A2(\bmul/two11 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2680 (.X(pprow11[5]), 
	.A2(n2008), 
	.A1(net2269));
   SEN_AOI22_1 U2681 (.X(n2008), 
	.B2(\bmul/one11 ), 
	.B1(n854), 
	.A2(\bmul/two11 ), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2682 (.X(pprow11[6]), 
	.A2(n2007), 
	.A1(net2269));
   SEN_AOI22_1 U2683 (.X(n2007), 
	.B2(\bmul/one11 ), 
	.B1(n856), 
	.A2(\bmul/two11 ), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2684 (.X(pprow11[7]), 
	.A2(n2006), 
	.A1(net2269));
   SEN_AOI22_1 U2685 (.X(n2006), 
	.B2(\bmul/one11 ), 
	.B1(B[7]), 
	.A2(\bmul/two11 ), 
	.A1(B[6]));
   SEN_NR2_1 U2686 (.X(\bmul/two4 ), 
	.A2(n2025), 
	.A1(n772));
   SEN_EO2_S_0P5 U2687 (.X(n697), 
	.A2(net82141), 
	.A1(net85926));
   SEN_NR2_1 U2688 (.X(n824), 
	.A2(n2025), 
	.A1(n772));
   SEN_EO2_S_0P5 U2689 (.X(pprow12[1]), 
	.A2(n2018), 
	.A1(n1489));
   SEN_AOI22_1 U2690 (.X(n2018), 
	.B2(\bmul/one12 ), 
	.B1(n846), 
	.A2(\bmul/two12 ), 
	.A1(n830));
   SEN_EO2_S_0P5 U2691 (.X(pprow12[2]), 
	.A2(n2017), 
	.A1(n1489));
   SEN_AOI22_1 U2692 (.X(n2017), 
	.B2(\bmul/one12 ), 
	.B1(n848), 
	.A2(\bmul/two12 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2693 (.X(pprow12[3]), 
	.A2(n2016), 
	.A1(n1489));
   SEN_AOI22_1 U2694 (.X(n2016), 
	.B2(\bmul/one12 ), 
	.B1(n850), 
	.A2(\bmul/two12 ), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2695 (.X(pprow12[4]), 
	.A2(n2015), 
	.A1(n1489));
   SEN_AOI22_1 U2696 (.X(n2015), 
	.B2(\bmul/one12 ), 
	.B1(n852), 
	.A2(\bmul/two12 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2697 (.X(pprow12[5]), 
	.A2(n2014), 
	.A1(n1489));
   SEN_AOI22_1 U2698 (.X(n2014), 
	.B2(\bmul/one12 ), 
	.B1(n854), 
	.A2(\bmul/two12 ), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2699 (.X(pprow5[1]), 
	.A2(n1924), 
	.A1(n819));
   SEN_AOI22_1 U2700 (.X(n1924), 
	.B2(\bmul/one5 ), 
	.B1(n846), 
	.A2(\bmul/two5 ), 
	.A1(n830));
   SEN_EO2_S_0P5 U2701 (.X(pprow5[2]), 
	.A2(n1923), 
	.A1(n819));
   SEN_AOI22_1 U2702 (.X(n1923), 
	.B2(\bmul/one5 ), 
	.B1(n848), 
	.A2(\bmul/two5 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2703 (.X(pprow5[3]), 
	.A2(n1922), 
	.A1(n819));
   SEN_AOI22_1 U2704 (.X(n1922), 
	.B2(\bmul/one5 ), 
	.B1(n850), 
	.A2(\bmul/two5 ), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2705 (.X(pprow5[4]), 
	.A2(n1921), 
	.A1(n819));
   SEN_AOI22_1 U2706 (.X(n1921), 
	.B2(n613), 
	.B1(n852), 
	.A2(\bmul/two5 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2707 (.X(pprow5[5]), 
	.A2(n1920), 
	.A1(n819));
   SEN_AOI22_1 U2708 (.X(n1920), 
	.B2(\bmul/one5 ), 
	.B1(n854), 
	.A2(\bmul/two5 ), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2709 (.X(pprow5[6]), 
	.A2(n1919), 
	.A1(n819));
   SEN_AOI22_1 U2710 (.X(n1919), 
	.B2(n613), 
	.B1(n856), 
	.A2(\bmul/two5 ), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2711 (.X(pprow5[7]), 
	.A2(n1918), 
	.A1(n819));
   SEN_AOI22_1 U2712 (.X(n1918), 
	.B2(n613), 
	.B1(B[7]), 
	.A2(\bmul/two5 ), 
	.A1(B[6]));
   SEN_EO2_S_0P5 U2713 (.X(pprow5[11]), 
	.A2(n1933), 
	.A1(n819));
   SEN_AOI22_1 U2714 (.X(n1933), 
	.B2(n613), 
	.B1(n789), 
	.A2(\bmul/two5 ), 
	.A1(n788));
   SEN_EO2_S_0P5 U2715 (.X(pprow5[12]), 
	.A2(n1932), 
	.A1(n819));
   SEN_AOI22_1 U2716 (.X(n1932), 
	.B2(\bmul/one5 ), 
	.B1(n790), 
	.A2(\bmul/two5 ), 
	.A1(n789));
   SEN_EO2_S_0P5 U2717 (.X(pprow5[13]), 
	.A2(n1931), 
	.A1(n819));
   SEN_AOI22_1 U2718 (.X(n1931), 
	.B2(\bmul/one5 ), 
	.B1(n791), 
	.A2(\bmul/two5 ), 
	.A1(n790));
   SEN_EO2_S_0P5 U2719 (.X(pprow5[14]), 
	.A2(n1930), 
	.A1(n819));
   SEN_AOI22_1 U2720 (.X(n1930), 
	.B2(\bmul/one5 ), 
	.B1(n792), 
	.A2(\bmul/two5 ), 
	.A1(n791));
   SEN_EO2_S_0P5 U2721 (.X(pprow5[15]), 
	.A2(n1929), 
	.A1(n608));
   SEN_AOI22_1 U2722 (.X(n1929), 
	.B2(n613), 
	.B1(n793), 
	.A2(n607), 
	.A1(n792));
   SEN_EO2_S_0P5 U2723 (.X(pprow5[16]), 
	.A2(n1928), 
	.A1(n608));
   SEN_AOI22_1 U2724 (.X(n1928), 
	.B2(n613), 
	.B1(n794), 
	.A2(n607), 
	.A1(n793));
   SEN_EO2_S_0P5 U2725 (.X(pprow5[17]), 
	.A2(n1927), 
	.A1(n608));
   SEN_AOI22_1 U2726 (.X(n1927), 
	.B2(n613), 
	.B1(n795), 
	.A2(n607), 
	.A1(n794));
   SEN_EO2_S_0P5 U2727 (.X(pprow5[18]), 
	.A2(n1926), 
	.A1(n608));
   SEN_AOI22_1 U2728 (.X(n1926), 
	.B2(n613), 
	.B1(n796), 
	.A2(n607), 
	.A1(n795));
   SEN_EO2_S_0P5 U2729 (.X(pprow5[19]), 
	.A2(n1925), 
	.A1(n608));
   SEN_AOI22_1 U2730 (.X(n1925), 
	.B2(n613), 
	.B1(n797), 
	.A2(n607), 
	.A1(n796));
   SEN_EO2_S_0P5 U2731 (.X(pprow14[0]), 
	.A2(\bmul/ppgen14/n35 ), 
	.A1(n1836));
   SEN_ND2_G_1 U2732 (.X(\bmul/ppgen14/n35 ), 
	.A2(\bmul/one14 ), 
	.A1(n829));
   SEN_EO2_S_0P5 U2733 (.X(pprow6[1]), 
	.A2(n1944), 
	.A1(n1015));
   SEN_AOI22_1 U2734 (.X(n1944), 
	.B2(\bmul/one6 ), 
	.B1(n846), 
	.A2(n606), 
	.A1(n830));
   SEN_EO2_S_0P5 U2735 (.X(pprow6[2]), 
	.A2(n1943), 
	.A1(n1841));
   SEN_AOI22_1 U2736 (.X(n1943), 
	.B2(\bmul/one6 ), 
	.B1(n848), 
	.A2(\bmul/two6 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2737 (.X(pprow6[3]), 
	.A2(n1942), 
	.A1(n1015));
   SEN_AOI22_1 U2738 (.X(n1942), 
	.B2(\bmul/one6 ), 
	.B1(n850), 
	.A2(n606), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2739 (.X(pprow6[4]), 
	.A2(n1941), 
	.A1(n1841));
   SEN_AOI22_1 U2740 (.X(n1941), 
	.B2(\bmul/one6 ), 
	.B1(n852), 
	.A2(\bmul/two6 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2741 (.X(pprow6[5]), 
	.A2(n1940), 
	.A1(n1841));
   SEN_AOI22_1 U2742 (.X(n1940), 
	.B2(\bmul/one6 ), 
	.B1(n854), 
	.A2(\bmul/two6 ), 
	.A1(n852));
   SEN_EO2_S_0P5 U2743 (.X(pprow6[6]), 
	.A2(n1939), 
	.A1(n1841));
   SEN_AOI22_1 U2744 (.X(n1939), 
	.B2(\bmul/one6 ), 
	.B1(n856), 
	.A2(\bmul/two6 ), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2745 (.X(pprow6[7]), 
	.A2(n1938), 
	.A1(n1841));
   SEN_AOI22_1 U2746 (.X(n1938), 
	.B2(\bmul/one6 ), 
	.B1(B[7]), 
	.A2(\bmul/two6 ), 
	.A1(B[6]));
   SEN_EO2_S_0P5 U2747 (.X(pprow6[11]), 
	.A2(n1951), 
	.A1(n1841));
   SEN_AOI22_1 U2748 (.X(n1951), 
	.B2(n612), 
	.B1(n789), 
	.A2(\bmul/two6 ), 
	.A1(n788));
   SEN_EO2_S_0P5 U2749 (.X(pprow6[12]), 
	.A2(n1950), 
	.A1(n1841));
   SEN_AOI22_1 U2750 (.X(n1950), 
	.B2(\bmul/one6 ), 
	.B1(n790), 
	.A2(\bmul/two6 ), 
	.A1(n789));
   SEN_EO2_S_0P5 U2751 (.X(pprow6[13]), 
	.A2(n1949), 
	.A1(n1841));
   SEN_AOI22_1 U2752 (.X(n1949), 
	.B2(\bmul/one6 ), 
	.B1(n791), 
	.A2(\bmul/two6 ), 
	.A1(n790));
   SEN_EO2_S_0P5 U2753 (.X(pprow6[14]), 
	.A2(n1948), 
	.A1(n1841));
   SEN_AOI22_1 U2754 (.X(n1948), 
	.B2(n612), 
	.B1(n792), 
	.A2(\bmul/two6 ), 
	.A1(n791));
   SEN_EO2_S_0P5 U2755 (.X(pprow6[15]), 
	.A2(n1947), 
	.A1(n1841));
   SEN_AOI22_1 U2756 (.X(n1947), 
	.B2(n612), 
	.B1(n793), 
	.A2(\bmul/two6 ), 
	.A1(n792));
   SEN_EO2_S_0P5 U2757 (.X(pprow6[16]), 
	.A2(n1946), 
	.A1(n1841));
   SEN_AOI22_1 U2758 (.X(n1946), 
	.B2(n612), 
	.B1(n794), 
	.A2(\bmul/two6 ), 
	.A1(n793));
   SEN_EO2_S_0P5 U2759 (.X(pprow6[17]), 
	.A2(n1945), 
	.A1(n1841));
   SEN_AOI22_1 U2760 (.X(n1945), 
	.B2(n612), 
	.B1(n795), 
	.A2(\bmul/two6 ), 
	.A1(n794));
   SEN_EO2_S_0P5 U2761 (.X(pprow13[1]), 
	.A2(n2022), 
	.A1(n1837));
   SEN_AOI22_1 U2762 (.X(n2022), 
	.B2(\bmul/one13 ), 
	.B1(n846), 
	.A2(\bmul/two13 ), 
	.A1(n830));
   SEN_EO2_S_0P5 U2763 (.X(pprow13[2]), 
	.A2(n2021), 
	.A1(n1837));
   SEN_AOI22_1 U2764 (.X(n2021), 
	.B2(\bmul/one13 ), 
	.B1(n848), 
	.A2(\bmul/two13 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2765 (.X(pprow13[3]), 
	.A2(n2020), 
	.A1(n1837));
   SEN_AOI22_1 U2766 (.X(n2020), 
	.B2(\bmul/one13 ), 
	.B1(n850), 
	.A2(\bmul/two13 ), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2767 (.X(pprow13[0]), 
	.A2(n2023), 
	.A1(n1837));
   SEN_ND2_G_1 U2768 (.X(n2023), 
	.A2(\bmul/one13 ), 
	.A1(n829));
   SEN_EO2_S_0P5 U2769 (.X(pprow8[1]), 
	.A2(n1978), 
	.A1(n817));
   SEN_AOI22_1 U2770 (.X(n1978), 
	.B2(\bmul/one8 ), 
	.B1(n846), 
	.A2(\bmul/two8 ), 
	.A1(n830));
   SEN_EO2_S_0P5 U2771 (.X(pprow8[2]), 
	.A2(n1977), 
	.A1(n817));
   SEN_AOI22_1 U2772 (.X(n1977), 
	.B2(\bmul/one8 ), 
	.B1(n848), 
	.A2(\bmul/two8 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2773 (.X(pprow8[3]), 
	.A2(n1976), 
	.A1(n817));
   SEN_AOI22_1 U2774 (.X(n1976), 
	.B2(\bmul/one8 ), 
	.B1(n850), 
	.A2(\bmul/two8 ), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2775 (.X(pprow8[4]), 
	.A2(n1975), 
	.A1(n817));
   SEN_AOI22_1 U2776 (.X(n1975), 
	.B2(\bmul/one8 ), 
	.B1(n852), 
	.A2(\bmul/two8 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2777 (.X(pprow8[5]), 
	.A2(n1974), 
	.A1(n817));
   SEN_AOI22_1 U2778 (.X(n1974), 
	.B2(\bmul/one8 ), 
	.B1(n854), 
	.A2(\bmul/two8 ), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2779 (.X(pprow8[6]), 
	.A2(n1973), 
	.A1(n817));
   SEN_AOI22_1 U2780 (.X(n1973), 
	.B2(\bmul/one8 ), 
	.B1(n856), 
	.A2(\bmul/two8 ), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2781 (.X(pprow8[7]), 
	.A2(n1972), 
	.A1(n817));
   SEN_AOI22_1 U2782 (.X(n1972), 
	.B2(\bmul/one8 ), 
	.B1(B[7]), 
	.A2(\bmul/two8 ), 
	.A1(B[6]));
   SEN_EO2_S_0P5 U2783 (.X(pprow8[11]), 
	.A2(n1981), 
	.A1(n817));
   SEN_AOI22_1 U2784 (.X(n1981), 
	.B2(\bmul/one8 ), 
	.B1(n789), 
	.A2(\bmul/two8 ), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2785 (.X(pprow8[12]), 
	.A2(n1980), 
	.A1(n817));
   SEN_AOI22_1 U2786 (.X(n1980), 
	.B2(\bmul/one8 ), 
	.B1(n790), 
	.A2(\bmul/two8 ), 
	.A1(n610));
   SEN_EO2_S_0P5 U2787 (.X(pprow8[13]), 
	.A2(n1979), 
	.A1(n817));
   SEN_AOI22_1 U2788 (.X(n1979), 
	.B2(\bmul/one8 ), 
	.B1(n791), 
	.A2(\bmul/two8 ), 
	.A1(n605));
   SEN_EO2_S_0P5 U2789 (.X(pprow4[7]), 
	.A2(n1896), 
	.A1(n820));
   SEN_AOI22_1 U2790 (.X(n1896), 
	.B2(n773), 
	.B1(B[7]), 
	.A2(n824), 
	.A1(B[6]));
   SEN_EO2_S_0P5 U2791 (.X(pprow4[8]), 
	.A2(n1895), 
	.A1(n820));
   SEN_AOI22_0P5 U2792 (.X(n1895), 
	.B2(n784), 
	.B1(n773), 
	.A2(\bmul/two4 ), 
	.A1(B[7]));
   SEN_EO2_S_0P5 U2793 (.X(pprow4[10]), 
	.A2(n1914), 
	.A1(n820));
   SEN_AOI22_0P5 U2794 (.X(n1914), 
	.B2(n824), 
	.B1(n786), 
	.A2(n773), 
	.A1(n788));
   SEN_EO2_S_0P5 U2795 (.X(pprow4[11]), 
	.A2(n1913), 
	.A1(n820));
   SEN_AOI22_1 U2796 (.X(n1913), 
	.B2(n772), 
	.B1(n789), 
	.A2(\bmul/two4 ), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2797 (.X(pprow4[12]), 
	.A2(n1912), 
	.A1(n820));
   SEN_AOI22_1 U2798 (.X(n1912), 
	.B2(n772), 
	.B1(n790), 
	.A2(n824), 
	.A1(n610));
   SEN_EO2_S_0P5 U2799 (.X(pprow4[13]), 
	.A2(n1911), 
	.A1(n820));
   SEN_AOI22_1 U2800 (.X(n1911), 
	.B2(n772), 
	.B1(n791), 
	.A2(\bmul/two4 ), 
	.A1(n790));
   SEN_EO2_S_0P5 U2801 (.X(pprow4[14]), 
	.A2(n1910), 
	.A1(n820));
   SEN_AOI22_1 U2802 (.X(n1910), 
	.B2(n772), 
	.B1(n792), 
	.A2(n824), 
	.A1(n791));
   SEN_EO2_S_0P5 U2803 (.X(pprow4[15]), 
	.A2(n1909), 
	.A1(n820));
   SEN_AOI22_1 U2804 (.X(n1909), 
	.B2(n772), 
	.B1(n793), 
	.A2(\bmul/two4 ), 
	.A1(n792));
   SEN_EO2_S_0P5 U2805 (.X(pprow4[16]), 
	.A2(n1908), 
	.A1(n614));
   SEN_AOI22_1 U2806 (.X(n1908), 
	.B2(n772), 
	.B1(n794), 
	.A2(n824), 
	.A1(n793));
   SEN_EO2_S_0P5 U2807 (.X(pprow4[17]), 
	.A2(n1907), 
	.A1(n614));
   SEN_AOI22_1 U2808 (.X(n1907), 
	.B2(n772), 
	.B1(n795), 
	.A2(\bmul/two4 ), 
	.A1(n794));
   SEN_EO2_S_0P5 U2809 (.X(pprow4[18]), 
	.A2(n1906), 
	.A1(n614));
   SEN_AOI22_1 U2810 (.X(n1906), 
	.B2(n772), 
	.B1(n796), 
	.A2(n824), 
	.A1(n795));
   SEN_EO2_S_0P5 U2811 (.X(pprow4[19]), 
	.A2(n1905), 
	.A1(n614));
   SEN_AOI22_1 U2812 (.X(n1905), 
	.B2(n772), 
	.B1(n797), 
	.A2(\bmul/two4 ), 
	.A1(n796));
   SEN_EO2_S_0P5 U2813 (.X(pprow4[20]), 
	.A2(n1903), 
	.A1(n614));
   SEN_AOI22_1 U2814 (.X(n1903), 
	.B2(n772), 
	.B1(n798), 
	.A2(\bmul/two4 ), 
	.A1(n797));
   SEN_EO2_S_0P5 U2815 (.X(pprow4[21]), 
	.A2(n1902), 
	.A1(n614));
   SEN_AOI22_1 U2816 (.X(n1902), 
	.B2(n772), 
	.B1(n799), 
	.A2(n824), 
	.A1(n798));
   SEN_EO2_S_0P5 U2817 (.X(pprow5[0]), 
	.A2(n1935), 
	.A1(n819));
   SEN_ND2_G_1 U2818 (.X(n1935), 
	.A2(n613), 
	.A1(n829));
   SEN_EO2_S_0P5 U2819 (.X(pprow5[8]), 
	.A2(n1917), 
	.A1(n819));
   SEN_AOI22_1 U2820 (.X(n1917), 
	.B2(n784), 
	.B1(\bmul/one5 ), 
	.A2(\bmul/two5 ), 
	.A1(B[7]));
   SEN_EO2_S_0P5 U2821 (.X(pprow5[9]), 
	.A2(n1916), 
	.A1(n819));
   SEN_AOI22_1 U2822 (.X(n1916), 
	.B2(n786), 
	.B1(\bmul/one5 ), 
	.A2(n784), 
	.A1(\bmul/two5 ));
   SEN_EO2_S_0P5 U2823 (.X(pprow5[10]), 
	.A2(n1934), 
	.A1(n608));
   SEN_AOI22_1 U2824 (.X(n1934), 
	.B2(\bmul/two5 ), 
	.B1(B[9]), 
	.A2(n613), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2825 (.X(pprow10[0]), 
	.A2(n2005), 
	.A1(net2268));
   SEN_ND2_G_1 U2826 (.X(n2005), 
	.A2(\bmul/one10 ), 
	.A1(n829));
   SEN_EO2_S_0P5 U2827 (.X(pprow10[1]), 
	.A2(n2004), 
	.A1(net2268));
   SEN_AOI22_1 U2828 (.X(n2004), 
	.B2(\bmul/one10 ), 
	.B1(B[1]), 
	.A2(\bmul/two10 ), 
	.A1(n830));
   SEN_EO2_S_0P5 U2829 (.X(pprow10[2]), 
	.A2(n2003), 
	.A1(net2268));
   SEN_AOI22_1 U2830 (.X(n2003), 
	.B2(\bmul/one10 ), 
	.B1(n848), 
	.A2(\bmul/two10 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2831 (.X(pprow10[3]), 
	.A2(n2002), 
	.A1(net2268));
   SEN_AOI22_1 U2832 (.X(n2002), 
	.B2(\bmul/one10 ), 
	.B1(n850), 
	.A2(\bmul/two10 ), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2833 (.X(pprow10[4]), 
	.A2(n2001), 
	.A1(net2268));
   SEN_AOI22_1 U2834 (.X(n2001), 
	.B2(\bmul/one10 ), 
	.B1(n852), 
	.A2(\bmul/two10 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2835 (.X(pprow10[5]), 
	.A2(n2000), 
	.A1(net2268));
   SEN_AOI22_1 U2836 (.X(n2000), 
	.B2(\bmul/one10 ), 
	.B1(n854), 
	.A2(\bmul/two10 ), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2837 (.X(pprow10[6]), 
	.A2(n1999), 
	.A1(net2268));
   SEN_AOI22_1 U2838 (.X(n1999), 
	.B2(\bmul/one10 ), 
	.B1(n856), 
	.A2(\bmul/two10 ), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2839 (.X(pprow10[7]), 
	.A2(n1998), 
	.A1(net2268));
   SEN_AOI22_1 U2840 (.X(n1998), 
	.B2(\bmul/one10 ), 
	.B1(B[7]), 
	.A2(\bmul/two10 ), 
	.A1(B[6]));
   SEN_EO2_S_0P5 U2841 (.X(pprow10[8]), 
	.A2(n1997), 
	.A1(net2268));
   SEN_AOI22_1 U2842 (.X(n1997), 
	.B2(n784), 
	.B1(\bmul/one10 ), 
	.A2(\bmul/two10 ), 
	.A1(n615));
   SEN_EO2_S_0P5 U2843 (.X(pprow10[9]), 
	.A2(n1996), 
	.A1(net2268));
   SEN_AOI22_1 U2844 (.X(n1996), 
	.B2(n786), 
	.B1(\bmul/one10 ), 
	.A2(B[8]), 
	.A1(\bmul/two10 ));
   SEN_EO2_S_0P5 U2845 (.X(pprow6[0]), 
	.A2(n1953), 
	.A1(n1841));
   SEN_ND2_G_1 U2846 (.X(n1953), 
	.A2(n612), 
	.A1(n829));
   SEN_EO2_S_0P5 U2847 (.X(pprow6[8]), 
	.A2(n1937), 
	.A1(n1841));
   SEN_AOI22_1 U2848 (.X(n1937), 
	.B2(n784), 
	.B1(n612), 
	.A2(n606), 
	.A1(n615));
   SEN_EO2_S_0P5 U2849 (.X(pprow6[10]), 
	.A2(n1952), 
	.A1(n1015));
   SEN_AOI22_1 U2850 (.X(n1952), 
	.B2(\bmul/two6 ), 
	.B1(B[9]), 
	.A2(n612), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2851 (.X(pprow7[1]), 
	.A2(n1962), 
	.A1(n818));
   SEN_AOI22_1 U2852 (.X(n1962), 
	.B2(\bmul/one7 ), 
	.B1(n846), 
	.A2(\bmul/two7 ), 
	.A1(n830));
   SEN_EO2_S_0P5 U2853 (.X(pprow7[2]), 
	.A2(n1961), 
	.A1(n818));
   SEN_AOI22_1 U2854 (.X(n1961), 
	.B2(\bmul/one7 ), 
	.B1(n848), 
	.A2(\bmul/two7 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2855 (.X(pprow7[3]), 
	.A2(n1960), 
	.A1(n818));
   SEN_AOI22_1 U2856 (.X(n1960), 
	.B2(\bmul/one7 ), 
	.B1(n850), 
	.A2(\bmul/two7 ), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2857 (.X(pprow7[4]), 
	.A2(n1959), 
	.A1(n818));
   SEN_AOI22_1 U2858 (.X(n1959), 
	.B2(\bmul/one7 ), 
	.B1(n852), 
	.A2(\bmul/two7 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2859 (.X(pprow7[5]), 
	.A2(n1958), 
	.A1(n1840));
   SEN_AOI22_1 U2860 (.X(n1958), 
	.B2(\bmul/one7 ), 
	.B1(n854), 
	.A2(\bmul/two7 ), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2861 (.X(pprow7[6]), 
	.A2(n1957), 
	.A1(n818));
   SEN_AOI22_1 U2862 (.X(n1957), 
	.B2(\bmul/one7 ), 
	.B1(n856), 
	.A2(\bmul/two7 ), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2863 (.X(pprow7[8]), 
	.A2(n1955), 
	.A1(n818));
   SEN_AOI22_1 U2864 (.X(n1955), 
	.B2(n784), 
	.B1(n611), 
	.A2(\bmul/two7 ), 
	.A1(n615));
   SEN_EO2_S_0P5 U2865 (.X(pprow7[9]), 
	.A2(n1954), 
	.A1(n818));
   SEN_AOI22_1 U2866 (.X(n1954), 
	.B2(n786), 
	.B1(n611), 
	.A2(B[8]), 
	.A1(\bmul/two7 ));
   SEN_EO2_S_0P5 U2867 (.X(pprow7[10]), 
	.A2(n1968), 
	.A1(n818));
   SEN_AOI22_1 U2868 (.X(n1968), 
	.B2(\bmul/two7 ), 
	.B1(B[9]), 
	.A2(n611), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2869 (.X(pprow7[11]), 
	.A2(n1967), 
	.A1(n818));
   SEN_AOI22_1 U2870 (.X(n1967), 
	.B2(n611), 
	.B1(n789), 
	.A2(\bmul/two7 ), 
	.A1(n788));
   SEN_EO2_S_0P5 U2871 (.X(pprow7[12]), 
	.A2(n1966), 
	.A1(n818));
   SEN_AOI22_1 U2872 (.X(n1966), 
	.B2(\bmul/one7 ), 
	.B1(n790), 
	.A2(\bmul/two7 ), 
	.A1(n610));
   SEN_EO2_S_0P5 U2873 (.X(pprow7[13]), 
	.A2(n1965), 
	.A1(n818));
   SEN_AOI22_1 U2874 (.X(n1965), 
	.B2(\bmul/one7 ), 
	.B1(n791), 
	.A2(\bmul/two7 ), 
	.A1(n790));
   SEN_EO2_S_0P5 U2875 (.X(pprow7[14]), 
	.A2(n1964), 
	.A1(n818));
   SEN_AOI22_1 U2876 (.X(n1964), 
	.B2(\bmul/one7 ), 
	.B1(n792), 
	.A2(\bmul/two7 ), 
	.A1(n791));
   SEN_EO2_S_0P5 U2877 (.X(pprow7[15]), 
	.A2(n1963), 
	.A1(n818));
   SEN_AOI22_1 U2878 (.X(n1963), 
	.B2(n611), 
	.B1(n793), 
	.A2(\bmul/two7 ), 
	.A1(n792));
   SEN_EO2_S_0P5 U2879 (.X(pprow8[0]), 
	.A2(n1983), 
	.A1(n817));
   SEN_ND2_G_1 U2880 (.X(n1983), 
	.A2(\bmul/one8 ), 
	.A1(n829));
   SEN_EO2_S_0P5 U2881 (.X(pprow8[8]), 
	.A2(n1971), 
	.A1(n817));
   SEN_AOI22_1 U2882 (.X(n1971), 
	.B2(n784), 
	.B1(\bmul/one8 ), 
	.A2(\bmul/two8 ), 
	.A1(n615));
   SEN_EO2_S_0P5 U2883 (.X(pprow8[9]), 
	.A2(n1970), 
	.A1(n817));
   SEN_AOI22_1 U2884 (.X(n1970), 
	.B2(n786), 
	.B1(\bmul/one8 ), 
	.A2(B[8]), 
	.A1(\bmul/two8 ));
   SEN_EO2_S_0P5 U2885 (.X(pprow8[10]), 
	.A2(n1982), 
	.A1(n817));
   SEN_AOI22_1 U2886 (.X(n1982), 
	.B2(\bmul/two8 ), 
	.B1(B[9]), 
	.A2(\bmul/one8 ), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2887 (.X(pprow9[0]), 
	.A2(n1995), 
	.A1(n1838));
   SEN_ND2_G_1 U2888 (.X(n1995), 
	.A2(\bmul/one9 ), 
	.A1(n829));
   SEN_EO2_S_0P5 U2889 (.X(pprow9[1]), 
	.A2(n1992), 
	.A1(n1838));
   SEN_AOI22_1 U2890 (.X(n1992), 
	.B2(\bmul/one9 ), 
	.B1(n846), 
	.A2(\bmul/two9 ), 
	.A1(n830));
   SEN_EO2_S_0P5 U2891 (.X(pprow9[2]), 
	.A2(n1991), 
	.A1(n1838));
   SEN_AOI22_1 U2892 (.X(n1991), 
	.B2(\bmul/one9 ), 
	.B1(n848), 
	.A2(\bmul/two9 ), 
	.A1(B[1]));
   SEN_EO2_S_0P5 U2893 (.X(pprow9[3]), 
	.A2(n1990), 
	.A1(n1838));
   SEN_AOI22_1 U2894 (.X(n1990), 
	.B2(\bmul/one9 ), 
	.B1(n850), 
	.A2(\bmul/two9 ), 
	.A1(B[2]));
   SEN_EO2_S_0P5 U2895 (.X(pprow9[4]), 
	.A2(n1989), 
	.A1(n1838));
   SEN_AOI22_1 U2896 (.X(n1989), 
	.B2(\bmul/one9 ), 
	.B1(n852), 
	.A2(\bmul/two9 ), 
	.A1(B[3]));
   SEN_EO2_S_0P5 U2897 (.X(pprow9[5]), 
	.A2(n1988), 
	.A1(n1838));
   SEN_AOI22_1 U2898 (.X(n1988), 
	.B2(\bmul/one9 ), 
	.B1(n854), 
	.A2(\bmul/two9 ), 
	.A1(B[4]));
   SEN_EO2_S_0P5 U2899 (.X(pprow9[6]), 
	.A2(n1987), 
	.A1(n1838));
   SEN_AOI22_1 U2900 (.X(n1987), 
	.B2(\bmul/one9 ), 
	.B1(n856), 
	.A2(\bmul/two9 ), 
	.A1(B[5]));
   SEN_EO2_S_0P5 U2901 (.X(pprow9[7]), 
	.A2(n1986), 
	.A1(n1838));
   SEN_AOI22_1 U2902 (.X(n1986), 
	.B2(\bmul/one9 ), 
	.B1(n615), 
	.A2(\bmul/two9 ), 
	.A1(B[6]));
   SEN_EO2_S_0P5 U2903 (.X(pprow9[8]), 
	.A2(n1985), 
	.A1(n1838));
   SEN_AOI22_1 U2904 (.X(n1985), 
	.B2(n784), 
	.B1(\bmul/one9 ), 
	.A2(\bmul/two9 ), 
	.A1(n615));
   SEN_EO2_S_0P5 U2905 (.X(pprow9[9]), 
	.A2(n1984), 
	.A1(n1838));
   SEN_AOI22_1 U2906 (.X(n1984), 
	.B2(n786), 
	.B1(\bmul/one9 ), 
	.A2(B[8]), 
	.A1(\bmul/two9 ));
   SEN_EO2_S_0P5 U2907 (.X(pprow9[10]), 
	.A2(n1994), 
	.A1(n1838));
   SEN_AOI22_1 U2908 (.X(n1994), 
	.B2(\bmul/two9 ), 
	.B1(B[9]), 
	.A2(\bmul/one9 ), 
	.A1(n788));
   SEN_EO2_S_0P5 U2909 (.X(pprow9[11]), 
	.A2(n1993), 
	.A1(n1838));
   SEN_AOI22_1 U2910 (.X(n1993), 
	.B2(\bmul/one9 ), 
	.B1(n789), 
	.A2(\bmul/two9 ), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2911 (.X(pprow1[7]), 
	.A2(\bmul/ppgen1/n4 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U2912 (.X(\bmul/ppgen1/n4 ), 
	.B2(n836), 
	.B1(B[7]), 
	.A2(n839), 
	.A1(n856));
   SEN_EO2_S_0P5 U2913 (.X(pprow1[16]), 
	.A2(\bmul/ppgen1/n28 ), 
	.A1(net84586));
   SEN_AOI22_T_0P5 U2914 (.X(\bmul/ppgen1/n28 ), 
	.B2(n835), 
	.B1(n794), 
	.A2(n838), 
	.A1(n793));
   SEN_EO2_S_0P5 U2915 (.X(pprow1[12]), 
	.A2(\bmul/ppgen1/n32 ), 
	.A1(net84586));
   SEN_AOI22_0P5 U2916 (.X(\bmul/ppgen1/n32 ), 
	.B2(n835), 
	.B1(n790), 
	.A2(n838), 
	.A1(n789));
   SEN_EO2_S_0P5 U2917 (.X(pprow1[14]), 
	.A2(\bmul/ppgen1/n30 ), 
	.A1(net84586));
   SEN_AOI22_0P5 U2918 (.X(\bmul/ppgen1/n30 ), 
	.B2(n835), 
	.B1(B[14]), 
	.A2(n838), 
	.A1(n791));
   SEN_EO2_S_0P5 U2919 (.X(pprow1[17]), 
	.A2(\bmul/ppgen1/n27 ), 
	.A1(net84586));
   SEN_AOI22_0P5 U2920 (.X(\bmul/ppgen1/n27 ), 
	.B2(n835), 
	.B1(n795), 
	.A2(n838), 
	.A1(n794));
   SEN_EO2_S_0P5 U2921 (.X(pprow1[18]), 
	.A2(\bmul/ppgen1/n26 ), 
	.A1(net84586));
   SEN_AOI22_0P5 U2922 (.X(\bmul/ppgen1/n26 ), 
	.B2(n835), 
	.B1(n796), 
	.A2(n838), 
	.A1(n795));
   SEN_EO2_S_0P5 U2923 (.X(pprow1[19]), 
	.A2(\bmul/ppgen1/n25 ), 
	.A1(net84586));
   SEN_AOI22_0P5 U2924 (.X(\bmul/ppgen1/n25 ), 
	.B2(n835), 
	.B1(n797), 
	.A2(n838), 
	.A1(n796));
   SEN_EO2_S_0P5 U2925 (.X(pprow1[21]), 
	.A2(\bmul/ppgen1/n22 ), 
	.A1(net84586));
   SEN_AOI22_0P5 U2926 (.X(\bmul/ppgen1/n22 ), 
	.B2(n835), 
	.B1(n799), 
	.A2(n838), 
	.A1(n798));
   SEN_EO2_S_0P5 U2927 (.X(pprow1[22]), 
	.A2(\bmul/ppgen1/n21 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U2928 (.X(\bmul/ppgen1/n21 ), 
	.B2(n835), 
	.B1(n800), 
	.A2(n838), 
	.A1(n799));
   SEN_EO2_S_0P5 U2929 (.X(pprow1[24]), 
	.A2(\bmul/ppgen1/n19 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U2930 (.X(\bmul/ppgen1/n19 ), 
	.B2(n836), 
	.B1(n802), 
	.A2(n839), 
	.A1(n801));
   SEN_EO2_S_0P5 U2931 (.X(pprow0[10]), 
	.A2(\bmul/ppgen0/n34 ), 
	.A1(n827));
   SEN_AOI22_1 U2932 (.X(\bmul/ppgen0/n34 ), 
	.B2(n832), 
	.B1(B[9]), 
	.A2(n858), 
	.A1(n788));
   SEN_EO2_S_0P5 U2933 (.X(pprow0[23]), 
	.A2(\bmul/ppgen0/n20 ), 
	.A1(n828));
   SEN_AOI22_1 U2934 (.X(\bmul/ppgen0/n20 ), 
	.B2(n807), 
	.B1(n801), 
	.A2(n833), 
	.A1(n800));
   SEN_EO2_S_0P5 U2935 (.X(pprow0[24]), 
	.A2(\bmul/ppgen0/n19 ), 
	.A1(n828));
   SEN_AOI22_1 U2936 (.X(\bmul/ppgen0/n19 ), 
	.B2(A[0]), 
	.B1(n802), 
	.A2(n833), 
	.A1(n801));
   SEN_EO2_S_0P5 U2937 (.X(pprow0[25]), 
	.A2(\bmul/ppgen0/n18 ), 
	.A1(n828));
   SEN_AOI22_1 U2938 (.X(\bmul/ppgen0/n18 ), 
	.B2(A[0]), 
	.B1(n803), 
	.A2(n833), 
	.A1(n802));
   SEN_EO2_S_0P5 U2939 (.X(pprow0[26]), 
	.A2(\bmul/ppgen0/n17 ), 
	.A1(n828));
   SEN_AOI22_1 U2940 (.X(\bmul/ppgen0/n17 ), 
	.B2(A[0]), 
	.B1(n804), 
	.A2(n833), 
	.A1(n803));
   SEN_EO2_S_0P5 U2941 (.X(pprow0[27]), 
	.A2(\bmul/ppgen0/n16 ), 
	.A1(n828));
   SEN_AOI22_1 U2942 (.X(\bmul/ppgen0/n16 ), 
	.B2(A[0]), 
	.B1(n805), 
	.A2(n833), 
	.A1(n804));
   SEN_EO2_S_0P5 U2943 (.X(pprow0[28]), 
	.A2(\bmul/ppgen0/n15 ), 
	.A1(n828));
   SEN_AOI22_1 U2944 (.X(\bmul/ppgen0/n15 ), 
	.B2(A[0]), 
	.B1(n806), 
	.A2(n833), 
	.A1(n805));
   SEN_EO2_S_0P5 U2945 (.X(pprow3[10]), 
	.A2(n1892), 
	.A1(net84600));
   SEN_AOI22_1 U2946 (.X(n1892), 
	.B2(n823), 
	.B1(n786), 
	.A2(n845), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2947 (.X(pprow3[13]), 
	.A2(n1889), 
	.A1(net84600));
   SEN_AOI22_1 U2948 (.X(n1889), 
	.B2(n844), 
	.B1(n791), 
	.A2(n823), 
	.A1(n605));
   SEN_EO2_S_0P5 U2949 (.X(pprow3[14]), 
	.A2(n1888), 
	.A1(net84600));
   SEN_AOI22_1 U2950 (.X(n1888), 
	.B2(n844), 
	.B1(n792), 
	.A2(n823), 
	.A1(n609));
   SEN_EO2_S_0P5 U2951 (.X(pprow3[17]), 
	.A2(n1885), 
	.A1(net84600));
   SEN_AOI22_1 U2952 (.X(n1885), 
	.B2(n844), 
	.B1(n795), 
	.A2(n823), 
	.A1(n794));
   SEN_EO2_S_0P5 U2953 (.X(pprow3[18]), 
	.A2(n1884), 
	.A1(net84600));
   SEN_AOI22_1 U2954 (.X(n1884), 
	.B2(n844), 
	.B1(n796), 
	.A2(n823), 
	.A1(n795));
   SEN_EO2_S_0P5 U2955 (.X(pprow3[20]), 
	.A2(n1881), 
	.A1(net84600));
   SEN_AOI22_1 U2956 (.X(n1881), 
	.B2(n844), 
	.B1(n798), 
	.A2(n823), 
	.A1(n797));
   SEN_EO2_S_0P5 U2957 (.X(pprow3[21]), 
	.A2(n1880), 
	.A1(net84600));
   SEN_AOI22_1 U2958 (.X(n1880), 
	.B2(n844), 
	.B1(n799), 
	.A2(n823), 
	.A1(n798));
   SEN_EO2_S_0P5 U2959 (.X(pprow2[10]), 
	.A2(n1868), 
	.A1(n825));
   SEN_AOI22_1 U2960 (.X(n1868), 
	.B2(n842), 
	.B1(n786), 
	.A2(n841), 
	.A1(n788));
   SEN_EO2_S_0P5 U2961 (.X(pprow2[11]), 
	.A2(n1867), 
	.A1(n825));
   SEN_AOI22_1 U2962 (.X(n1867), 
	.B2(n840), 
	.B1(n789), 
	.A2(n842), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U2963 (.X(pprow2[12]), 
	.A2(n1866), 
	.A1(n825));
   SEN_AOI22_1 U2964 (.X(n1866), 
	.B2(n840), 
	.B1(n790), 
	.A2(n842), 
	.A1(n789));
   SEN_EO2_S_0P5 U2965 (.X(pprow2[13]), 
	.A2(n1865), 
	.A1(n825));
   SEN_AOI22_1 U2966 (.X(n1865), 
	.B2(n840), 
	.B1(n791), 
	.A2(n842), 
	.A1(n605));
   SEN_EO2_S_0P5 U2967 (.X(pprow2[14]), 
	.A2(n1864), 
	.A1(n825));
   SEN_AOI22_1 U2968 (.X(n1864), 
	.B2(n840), 
	.B1(n792), 
	.A2(n842), 
	.A1(n609));
   SEN_EO2_S_0P5 U2969 (.X(pprow2[15]), 
	.A2(n1863), 
	.A1(n825));
   SEN_AOI22_1 U2970 (.X(n1863), 
	.B2(n840), 
	.B1(n793), 
	.A2(n842), 
	.A1(n792));
   SEN_EO2_S_0P5 U2971 (.X(pprow2[16]), 
	.A2(n1862), 
	.A1(n825));
   SEN_AOI22_1 U2972 (.X(n1862), 
	.B2(n840), 
	.B1(n794), 
	.A2(n842), 
	.A1(n793));
   SEN_EO2_S_0P5 U2973 (.X(pprow2[17]), 
	.A2(n1861), 
	.A1(n825));
   SEN_AOI22_1 U2974 (.X(n1861), 
	.B2(n840), 
	.B1(n795), 
	.A2(n842), 
	.A1(n794));
   SEN_EO2_S_0P5 U2975 (.X(pprow2[18]), 
	.A2(n1860), 
	.A1(n825));
   SEN_AOI22_1 U2976 (.X(n1860), 
	.B2(n840), 
	.B1(n796), 
	.A2(n842), 
	.A1(n795));
   SEN_EO2_S_0P5 U2977 (.X(pprow2[19]), 
	.A2(n1859), 
	.A1(n825));
   SEN_AOI22_1 U2978 (.X(n1859), 
	.B2(n840), 
	.B1(n797), 
	.A2(n842), 
	.A1(n796));
   SEN_EO2_S_0P5 U2979 (.X(pprow2[20]), 
	.A2(n1857), 
	.A1(n825));
   SEN_AOI22_0P5 U2980 (.X(n1857), 
	.B2(n840), 
	.B1(n798), 
	.A2(n842), 
	.A1(n797));
   SEN_EO2_S_0P5 U2981 (.X(pprow2[21]), 
	.A2(n1856), 
	.A1(n825));
   SEN_AOI22_0P5 U2982 (.X(n1856), 
	.B2(n840), 
	.B1(n799), 
	.A2(n842), 
	.A1(n798));
   SEN_EO2_S_0P5 U2983 (.X(pprow7[7]), 
	.A2(n1956), 
	.A1(n818));
   SEN_AOI22_1 U2984 (.X(n1956), 
	.B2(\bmul/one7 ), 
	.B1(B[7]), 
	.A2(\bmul/two7 ), 
	.A1(B[6]));
   SEN_EO2_S_0P5 U2985 (.X(pprow2[7]), 
	.A2(n1846), 
	.A1(n826));
   SEN_AOI22_1 U2986 (.X(n1846), 
	.B2(n841), 
	.B1(B[7]), 
	.A2(n843), 
	.A1(B[6]));
   SEN_EO2_S_0P5 U2987 (.X(pprow2[8]), 
	.A2(n1845), 
	.A1(n826));
   SEN_AOI22_1 U2988 (.X(n1845), 
	.B2(n784), 
	.B1(n841), 
	.A2(n843), 
	.A1(n615));
   SEN_EO2_S_0P5 U2989 (.X(pprow2[9]), 
	.A2(n1844), 
	.A1(n826));
   SEN_AOI22_1 U2990 (.X(n1844), 
	.B2(n786), 
	.B1(n841), 
	.A2(B[8]), 
	.A1(n843));
   SEN_EO2_S_0P5 U2991 (.X(pprow2[22]), 
	.A2(n1855), 
	.A1(n826));
   SEN_AOI22_0P5 U2992 (.X(n1855), 
	.B2(n840), 
	.B1(n800), 
	.A2(n842), 
	.A1(n799));
   SEN_EO2_S_0P5 U2993 (.X(pprow2[24]), 
	.A2(n1853), 
	.A1(n826));
   SEN_AOI22_1 U2994 (.X(n1853), 
	.B2(n841), 
	.B1(n802), 
	.A2(n843), 
	.A1(n801));
   SEN_EO2_S_0P5 U2995 (.X(pprow2[25]), 
	.A2(n1852), 
	.A1(n826));
   SEN_AOI22_1 U2996 (.X(n1852), 
	.B2(n841), 
	.B1(n803), 
	.A2(n843), 
	.A1(n802));
   SEN_EO2_S_0P5 U2997 (.X(pprow3[7]), 
	.A2(n1872), 
	.A1(n202));
   SEN_AOI22_1 U2998 (.X(n1872), 
	.B2(n845), 
	.B1(B[7]), 
	.A2(n823), 
	.A1(n856));
   SEN_EO2_S_0P5 U2999 (.X(pprow3[9]), 
	.A2(n1870), 
	.A1(n202));
   SEN_AOI22_1 U3000 (.X(n1870), 
	.B2(n786), 
	.B1(n845), 
	.A2(B[8]), 
	.A1(n822));
   SEN_EO2_S_0P5 U3001 (.X(pprow0[8]), 
	.A2(\bmul/ppgen0/n4 ), 
	.A1(n1843));
   SEN_AOI22_1 U3002 (.X(\bmul/ppgen0/n4 ), 
	.B2(n784), 
	.B1(n858), 
	.A2(n834), 
	.A1(B[7]));
   SEN_EO2_S_0P5 U3003 (.X(pprow0[9]), 
	.A2(\bmul/ppgen0/n3 ), 
	.A1(n828));
   SEN_AOI22_1 U3004 (.X(\bmul/ppgen0/n3 ), 
	.B2(n786), 
	.B1(n858), 
	.A2(B[8]), 
	.A1(n834));
   SEN_EO2_S_0P5 U3005 (.X(pprow1[8]), 
	.A2(\bmul/ppgen1/n3 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U3006 (.X(\bmul/ppgen1/n3 ), 
	.B2(n784), 
	.B1(n837), 
	.A2(n839), 
	.A1(B[7]));
   SEN_ND4B_1 U3007 (.X(n962), 
	.B3(n996), 
	.B2(n291), 
	.B1(n961), 
	.A(n1195));
   SEN_EO2_S_0P5 U3008 (.X(Z[4]), 
	.A2(net84404), 
	.A1(n809));
   SEN_OAI21_S_0P5 U3009 (.X(n951), 
	.B(net84067), 
	.A2(n938), 
	.A1(n939));
   SEN_EO2_S_0P5 U3010 (.X(pprow4[9]), 
	.A2(n1894), 
	.A1(n614));
   SEN_AOI22_0P5 U3011 (.X(n1894), 
	.B2(n786), 
	.B1(n773), 
	.A2(n784), 
	.A1(\bmul/two4 ));
   SEN_EO2_S_0P5 U3012 (.X(pprow3[8]), 
	.A2(n1871), 
	.A1(n202));
   SEN_AOI22_1 U3013 (.X(n1871), 
	.B2(n784), 
	.B1(n845), 
	.A2(n822), 
	.A1(n615));
   SEN_EO2_S_0P5 U3014 (.X(pprow3[11]), 
	.A2(n1891), 
	.A1(net84600));
   SEN_AOI22_1 U3015 (.X(n1891), 
	.B2(n844), 
	.B1(n789), 
	.A2(n822), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U3016 (.X(pprow3[12]), 
	.A2(n1890), 
	.A1(net84600));
   SEN_AOI22_1 U3017 (.X(n1890), 
	.B2(n844), 
	.B1(n790), 
	.A2(n822), 
	.A1(n610));
   SEN_EO2_S_0P5 U3018 (.X(pprow3[15]), 
	.A2(n1887), 
	.A1(net84600));
   SEN_AOI22_1 U3019 (.X(n1887), 
	.B2(n844), 
	.B1(n793), 
	.A2(n822), 
	.A1(n792));
   SEN_EO2_S_0P5 U3020 (.X(pprow3[16]), 
	.A2(n1886), 
	.A1(net84600));
   SEN_AOI22_1 U3021 (.X(n1886), 
	.B2(n844), 
	.B1(n794), 
	.A2(n822), 
	.A1(n793));
   SEN_EO2_S_0P5 U3022 (.X(pprow3[19]), 
	.A2(n1883), 
	.A1(net84600));
   SEN_AOI22_1 U3023 (.X(n1883), 
	.B2(n844), 
	.B1(n797), 
	.A2(n822), 
	.A1(n796));
   SEN_EO2_S_0P5 U3024 (.X(pprow3[22]), 
	.A2(n1879), 
	.A1(n202));
   SEN_AOI22_1 U3025 (.X(n1879), 
	.B2(n844), 
	.B1(n800), 
	.A2(n822), 
	.A1(n799));
   SEN_EO2_S_0P5 U3026 (.X(pprow3[23]), 
	.A2(n1878), 
	.A1(n202));
   SEN_AOI22_1 U3027 (.X(n1878), 
	.B2(n845), 
	.B1(n801), 
	.A2(n822), 
	.A1(n800));
   SEN_EO2_S_0P5 U3028 (.X(pprow1[11]), 
	.A2(\bmul/ppgen1/n33 ), 
	.A1(net84586));
   SEN_AOI22_T_0P5 U3029 (.X(\bmul/ppgen1/n33 ), 
	.B2(n835), 
	.B1(n789), 
	.A2(n838), 
	.A1(n788));
   SEN_EO2_S_0P5 U3030 (.X(pprow1[13]), 
	.A2(\bmul/ppgen1/n31 ), 
	.A1(net84586));
   SEN_AOI22_T_0P5 U3031 (.X(\bmul/ppgen1/n31 ), 
	.B2(n835), 
	.B1(n791), 
	.A2(n838), 
	.A1(n790));
   SEN_EO2_S_0P5 U3032 (.X(pprow1[15]), 
	.A2(\bmul/ppgen1/n29 ), 
	.A1(net84586));
   SEN_AOI22_0P5 U3033 (.X(\bmul/ppgen1/n29 ), 
	.B2(n836), 
	.B1(n793), 
	.A2(n838), 
	.A1(n792));
   SEN_EO2_S_0P5 U3034 (.X(pprow1[20]), 
	.A2(\bmul/ppgen1/n23 ), 
	.A1(net84586));
   SEN_AOI22_1 U3035 (.X(\bmul/ppgen1/n23 ), 
	.B2(n835), 
	.B1(n798), 
	.A2(n838), 
	.A1(n797));
   SEN_EO2_S_0P5 U3036 (.X(pprow1[23]), 
	.A2(\bmul/ppgen1/n20 ), 
	.A1(net84588));
   SEN_AOI22_1 U3037 (.X(\bmul/ppgen1/n20 ), 
	.B2(n835), 
	.B1(n801), 
	.A2(n839), 
	.A1(n800));
   SEN_EO2_S_0P5 U3038 (.X(pprow1[25]), 
	.A2(\bmul/ppgen1/n18 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U3039 (.X(\bmul/ppgen1/n18 ), 
	.B2(n836), 
	.B1(n803), 
	.A2(n839), 
	.A1(n802));
   SEN_EO2_S_0P5 U3040 (.X(pprow1[26]), 
	.A2(\bmul/ppgen1/n17 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U3041 (.X(\bmul/ppgen1/n17 ), 
	.B2(n836), 
	.B1(n804), 
	.A2(n839), 
	.A1(n803));
   SEN_EO2_S_0P5 U3042 (.X(pprow1[27]), 
	.A2(\bmul/ppgen1/n16 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U3043 (.X(\bmul/ppgen1/n16 ), 
	.B2(n836), 
	.B1(n805), 
	.A2(n839), 
	.A1(n804));
   SEN_EO2_S_0P5 U3044 (.X(pprow1[28]), 
	.A2(\bmul/ppgen1/n15 ), 
	.A1(net84588));
   SEN_AOI22_0P5 U3045 (.X(\bmul/ppgen1/n15 ), 
	.B2(n836), 
	.B1(n806), 
	.A2(n839), 
	.A1(n805));
   SEN_EO2_S_0P5 U3046 (.X(pprow0[11]), 
	.A2(\bmul/ppgen0/n33 ), 
	.A1(n827));
   SEN_AOI22_1 U3047 (.X(\bmul/ppgen0/n33 ), 
	.B2(n858), 
	.B1(n789), 
	.A2(n832), 
	.A1(B[10]));
   SEN_EO2_S_0P5 U3048 (.X(pprow0[12]), 
	.A2(\bmul/ppgen0/n32 ), 
	.A1(n827));
   SEN_AOI22_1 U3049 (.X(\bmul/ppgen0/n32 ), 
	.B2(n858), 
	.B1(n790), 
	.A2(n832), 
	.A1(n610));
   SEN_EO2_S_0P5 U3050 (.X(pprow0[13]), 
	.A2(\bmul/ppgen0/n31 ), 
	.A1(n827));
   SEN_AOI22_1 U3051 (.X(\bmul/ppgen0/n31 ), 
	.B2(n858), 
	.B1(n791), 
	.A2(n832), 
	.A1(n605));
   SEN_EO2_S_0P5 U3052 (.X(pprow0[14]), 
	.A2(\bmul/ppgen0/n30 ), 
	.A1(n827));
   SEN_AOI22_1 U3053 (.X(\bmul/ppgen0/n30 ), 
	.B2(n807), 
	.B1(n792), 
	.A2(n832), 
	.A1(n609));
   SEN_EO2_S_0P5 U3054 (.X(pprow0[15]), 
	.A2(\bmul/ppgen0/n29 ), 
	.A1(n827));
   SEN_AOI22_1 U3055 (.X(\bmul/ppgen0/n29 ), 
	.B2(A[0]), 
	.B1(n793), 
	.A2(n832), 
	.A1(n792));
   SEN_EO2_S_0P5 U3056 (.X(pprow0[16]), 
	.A2(\bmul/ppgen0/n28 ), 
	.A1(n827));
   SEN_AOI22_1 U3057 (.X(\bmul/ppgen0/n28 ), 
	.B2(A[0]), 
	.B1(n794), 
	.A2(n832), 
	.A1(n793));
   SEN_EO2_S_0P5 U3058 (.X(pprow0[17]), 
	.A2(\bmul/ppgen0/n27 ), 
	.A1(n827));
   SEN_AOI22_1 U3059 (.X(\bmul/ppgen0/n27 ), 
	.B2(A[0]), 
	.B1(n795), 
	.A2(n832), 
	.A1(n794));
   SEN_EO2_S_0P5 U3060 (.X(pprow0[18]), 
	.A2(\bmul/ppgen0/n26 ), 
	.A1(n827));
   SEN_AOI22_1 U3061 (.X(\bmul/ppgen0/n26 ), 
	.B2(A[0]), 
	.B1(n796), 
	.A2(n832), 
	.A1(n795));
   SEN_EO2_S_0P5 U3062 (.X(pprow0[19]), 
	.A2(\bmul/ppgen0/n25 ), 
	.A1(n827));
   SEN_AOI22_1 U3063 (.X(\bmul/ppgen0/n25 ), 
	.B2(A[0]), 
	.B1(n797), 
	.A2(n832), 
	.A1(n796));
   SEN_EO2_S_0P5 U3064 (.X(pprow0[20]), 
	.A2(\bmul/ppgen0/n23 ), 
	.A1(n827));
   SEN_AOI22_1 U3065 (.X(\bmul/ppgen0/n23 ), 
	.B2(n858), 
	.B1(n798), 
	.A2(n832), 
	.A1(n797));
   SEN_EO2_S_0P5 U3066 (.X(pprow0[21]), 
	.A2(\bmul/ppgen0/n22 ), 
	.A1(n827));
   SEN_AOI22_1 U3067 (.X(\bmul/ppgen0/n22 ), 
	.B2(A[0]), 
	.B1(n799), 
	.A2(n832), 
	.A1(n798));
   SEN_EO2_S_0P5 U3068 (.X(pprow0[22]), 
	.A2(\bmul/ppgen0/n21 ), 
	.A1(n828));
   SEN_AOI22_1 U3069 (.X(\bmul/ppgen0/n21 ), 
	.B2(n858), 
	.B1(n800), 
	.A2(n832), 
	.A1(n799));
   SEN_EO2_S_0P5 U3070 (.X(pprow2[23]), 
	.A2(n1854), 
	.A1(n826));
   SEN_AOI22_1 U3071 (.X(n1854), 
	.B2(n841), 
	.B1(n801), 
	.A2(n843), 
	.A1(n800));
   SEN_EO2_S_0P5 U3072 (.X(pprow1[10]), 
	.A2(\bmul/ppgen1/n34 ), 
	.A1(net84586));
   SEN_AOI22_0P5 U3073 (.X(\bmul/ppgen1/n34 ), 
	.B2(n838), 
	.B1(n786), 
	.A2(n837), 
	.A1(n788));
   SEN_EO2_S_0P5 U3074 (.X(pprow0[7]), 
	.A2(\bmul/ppgen0/n5 ), 
	.A1(n1843));
   SEN_AOI22_1 U3075 (.X(\bmul/ppgen0/n5 ), 
	.B2(A[0]), 
	.B1(n615), 
	.A2(n834), 
	.A1(n856));
   SEN_ND2_S_0P5 U3076 (.X(n1187), 
	.A2(n1146), 
	.A1(n1171));
   SEN_INV_1 U3077 (.X(n1780), 
	.A(n1776));
   SEN_ND2_S_0P5 U3078 (.X(n1540), 
	.A2(n1538), 
	.A1(n1539));
   SEN_EO2_S_0P5 U3079 (.X(pprow12[0]), 
	.A2(n2019), 
	.A1(n1489));
   SEN_ND2_G_1 U3080 (.X(n2019), 
	.A2(\bmul/one12 ), 
	.A1(n829));
   SEN_INV_2 U3081 (.X(n1227), 
	.A(n1231));
   SEN_INV_S_1 U3082 (.X(n1015), 
	.A(n811));
   SEN_EO2_S_0P5 U3083 (.X(pprow7[0]), 
	.A2(n1969), 
	.A1(n818));
   SEN_ND2_G_1 U3084 (.X(n1969), 
	.A2(n611), 
	.A1(n829));
   SEN_BUF_S_1 U3085 (.X(n823), 
	.A(\bmul/two3 ));
   SEN_NR2_S_0P5 U3086 (.X(\bmul/two3 ), 
	.A2(n2024), 
	.A1(n845));
   SEN_INV_2 U3087 (.X(n1746), 
	.A(n1750));
   SEN_INV_S_0P5 U3088 (.X(net2259), 
	.A(net84654));
   SEN_INV_S_1 U3089 (.X(n896), 
	.A(n893));
   SEN_BUF_S_1 U3090 (.X(n822), 
	.A(n821));
   SEN_NR2_S_0P5 U3091 (.X(n821), 
	.A2(n2024), 
	.A1(n845));
   SEN_INV_S_1 U3092 (.X(n836), 
	.A(n755));
   SEN_INV_1 U3093 (.X(n1013), 
	.A(n1014));
   SEN_BUF_S_1 U3094 (.X(n859), 
	.A(n860));
   SEN_AO21_1 U3095 (.X(n921), 
	.B(n938), 
	.A2(n915), 
	.A1(n614));
   SEN_AO21_DG_1 U3096 (.X(net82772), 
	.B(n1536), 
	.A2(n1488), 
	.A1(n1489));
   SEN_ND2_G_1 U3097 (.X(n1431), 
	.A2(n1428), 
	.A1(n1429));
   SEN_INV_S_1 U3098 (.X(n843), 
	.A(n764));
   SEN_INV_S_1 U3099 (.X(n938), 
	.A(n914));
   SEN_INV_0P8 U3100 (.X(n773), 
	.A(n771));
   SEN_INV_S_1 U3101 (.X(n829), 
	.A(n831));
   SEN_INV_S_0P5 U3102 (.X(n837), 
	.A(n755));
   SEN_AN2_S_0P5 U3103 (.X(net83644), 
	.A2(net83646), 
	.A1(net83645));
   SEN_EO2_S_0P5 U3104 (.X(pprow1[9]), 
	.A2(\bmul/ppgen1/n2 ), 
	.A1(net84586));
   SEN_AOI22_1 U3105 (.X(\bmul/ppgen1/n2 ), 
	.B2(n786), 
	.B1(n837), 
	.A2(n784), 
	.A1(n839));
   SEN_INV_S_1 U3106 (.X(net2268), 
	.A(net84636));
   SEN_EN2_0P5 U3107 (.X(\dp_cluster_0/N288 ), 
	.A2(n861), 
	.A1(n808));
   SEN_INV_S_0P5 U3108 (.X(n1840), 
	.A(n437));
   SEN_INV_S_0P5 U3109 (.X(n1839), 
	.A(n813));
   SEN_INV_S_1 U3110 (.X(n788), 
	.A(n787));
   SEN_AN2_S_1 U3111 (.X(n1693), 
	.A2(pprow11_qual[3]), 
	.A1(pprow10_qual[5]));
   SEN_EN2_0P5 U3112 (.X(n2032), 
	.A2(net84634), 
	.A1(A[22]));
   SEN_EO2_S_0P5 U3113 (.X(n707), 
	.A2(pprow5_qual[8]), 
	.A1(pprow4_qual[10]));
   SEN_EO2_S_0P5 U3114 (.X(n710), 
	.A2(pprow1_qual[18]), 
	.A1(pprow1_qual[20]));
   SEN_EO2_S_0P5 U3115 (.X(n1685), 
	.A2(pprow7_qual[12]), 
	.A1(pprow6_qual[14]));
   SEN_EO2_S_0P5 U3116 (.X(n711), 
	.A2(pprow9_qual[8]), 
	.A1(pprow8_qual[10]));
   SEN_NR2_1 U3117 (.X(\bmul/two12 ), 
	.A2(n2033), 
	.A1(\bmul/one12 ));
   SEN_EN2_0P5 U3118 (.X(n2033), 
	.A2(n815), 
	.A1(A[24]));
   SEN_EO2_S_0P5 U3119 (.X(n717), 
	.A2(pprow3_qual[22]), 
	.A1(pprow2_qual[24]));
   SEN_EO2_S_0P5 U3120 (.X(n1470), 
	.A2(pprow7_qual[8]), 
	.A1(pprow6_qual[10]));
   SEN_EN2_0P5 U3121 (.X(n2026), 
	.A2(n399), 
	.A1(A[10]));
   SEN_EO2_S_0P5 U3122 (.X(n993), 
	.A2(C[12]), 
	.A1(net84026));
   SEN_EN2_0P5 U3123 (.X(n2024), 
	.A2(net90815), 
	.A1(A[6]));
   SEN_INV_S_0P5 U3124 (.X(n1220), 
	.A(n1239));
   SEN_EN2_0P5 U3125 (.X(n1303), 
	.A2(pprow9_qual[0]), 
	.A1(pprow8_qual[2]));
   SEN_EO2_2 U3126 (.X(n1475), 
	.A2(n1468), 
	.A1(n1402));
   SEN_EN2_0P5 U3127 (.X(n1402), 
	.A2(pprow9_qual[3]), 
	.A1(pprow8_qual[5]));
   SEN_EO2_S_0P5 U3128 (.X(n718), 
	.A2(pprow9_qual[4]), 
	.A1(pprow8_qual[6]));
   SEN_EO2_S_0P5 U3129 (.X(n1591), 
	.A2(pprow11_qual[2]), 
	.A1(pprow10_qual[4]));
   SEN_EN2_0P5 U3130 (.X(n719), 
	.A2(pprow11_qual[5]), 
	.A1(pprow10_qual[7]));
   SEN_EO2_S_0P5 U3131 (.X(n720), 
	.A2(pprow9_qual[2]), 
	.A1(pprow8_qual[4]));
   SEN_EO2_S_0P5 U3132 (.X(n722), 
	.A2(pprow1_qual[13]), 
	.A1(pprow1_qual[15]));
   SEN_EO2_S_0P5 U3133 (.X(\bmul/one14 ), 
	.A2(n816), 
	.A1(A[28]));
   SEN_EO2_S_0P5 U3134 (.X(n723), 
	.A2(pprow5_qual[11]), 
	.A1(pprow4_qual[13]));
   SEN_EO2_1 U3135 (.X(n724), 
	.A2(pprow5_qual[1]), 
	.A1(pprow4_qual[3]));
   SEN_EN2_0P5 U3136 (.X(n2027), 
	.A2(n811), 
	.A1(A[12]));
   SEN_EN2_0P5 U3137 (.X(n728), 
	.A2(pprow9_qual[9]), 
	.A1(pprow8_qual[11]));
   SEN_EO2_S_0P5 U3138 (.X(n1181), 
	.A2(pprow5_qual[5]), 
	.A1(pprow4_qual[7]));
   SEN_EO2_S_0P5 U3139 (.X(n731), 
	.A2(pprow11_qual[3]), 
	.A1(pprow10_qual[5]));
   SEN_EN2_0P5 U3140 (.X(n912), 
	.A2(n530), 
	.A1(n527));
   SEN_EO2_S_0P5 U3141 (.X(n732), 
	.A2(pprow9_qual[5]), 
	.A1(pprow8_qual[7]));
   SEN_EO2_S_0P5 U3142 (.X(n733), 
	.A2(pprow7_qual[14]), 
	.A1(pprow6_qual[16]));
   SEN_EN2_0P5 U3143 (.X(n974), 
	.A2(pprow1_qual[7]), 
	.A1(pprow1_qual[9]));
   SEN_EO2_S_0P5 U3144 (.X(n1791), 
	.A2(C[29]), 
	.A1(n1789));
   SEN_EO2_S_0P5 U3145 (.X(n734), 
	.A2(pprow11_qual[6]), 
	.A1(pprow10_qual[8]));
   SEN_AN2_1 U3146 (.X(n1589), 
	.A2(pprow11_qual[1]), 
	.A1(pprow10_qual[3]));
   SEN_EO2_S_0P5 U3147 (.X(n735), 
	.A2(pprow9_qual[6]), 
	.A1(pprow8_qual[8]));
   SEN_EN2_0P5 U3148 (.X(n2028), 
	.A2(n437), 
	.A1(A[14]));
   SEN_AN2_S_1 U3149 (.X(net82486), 
	.A2(pprow7_qual[11]), 
	.A1(pprow6_qual[13]));
   SEN_INV_S_0P5 U3150 (.X(n1110), 
	.A(n1190));
   SEN_AN2_S_1 U3151 (.X(n1498), 
	.A2(pprow9_qual[4]), 
	.A1(pprow8_qual[6]));
   SEN_EO2_S_0P5 U3152 (.X(n739), 
	.A2(pprow7_qual[13]), 
	.A1(pprow6_qual[15]));
   SEN_AN2_S_1 U3153 (.X(n1669), 
	.A2(pprow5_qual[15]), 
	.A1(pprow4_qual[17]));
   SEN_ND2_G_1 U3154 (.X(n1761), 
	.A2(C[28]), 
	.A1(pprow0_qual[28]));
   SEN_AN2_S_1 U3155 (.X(n1717), 
	.A2(pprow9_qual[8]), 
	.A1(pprow8_qual[10]));
   SEN_EO2_S_0P5 U3156 (.X(n1695), 
	.A2(pprow11_qual[4]), 
	.A1(pprow10_qual[6]));
   SEN_EN2_0P5 U3157 (.X(n888), 
	.A2(net90815), 
	.A1(pprow2_qual[0]));
   SEN_EO2_S_0P5 U3158 (.X(n1750), 
	.A2(n1691), 
	.A1(n1692));
   SEN_EN2_0P5 U3159 (.X(n1692), 
	.A2(pprow13_qual[0]), 
	.A1(pprow12_qual[2]));
   SEN_EN2_0P5 U3160 (.X(net82181), 
	.A2(\bmul/neg15 ), 
	.A1(pprow14_qual[0]));
   SEN_EO2_S_0P5 U3161 (.X(n1609), 
	.A2(pprow9_qual[7]), 
	.A1(pprow8_qual[9]));
   SEN_EN2_0P5 U3162 (.X(n2029), 
	.A2(n813), 
	.A1(A[16]));
   SEN_NR2_1 U3163 (.X(\bmul/two13 ), 
	.A2(n2034), 
	.A1(\bmul/one13 ));
   SEN_EN2_0P5 U3164 (.X(n2034), 
	.A2(n816), 
	.A1(A[26]));
   SEN_EO2_S_0P5 U3165 (.X(n1671), 
	.A2(pprow5_qual[16]), 
	.A1(pprow4_qual[18]));
   SEN_EN2_0P5 U3166 (.X(n865), 
	.A2(pprow1_qual[0]), 
	.A1(pprow1_qual[2]));
   SEN_EN2_0P5 U3167 (.X(n1087), 
	.A2(n255), 
	.A1(pprow4_qual[5]));
   SEN_EN2_0P5 U3168 (.X(n1077), 
	.A2(n437), 
	.A1(pprow6_qual[0]));
   SEN_INV_S_1 U3169 (.X(n1763), 
	.A(C[28]));
   SEN_INV_S_1 U3170 (.X(n1534), 
	.A(pprow11_qual[0]));
   SEN_ND2_G_1 U3171 (.X(n1681), 
	.A2(pprow9_qual[7]), 
	.A1(pprow8_qual[9]));
   SEN_INV_S_1 U3172 (.X(n1684), 
	.A(pprow8_qual[9]));
   SEN_ND2_G_1 U3173 (.X(n1556), 
	.A2(pprow9_qual[5]), 
	.A1(pprow8_qual[7]));
   SEN_ND2_G_1 U3174 (.X(n1719), 
	.A2(pprow7_qual[12]), 
	.A1(pprow6_qual[14]));
   SEN_INV_S_1 U3175 (.X(n1721), 
	.A(pprow6_qual[14]));
   SEN_INV_S_1 U3176 (.X(n1720), 
	.A(pprow7_qual[12]));
   SEN_EN2_0P5 U3177 (.X(n2030), 
	.A2(n814), 
	.A1(A[18]));
   SEN_ND2_G_1 U3178 (.X(n1601), 
	.A2(n561), 
	.A1(n1599));
   SEN_ND2_G_1 U3179 (.X(n1706), 
	.A2(n1703), 
	.A1(n1704));
   SEN_EO2_S_0P5 U3180 (.X(pprow14[1]), 
	.A2(\bmul/ppgen14/n24 ), 
	.A1(n1836));
   SEN_AOI22_1 U3181 (.X(\bmul/ppgen14/n24 ), 
	.B2(\bmul/one14 ), 
	.B1(n846), 
	.A2(\bmul/two14 ), 
	.A1(n830));
   SEN_NR2_1 U3182 (.X(\bmul/two14 ), 
	.A2(n2035), 
	.A1(\bmul/one14 ));
   SEN_EN2_0P5 U3183 (.X(n2035), 
	.A2(\bmul/neg14 ), 
	.A1(A[28]));
   SEN_AN2_S_1 U3184 (.X(n1792), 
	.A2(pprow7_qual[13]), 
	.A1(pprow6_qual[15]));
   SEN_ND2_G_1 U3185 (.X(n1812), 
	.A2(pprow7_qual[14]), 
	.A1(pprow6_qual[16]));
   SEN_INV_S_1 U3186 (.X(n1815), 
	.A(pprow6_qual[16]));
   SEN_INV_S_1 U3187 (.X(n1814), 
	.A(pprow7_qual[14]));
   SEN_ND2_G_1 U3188 (.X(n1639), 
	.A2(C[26]), 
	.A1(pprow0_qual[26]));
   SEN_OR2_1 U3189 (.X(n748), 
	.A2(pprow4_qual[12]), 
	.A1(pprow5_qual[10]));
   SEN_EN2_0P5 U3190 (.X(n1168), 
	.A2(pprow7_qual[1]), 
	.A1(pprow6_qual[3]));
   SEN_EN2_0P5 U3191 (.X(n2031), 
	.A2(net84636), 
	.A1(A[20]));
   SEN_EO2_S_0P5 U3192 (.X(pprow1[29]), 
	.A2(\bmul/ppgen1/n14 ), 
	.A1(net84588));
   SEN_AOI22_1 U3193 (.X(\bmul/ppgen1/n14 ), 
	.B2(n836), 
	.B1(B[29]), 
	.A2(n839), 
	.A1(n806));
   SEN_EO2_S_0P5 U3194 (.X(pprow0[29]), 
	.A2(\bmul/ppgen0/n14 ), 
	.A1(n828));
   SEN_AOI22_1 U3195 (.X(\bmul/ppgen0/n14 ), 
	.B2(A[0]), 
	.B1(B[29]), 
	.A2(n833), 
	.A1(n806));
   SEN_EO2_S_0P5 U3196 (.X(pprow0[30]), 
	.A2(\bmul/ppgen0/n12 ), 
	.A1(n828));
   SEN_AOI22_1 U3197 (.X(\bmul/ppgen0/n12 ), 
	.B2(A[0]), 
	.B1(B[30]), 
	.A2(n833), 
	.A1(B[29]));
   SEN_EO2_S_0P5 U3198 (.X(pprow0[31]), 
	.A2(\bmul/ppgen0/n11 ), 
	.A1(n828));
   SEN_AOI22_1 U3199 (.X(\bmul/ppgen0/n11 ), 
	.B2(n807), 
	.B1(B[31]), 
	.A2(n833), 
	.A1(B[30]));
   SEN_ND2_G_1 U3200 (.X(n1800), 
	.A2(n1797), 
	.A1(n1798));
   SEN_OR2_1 U3201 (.X(net82701), 
	.A2(pprow3_qual[15]), 
	.A1(pprow2_qual[17]));
   SEN_EN2_0P5 U3202 (.X(n751), 
	.A2(pprow13_qual[2]), 
	.A1(pprow12_qual[4]));
   SEN_ND2_G_1 U3203 (.X(n1788), 
	.A2(pprow0_qual[29]), 
	.A1(C[29]));
   SEN_INV_S_1 U3204 (.X(n1790), 
	.A(C[29]));
   SEN_ND2_G_1 U3205 (.X(n1801), 
	.A2(pprow4_qual[19]), 
	.A1(pprow5_qual[17]));
   SEN_OR2_1 U3206 (.X(n754), 
	.A2(pprow4_qual[13]), 
	.A1(pprow5_qual[11]));
   SEN_EN2_0P5 U3207 (.X(n755), 
	.A2(n808), 
	.A1(A[2]));
   SEN_ND2_S_0P5 U3208 (.X(n1361), 
	.A2(n525), 
	.A1(pprow1_qual[18]));
   SEN_ND2_G_1 U3209 (.X(net82166), 
	.A2(pprow0_qual[30]), 
	.A1(C[30]));
   SEN_INV_S_1 U3211 (.X(n1732), 
	.A(pprow2_qual[22]));
   SEN_INV_S_1 U3212 (.X(n1803), 
	.A(pprow4_qual[19]));
   SEN_ND2_G_1 U3213 (.X(n1731), 
	.A2(pprow2_qual[22]), 
	.A1(pprow3_qual[20]));
   SEN_EN2_0P5 U3214 (.X(n758), 
	.A2(pprow9_qual[10]), 
	.A1(pprow8_qual[12]));
   SEN_INV_S_1 U3215 (.X(net82163), 
	.A(C[30]));
   SEN_INV_S_1 U3216 (.X(n1258), 
	.A(n1292));
   SEN_EO2_S_0P5 U3217 (.X(n759), 
	.A2(pprow1_qual[21]), 
	.A1(pprow1_qual[23]));
   SEN_AO21_1 U3218 (.X(n1690), 
	.B(n1691), 
	.A2(n1637), 
	.A1(n1638));
   SEN_INV_S_1 U3219 (.X(n1638), 
	.A(pprow12_qual[1]));
   SEN_EN2_0P5 U3220 (.X(n760), 
	.A2(net84654), 
	.A1(A[4]));
   SEN_EN2_0P5 U3221 (.X(n761), 
	.A2(n809), 
	.A1(A[6]));
   SEN_ND2_G_1 U3222 (.X(n1794), 
	.A2(pprow9_qual[9]), 
	.A1(pprow8_qual[11]));
   SEN_NR2_1 U3223 (.X(n1795), 
	.A2(pprow8_qual[11]), 
	.A1(pprow9_qual[9]));
   SEN_ND2B_1 U3224 (.X(n762), 
	.B(n763), 
	.A(n837));
   SEN_INV_S_1 U3225 (.X(net82511), 
	.A(pprow2_qual[21]));
   SEN_INV_2 U3226 (.X(n1166), 
	.A(n1101));
   SEN_INV_S_1 U3227 (.X(n1797), 
	.A(pprow2_qual[23]));
   SEN_INV_S_1 U3228 (.X(n1789), 
	.A(pprow0_qual[29]));
   SEN_INV_S_1 U3230 (.X(n1764), 
	.A(pprow0_qual[28]));
   SEN_INV_S_1 U3231 (.X(n1733), 
	.A(pprow3_qual[20]));
   SEN_INV_S_1 U3232 (.X(n1804), 
	.A(pprow5_qual[17]));
   SEN_ND2B_1 U3233 (.X(n764), 
	.B(n765), 
	.A(n841));
   SEN_EO2_S_0P5 U3234 (.X(n765), 
	.A2(n809), 
	.A1(A[4]));
   SEN_INV_S_2 U3236 (.X(n941), 
	.A(pprow2_qual[3]));
   SEN_INV_S_1 U3237 (.X(net82510), 
	.A(pprow3_qual[19]));
   SEN_OA21_2 U3238 (.X(n766), 
	.B(n1166), 
	.A2(pprow6_qual[2]), 
	.A1(pprow7_qual[0]));
   SEN_OR2_1 U3239 (.X(n1390), 
	.A2(pprow3_qual[13]), 
	.A1(pprow2_qual[15]));
   SEN_AO21_DG_1 U3240 (.X(n893), 
	.B(n913), 
	.A2(n934), 
	.A1(n892));
   SEN_INV_S_1 U3241 (.X(n1599), 
	.A(pprow0_qual[25]));
   SEN_INV_S_1 U3242 (.X(n1704), 
	.A(pprow0_qual[27]));
   SEN_INV_S_1 U3244 (.X(n1798), 
	.A(pprow3_qual[21]));
   SEN_ND2_G_1 U3245 (.X(net82130), 
	.A2(n1783), 
	.A1(n1784));
   SEN_OAI21_G_1 U3246 (.X(n1783), 
	.B(n1782), 
	.A2(pprow12_qual[3]), 
	.A1(pprow13_qual[1]));
   SEN_ND2_G_1 U3247 (.X(n1726), 
	.A2(pprow5_qual[16]), 
	.A1(pprow4_qual[18]));
   SEN_INV_S_1 U3248 (.X(n1729), 
	.A(pprow4_qual[18]));
   SEN_INV_S_0P5 U3249 (.X(n1029), 
	.A(pprow4_qual[1]));
   SEN_INV_S_1 U3250 (.X(n872), 
	.A(pprow0_qual[4]));
   SEN_INV_S_1 U3251 (.X(n1728), 
	.A(pprow5_qual[16]));
   SEN_INV_S_1 U3252 (.X(n1541), 
	.A(pprow0_qual[24]));
   SEN_OR2_DG_1 U3253 (.X(n770), 
	.A2(pprow1_qual[18]), 
	.A1(n525));
   SEN_EN2_0P5 U3254 (.X(n771), 
	.A2(net90815), 
	.A1(A[8]));
   SEN_BUF_S_1 U3255 (.X(n809), 
	.A(\bmul/neg2 ));
   SEN_INV_S_1 U3256 (.X(net82171), 
	.A(pprow1_qual[28]));
   SEN_INV_S_1 U3257 (.X(n847), 
	.A(B[1]));
   SEN_INV_S_1 U3258 (.X(n849), 
	.A(B[2]));
   SEN_INV_S_1 U3259 (.X(n851), 
	.A(B[3]));
   SEN_INV_S_1 U3260 (.X(n853), 
	.A(B[4]));
   SEN_INV_S_1 U3261 (.X(n855), 
	.A(B[5]));
   SEN_INV_S_1 U3262 (.X(n857), 
	.A(B[6]));
   SEN_OR2_1 U3263 (.X(net85748), 
	.A2(pprow1_qual[28]), 
	.A1(pprow1_qual[26]));
   SEN_INV_S_1 U3264 (.X(n860), 
	.A(n807));
   SEN_BUF_S_1 U3265 (.X(n807), 
	.A(A[0]));
   SEN_INV_S_1 U3266 (.X(n831), 
	.A(\bmul/ppgen15/twoscomp[0] ));
   SEN_INV_S_1 U3267 (.X(n1836), 
	.A(\bmul/neg14 ));
   SEN_INV_S_1 U3268 (.X(n782), 
	.A(B[7]));
   SEN_INV_S_1 U3269 (.X(n785), 
	.A(B[9]));
   SEN_INV_S_1 U3270 (.X(n787), 
	.A(B[10]));
   SEN_INV_S_1 U3271 (.X(n783), 
	.A(B[8]));
   SEN_BUF_S_1 U3272 (.X(n792), 
	.A(B[14]));
   SEN_BUF_S_1 U3273 (.X(n793), 
	.A(B[15]));
   SEN_BUF_S_1 U3274 (.X(n794), 
	.A(B[16]));
   SEN_BUF_S_1 U3275 (.X(n795), 
	.A(B[17]));
   SEN_BUF_S_1 U3276 (.X(n796), 
	.A(B[18]));
   SEN_BUF_S_1 U3277 (.X(n797), 
	.A(B[19]));
   SEN_BUF_S_1 U3278 (.X(n798), 
	.A(B[20]));
   SEN_BUF_S_1 U3279 (.X(n799), 
	.A(B[21]));
   SEN_BUF_S_1 U3280 (.X(n800), 
	.A(B[22]));
   SEN_BUF_S_1 U3281 (.X(n801), 
	.A(B[23]));
   SEN_BUF_S_1 U3282 (.X(n802), 
	.A(B[24]));
   SEN_BUF_S_1 U3283 (.X(n803), 
	.A(B[25]));
   SEN_BUF_S_1 U3284 (.X(n804), 
	.A(B[26]));
   SEN_BUF_S_1 U3285 (.X(n805), 
	.A(B[27]));
   SEN_BUF_S_1 U3286 (.X(n806), 
	.A(B[28]));
   SEN_EN2_0P5 U3287 (.X(n1063), 
	.A2(pprow1_qual[10]), 
	.A1(pprow1_qual[12]));
   SEN_ND2_1P5 U3288 (.X(n1148), 
	.A2(pprow1_qual[8]), 
	.A1(pprow1_qual[10]));
   SEN_ND2_S_0P5 U3289 (.X(n1146), 
	.A2(n1145), 
	.A1(n1839));
   SEN_EN2_0P5 U3290 (.X(n883), 
	.A2(n887), 
	.A1(n886));
   SEN_EN3_0P5 U3291 (.X(Z[8]), 
	.A3(n464), 
	.A2(n916), 
	.A1(n917));
   SEN_EN3_0P5 U3292 (.X(Z[7]), 
	.A3(n895), 
	.A2(n893), 
	.A1(n258));
   SEN_NR2_S_0P5 U3293 (.X(n970), 
	.A2(n995), 
	.A1(n704));
   SEN_ND2_S_0P5 U3294 (.X(n779), 
	.A2(n876), 
	.A1(n904));
   SEN_INV_4 U3295 (.X(net82260), 
	.A(net82251));
   SEN_ND2B_6 U3296 (.X(n1506), 
	.B(n1504), 
	.A(n1505));
   SEN_AN3B_4 U3297 (.X(n1774), 
	.B2(n1767), 
	.B1(n384), 
	.A(n1766));
   SEN_EN2_0P5 U3298 (.X(n1115), 
	.A2(pprow1_qual[11]), 
	.A1(pprow1_qual[13]));
   SEN_ND4B_1 U3299 (.X(n1251), 
	.B3(n434), 
	.B2(n555), 
	.B1(n556), 
	.A(n1357));
   SEN_INV_S_3 U3300 (.X(n1122), 
	.A(n1121));
   SEN_ND2_4 U3301 (.X(n1171), 
	.A2(n1144), 
	.A1(n813));
   SEN_ND2_4 U3302 (.X(n1438), 
	.A2(n1207), 
	.A1(n1206));
   SEN_INV_S_4 U3303 (.X(n1219), 
	.A(pprow5_qual[5]));
   SEN_AOI311_4 U3304 (.X(n1222), 
	.B2(n1220), 
	.B1(n1221), 
	.A3(n1311), 
	.A2(n552), 
	.A1(n703));
   SEN_NR2B_4 U3305 (.X(n1391), 
	.B(net83111), 
	.A(n1390));
   SEN_OAI221_4 U3306 (.X(n1773), 
	.C(n1770), 
	.B2(net82284), 
	.B1(net95872), 
	.A2(net82284), 
	.A1(n1771));
   SEN_EO2_2 U274 (.X(net82119), 
	.A2(net82124), 
	.A1(net82123));
   SEN_EO2_S_0P5 U1696 (.X(net82122), 
	.A2(pprow1_qual[29]), 
	.A1(pprow0_qual[31]));
   SEN_ND2_S_0P5 U1259 (.X(net91410), 
	.A2(net91386), 
	.A1(net91394));
   SEN_INV_S_1 U1257 (.X(net91394), 
	.A(pprow1_qual[27]));
   SEN_EN2_5 U1695 (.X(net82120), 
	.A2(net91394), 
	.A1(net82122));
   SEN_EO3_4 U1694 (.X(net82115), 
	.A3(C[31]), 
	.A2(net82120), 
	.A1(net82119));
   SEN_EN2_0P5 U1693 (.X(n175), 
	.A2(pprow11_qual[7]), 
	.A1(pprow10_qual[9]));
   SEN_EO2_S_0P5 U1692 (.X(net82116), 
	.A2(n175), 
	.A1(pprow12_qual[5]));
   SEN_EO3_4 U1691 (.X(n177), 
	.A3(net82116), 
	.A2(net82115), 
	.A1(net82114));
   SEN_EN2_0P5 U1690 (.X(n174), 
	.A2(pprow5_qual[19]), 
	.A1(pprow4_qual[21]));
   SEN_EO2_S_0P5 U1689 (.X(n171), 
	.A2(n174), 
	.A1(pprow6_qual[17]));
   SEN_AN2_S_1 U1688 (.X(n176), 
	.A2(pprow14_qual[0]), 
	.A1(\bmul/neg15 ));
   SEN_EO3_1 U1687 (.X(n172), 
	.A3(pprow3_qual[23]), 
	.A2(pprow2_qual[25]), 
	.A1(n176));
   SEN_EO2_DG_8 U1686 (.X(n178), 
	.A2(n172), 
	.A1(n171));
   SEN_EN3_6 U360 (.X(n163), 
	.A3(n178), 
	.A2(n177), 
	.A1(n46));
   SEN_ND2_T_6 U1685 (.X(n170), 
	.A2(net82102), 
	.A1(net85897));
   SEN_OA2BB2_8 U1684 (.X(net82087), 
	.B2(net85897), 
	.B1(net82102), 
	.A2(n170), 
	.A1(net82100));
   SEN_INV_S_1 U1683 (.X(n167), 
	.A(pprow2_qual[24]));
   SEN_INV_S_1 U1682 (.X(n168), 
	.A(pprow3_qual[22]));
   SEN_ND2_G_1 U1681 (.X(n169), 
	.A2(pprow3_qual[22]), 
	.A1(pprow2_qual[24]));
   SEN_AOAI211_6 U1680 (.X(n164), 
	.C(n169), 
	.B(net82098), 
	.A2(n168), 
	.A1(n167));
   SEN_OR2_1 U1679 (.X(n173), 
	.A2(pprow5_qual[18]), 
	.A1(pprow4_qual[20]));
   SEN_INV_S_1 U2076 (.X(net90456), 
	.A(pprow4_qual[20]));
   SEN_EN2_DG_8 U158 (.X(n31), 
	.A2(net90456), 
	.A1(n166));
   SEN_INV_S_1 U1678 (.X(n166), 
	.A(pprow5_qual[18]));
   SEN_OA2BB2_8 U1677 (.X(n165), 
	.B2(n166), 
	.B1(net90456), 
	.A2(n173), 
	.A1(net82091));
   SEN_EO2_5 U30 (.X(net82088), 
	.A2(n165), 
	.A1(n164));
   SEN_EO3_4 U1140 (.X(net82085), 
	.A3(net82088), 
	.A2(net82087), 
	.A1(n163));
   SEN_EN3_6 U1676 (.X(net82073), 
	.A3(net82085), 
	.A2(net82084), 
	.A1(net82083));
   SEN_EO2_S_6 U1097 (.X(net82072), 
	.A2(net82073), 
	.A1(net82074));
   SEN_ND2_T_2 U455 (.X(net87948), 
	.A2(net87947), 
	.A1(net82064));
   SEN_INV_6 U460 (.X(net87946), 
	.A(net82064));
   SEN_EO2_S_6 U456 (.X(net82064), 
	.A2(net82072), 
	.A1(net82071));
   SEN_FDPQ_D_3 \pprow0_qual_reg[2]  (.Q(pprow0_qual[2]), 
	.D(pprow0[2]), 
	.CK(CLK));
   SEN_FDPQ_4 \pprow2_qual_reg[11]  (.Q(pprow2_qual[11]), 
	.D(pprow2[11]), 
	.CK(CLK));
   SEN_INV_6 U21 (.X(net83636), 
	.A(net83632));
   SEN_EN2_6 U22 (.X(net83632), 
	.A2(n2037), 
	.A1(n2036));
   SEN_INV_32 U32 (.X(n2036), 
	.A(n396));
   SEN_AO21B_6 U34 (.X(n2037), 
	.B(net101269), 
	.A2(net82999), 
	.A1(n565));
   SEN_INV_2P5 U36 (.X(n290), 
	.A(C[2]));
   SEN_INV_4 U37 (.X(n297), 
	.A(net83861));
   SEN_EO2_2 U40 (.X(n887), 
	.A2(net84371), 
	.A1(net84370));
   SEN_AO2BB2_8 U49 (.X(n895), 
	.B2(n886), 
	.B1(n887), 
	.A2(n889), 
	.A1(n890));
   SEN_INV_10 U51 (.X(n62), 
	.A(n63));
   SEN_BUF_S_1 U60 (.X(n2038), 
	.A(net83392));
   SEN_ND2_G_3 U66 (.X(net83392), 
	.A2(net83424), 
	.A1(n56));
   SEN_ND2_T_3 U67 (.X(net83174), 
	.A2(net83392), 
	.A1(n1268));
   SEN_ND2B_V1_3 U70 (.X(net83777), 
	.B(n185), 
	.A(net83573));
   SEN_INV_S_4 U72 (.X(net83380), 
	.A(net83381));
   SEN_AOI31_8 U75 (.X(n446), 
	.B(n448), 
	.A3(n249), 
	.A2(n447), 
	.A1(net84322));
   SEN_INV_3 U92 (.X(n398), 
	.A(net87796));
   SEN_NR2_T_6 U94 (.X(net83000), 
	.A2(net86560), 
	.A1(net83523));
   SEN_ND2_6 U96 (.X(n55), 
	.A2(n54), 
	.A1(n57));
   SEN_ND2_T_2 U102 (.X(n1269), 
	.A2(net83852), 
	.A1(net83851));
   SEN_BUF_2 U106 (.X(n301), 
	.A(net83851));
   SEN_AN2_6 U111 (.X(n2039), 
	.A2(n1452), 
	.A1(n1451));
   SEN_ND2_T_2 U121 (.X(n1630), 
	.A2(n1537), 
	.A1(n1536));
   SEN_BUF_1 U122 (.X(n2040), 
	.A(net82846));
   SEN_EO2_S_1 U131 (.X(n1537), 
	.A2(n736), 
	.A1(n1590));
   SEN_EO2_DG_1 U139 (.X(n656), 
	.A2(n1327), 
	.A1(n1449));
   SEN_AOI21_T_2 U152 (.X(net90917), 
	.B(n331), 
	.A2(n330), 
	.A1(n329));
   SEN_ND2B_V1DG_4 U155 (.X(net84193), 
	.B(n898), 
	.A(n901));
   SEN_AOI21_2 U166 (.X(n1586), 
	.B(n1579), 
	.A2(n1580), 
	.A1(n1581));
   SEN_INV_6 U169 (.X(n1449), 
	.A(n1328));
   SEN_INV_6 U170 (.X(n85), 
	.A(n83));
   SEN_EO2_3 U173 (.X(n1724), 
	.A2(n711), 
	.A1(n1718));
   SEN_INV_S_3 U174 (.X(net83373), 
	.A(net83374));
   SEN_NR3_T_5 U179 (.X(n2065), 
	.A3(n2067), 
	.A2(n2063), 
	.A1(n2066));
   SEN_INV_2 U185 (.X(n1073), 
	.A(n1065));
   SEN_AO21B_8 U192 (.X(n1722), 
	.B(n1678), 
	.A2(n1679), 
	.A1(n1680));
   SEN_INV_2 U196 (.X(net82616), 
	.A(n161));
   SEN_EO3_6 U199 (.X(n46), 
	.A3(n183), 
	.A2(n2041), 
	.A1(net82142));
   SEN_AOI22_T_6 U203 (.X(n2041), 
	.B2(pprow8_qual[12]), 
	.B1(pprow9_qual[10]), 
	.A2(n118), 
	.A1(n1816));
   SEN_BUF_1 U208 (.X(n2042), 
	.A(net94132));
   SEN_INV_8 U210 (.X(net94132), 
	.A(net85071));
   SEN_NR2_T_8 U220 (.X(n1261), 
	.A2(n1259), 
	.A1(n581));
   SEN_INV_S_0P5 U221 (.X(n2043), 
	.A(n199));
   SEN_ND2_T_4 U228 (.X(n199), 
	.A2(net83875), 
	.A1(n190));
   SEN_INV_6 U231 (.X(net95536), 
	.A(net94217));
   SEN_AN2_2 U232 (.X(n547), 
	.A2(n1724), 
	.A1(n1723));
   SEN_INV_AS_10 U235 (.X(n482), 
	.A(n486));
   SEN_ND2_G_1 U238 (.X(n53), 
	.A2(pprow0_qual[11]), 
	.A1(C[11]));
   SEN_INV_3 U242 (.X(net86560), 
	.A(net86559));
   SEN_EO2_8 U243 (.X(n1123), 
	.A2(n1099), 
	.A1(n1100));
   SEN_ND2B_3 U255 (.X(n889), 
	.B(n875), 
	.A(n874));
   SEN_BUF_AS_3 U263 (.X(n602), 
	.A(n1564));
   SEN_NR2_G_3 U280 (.X(n1564), 
	.A2(net82717), 
	.A1(n1561));
   SEN_INV_2P5 U283 (.X(net82970), 
	.A(net82965));
   SEN_BUF_6 U287 (.X(n552), 
	.A(n1306));
   SEN_ND2_S_8 U301 (.X(n1711), 
	.A2(n1659), 
	.A1(n645));
   SEN_EO2_G_4 U317 (.X(n1484), 
	.A2(n515), 
	.A1(n723));
   SEN_EO2_DG_1 U319 (.X(n1405), 
	.A2(n1401), 
	.A1(n720));
   SEN_INV_8 U324 (.X(n71), 
	.A(net90814));
   SEN_EN2_3 U331 (.X(net83634), 
	.A2(net83743), 
	.A1(n82));
   SEN_INV_6 U332 (.X(net83740), 
	.A(net83741));
   SEN_ND2_T_16 U333 (.X(net83741), 
	.A2(net83648), 
	.A1(net83647));
   SEN_ND2B_8 U335 (.X(net84152), 
	.B(n944), 
	.A(C[9]));
   SEN_ND2_T_2 U339 (.X(n1443), 
	.A2(n1327), 
	.A1(n1449));
   SEN_INV_AS_10 U340 (.X(n314), 
	.A(net83415));
   SEN_NR2_T_6 U342 (.X(net84238), 
	.A2(net84241), 
	.A1(n435));
   SEN_BUF_S_2 U345 (.X(n2044), 
	.A(net82967));
   SEN_ND2_8 U352 (.X(net82967), 
	.A2(n314), 
	.A1(n313));
   SEN_AN3B_4 U361 (.X(n1433), 
	.B2(n1428), 
	.B1(n1429), 
	.A(n1427));
   SEN_ND2_G_1 U362 (.X(n1594), 
	.A2(net82741), 
	.A1(n1549));
   SEN_EO2_S_0P5 U366 (.X(n1496), 
	.A2(n1549), 
	.A1(net82741));
   SEN_EO2_4 U373 (.X(n1549), 
	.A2(n1494), 
	.A1(n1495));
   SEN_ND2_S_2 U381 (.X(n1037), 
	.A2(n512), 
	.A1(n30));
   SEN_EO2_2 U385 (.X(net86454), 
	.A2(net82582), 
	.A1(net82581));
   SEN_AOAI211_3 U391 (.X(n1370), 
	.C(n1329), 
	.B(n1330), 
	.A2(n1331), 
	.A1(n1332));
   SEN_EO2_S_1 U403 (.X(n1487), 
	.A2(n1480), 
	.A1(n1523));
   SEN_NR2_G_4 U408 (.X(n1134), 
	.A2(net83786), 
	.A1(net83787));
   SEN_NR2_T_5 U420 (.X(n477), 
	.A2(n475), 
	.A1(n378));
   SEN_AN2_S_8 U423 (.X(n2045), 
	.A2(n1096), 
	.A1(n1097));
   SEN_INV_S_6 U427 (.X(n1096), 
	.A(n1095));
   SEN_INV_3 U430 (.X(n200), 
	.A(net84063));
   SEN_EO2_1 U438 (.X(n696), 
	.A2(n1723), 
	.A1(n1724));
   SEN_INV_4 U440 (.X(net95928), 
	.A(net84028));
   SEN_ND2_G_4 U481 (.X(net84028), 
	.A2(net83741), 
	.A1(net84029));
   SEN_BUF_S_4 U527 (.X(n436), 
	.A(n42));
   SEN_ND2_0P8 U529 (.X(n483), 
	.A2(net83301), 
	.A1(net83555));
   SEN_ND2_2 U532 (.X(n1265), 
	.A2(n1438), 
	.A1(n1264));
   SEN_BUF_S_6 U533 (.X(n300), 
	.A(n293));
   SEN_INV_10 U534 (.X(net82999), 
	.A(net83830));
   SEN_NR2B_V1_2 U537 (.X(n954), 
	.B(net84057), 
	.A(net84208));
   SEN_ND2_T_1 U539 (.X(n953), 
	.A2(net84058), 
	.A1(n438));
   SEN_EO2_6 U540 (.X(n2101), 
	.A2(n2065), 
	.A1(n2079));
   SEN_AN2_1P5 U545 (.X(n626), 
	.A2(n1175), 
	.A1(n1176));
   SEN_OR2_2 U564 (.X(n1176), 
	.A2(pprow5_qual[2]), 
	.A1(pprow4_qual[4]));
   SEN_EN2_S_3 U565 (.X(net83462), 
	.A2(n1222), 
	.A1(n122));
   SEN_INV_5 U568 (.X(n237), 
	.A(n300));
   SEN_INV_S_8 U596 (.X(net84734), 
	.A(n288));
   SEN_INV_0P65 U601 (.X(n238), 
	.A(net84393));
   SEN_ND2_2 U608 (.X(n278), 
	.A2(n281), 
	.A1(net84392));
   SEN_ND2_T_1P5 U613 (.X(n582), 
	.A2(net84471), 
	.A1(net88056));
   SEN_NR2B_V1_8 U616 (.X(n487), 
	.B(net83546), 
	.A(net83544));
   SEN_ND2_6 U624 (.X(net83546), 
	.A2(n1183), 
	.A1(net83685));
   SEN_NR2_S_1 U627 (.X(net83885), 
	.A2(net83782), 
	.A1(n1132));
   SEN_INV_1P25 U629 (.X(n2046), 
	.A(net88108));
   SEN_AN2_4 U637 (.X(net88108), 
	.A2(n482), 
	.A1(net83550));
   SEN_ND2_G_1 U638 (.X(n926), 
	.A2(pprow1_qual[1]), 
	.A1(pprow1_qual[3]));
   SEN_ND2_2 U644 (.X(n1001), 
	.A2(pprow1_qual[3]), 
	.A1(pprow1_qual[5]));
   SEN_ND2_3 U646 (.X(n906), 
	.A2(n904), 
	.A1(n942));
   SEN_OAI21_G_2 U647 (.X(n972), 
	.B(n962), 
	.A2(n963), 
	.A1(n964));
   SEN_ND2_8 U652 (.X(net83584), 
	.A2(net83962), 
	.A1(net83961));
   SEN_INV_6 U664 (.X(net84650), 
	.A(n201));
   SEN_NR2_T_6 U681 (.X(n1054), 
	.A2(n1053), 
	.A1(n617));
   SEN_INV_S_6 U686 (.X(n313), 
	.A(net83414));
   SEN_ND2_T_2 U689 (.X(net82998), 
	.A2(net82999), 
	.A1(net83000));
   SEN_OAI21B_8 U691 (.X(n1600), 
	.B(n21), 
	.A2(n1546), 
	.A1(n1545));
   SEN_ND2_T_6 U701 (.X(n1545), 
	.A2(n184), 
	.A1(n559));
   SEN_BUF_1 U707 (.X(n2047), 
	.A(net85837));
   SEN_EO2_2 U710 (.X(net85837), 
	.A2(net85838), 
	.A1(n238));
   SEN_AOAI211_8 U712 (.X(n1373), 
	.C(n1335), 
	.B(n1336), 
	.A2(n1337), 
	.A1(n1338));
   SEN_EN2_5 U716 (.X(net82717), 
	.A2(net82721), 
	.A1(n160));
   SEN_EO2_1 U722 (.X(net83018), 
	.A2(n1461), 
	.A1(n1462));
   SEN_ND2_G_3 U741 (.X(n536), 
	.A2(n1462), 
	.A1(n1461));
   SEN_INV_2 U742 (.X(n1580), 
	.A(n1462));
   SEN_ND2_T_8 U743 (.X(net94217), 
	.A2(net83169), 
	.A1(net95509));
   SEN_AN2_6 U755 (.X(n435), 
	.A2(n392), 
	.A1(net84730));
   SEN_ND2_T_2 U756 (.X(n2048), 
	.A2(net83549), 
	.A1(n243));
   SEN_ND2_6 U757 (.X(net83302), 
	.A2(net83549), 
	.A1(n243));
   SEN_INV_S_0P5 U766 (.X(net95817), 
	.A(n315));
   SEN_BUF_1 U769 (.X(n2049), 
	.A(n1208));
   SEN_OAI21_5 U773 (.X(net83833), 
	.B(net84355), 
	.A2(net84354), 
	.A1(net84391));
   SEN_EN2_5 U777 (.X(net84187), 
	.A2(net84111), 
	.A1(net86002));
   SEN_ND2_T_2 U785 (.X(n1471), 
	.A2(n1500), 
	.A1(n1505));
   SEN_NR2_S_5 U790 (.X(net95509), 
	.A2(net85071), 
	.A1(net83168));
   SEN_NR3_T_6 U796 (.X(net87627), 
	.A3(n440), 
	.A2(n441), 
	.A1(net95536));
   SEN_OAI21_T_4 U798 (.X(net83165), 
	.B(n55), 
	.A2(net83389), 
	.A1(net83390));
   SEN_ND2_T_5 U801 (.X(net83166), 
	.A2(net83390), 
	.A1(net83389));
   SEN_EN2_S_4 U804 (.X(net83390), 
	.A2(net83437), 
	.A1(net83436));
   SEN_BUF_S_6 U811 (.X(net85046), 
	.A(net83387));
   SEN_NR2_S_2 U815 (.X(n273), 
	.A2(net87846), 
	.A1(net84471));
   SEN_ND2_2 U825 (.X(net87846), 
	.A2(n289), 
	.A1(pprow0_qual[0]));
   SEN_ND2_S_6 U829 (.X(n507), 
	.A2(n30), 
	.A1(n512));
   SEN_INV_2 U830 (.X(n2050), 
	.A(n1228));
   SEN_INV_S_3 U833 (.X(n2051), 
	.A(n2050));
   SEN_EO2_2 U847 (.X(n1228), 
	.A2(n716), 
	.A1(n1235));
   SEN_INV_2 U853 (.X(net84415), 
	.A(net84384));
   SEN_EO2_3 U858 (.X(n880), 
	.A2(net84408), 
	.A1(net84407));
   SEN_ND2_T_2 U863 (.X(net83887), 
	.A2(net83962), 
	.A1(net83961));
   SEN_ND2_4 U871 (.X(net84056), 
	.A2(net84248), 
	.A1(net83961));
   SEN_ND2B_V1_4 U873 (.X(net83851), 
	.B(n990), 
	.A(n992));
   SEN_INV_2 U897 (.X(n990), 
	.A(n991));
   SEN_EO2_S_0P5 U908 (.X(n686), 
	.A2(n991), 
	.A1(n992));
   SEN_ND2_4 U921 (.X(net84042), 
	.A2(n991), 
	.A1(n992));
   SEN_EO2_4 U924 (.X(n991), 
	.A2(n973), 
	.A1(n974));
   SEN_EO2_S_6 U940 (.X(n1452), 
	.A2(n1261), 
	.A1(n1262));
   SEN_NR2_2 U941 (.X(n1259), 
	.A2(n1268), 
	.A1(net83422));
   SEN_INV_4 U945 (.X(net84235), 
	.A(net84236));
   SEN_ND2_6 U948 (.X(net84283), 
	.A2(net84236), 
	.A1(net84227));
   SEN_ND2_G_6 U950 (.X(net84236), 
	.A2(net84159), 
	.A1(net84358));
   SEN_ND2_6 U953 (.X(n1235), 
	.A2(n1216), 
	.A1(n1217));
   SEN_ND2_3 U956 (.X(n640), 
	.A2(net87769), 
	.A1(n638));
   SEN_ND2B_V1DG_8 U986 (.X(n1505), 
	.B(n1469), 
	.A(n767));
   SEN_INV_10 U992 (.X(n1338), 
	.A(n1333));
   SEN_EO2_DG_1 U1005 (.X(net83334), 
	.A2(n1238), 
	.A1(n1300));
   SEN_ND2_6 U1016 (.X(net83158), 
	.A2(net83163), 
	.A1(net83164));
   SEN_INV_5 U1023 (.X(net83171), 
	.A(net95543));
   SEN_EO2_DG_1 U1035 (.X(net82582), 
	.A2(n691), 
	.A1(n1612));
   SEN_INV_AS_10 U1045 (.X(n64), 
	.A(net82937));
   SEN_EN2_S_4 U1050 (.X(net86459), 
	.A2(n2053), 
	.A1(net82939));
   SEN_ND2_T_3 U1061 (.X(n1456), 
	.A2(n642), 
	.A1(n641));
   SEN_ND2_G_3 U1064 (.X(net82332), 
	.A2(n1771), 
	.A1(net82058));
   SEN_ND2_T_3 U1079 (.X(n1771), 
	.A2(net82333), 
	.A1(net82334));
   SEN_BUF_4 U1110 (.X(net101261), 
	.A(net82936));
   SEN_ND2_T_2 U1135 (.X(n976), 
	.A2(net84115), 
	.A1(net86698));
   SEN_ND3_8 U1148 (.X(n781), 
	.A3(n705), 
	.A2(n1522), 
	.A1(n1521));
   SEN_ND2B_6 U1174 (.X(n1521), 
	.B(n1519), 
	.A(n1520));
   SEN_OAI21_5 U1187 (.X(net83293), 
	.B(net83299), 
	.A2(net83298), 
	.A1(n25));
   SEN_INV_S_6 U1196 (.X(net83298), 
	.A(net83300));
   SEN_AOI22_T_6 U1199 (.X(n1341), 
	.B2(n1297), 
	.B1(n1298), 
	.A2(n1299), 
	.A1(n1300));
   SEN_INV_S_4 U1217 (.X(n1563), 
	.A(n1560));
   SEN_OAOI211_8 U1221 (.X(n1409), 
	.C(n1375), 
	.B(n1376), 
	.A2(n1377), 
	.A1(n1378));
   SEN_ND2_G_4 U1222 (.X(n1437), 
	.A2(n1208), 
	.A1(n1209));
   SEN_ND2_T_4 U1230 (.X(n1118), 
	.A2(n394), 
	.A1(net83507));
   SEN_OAOI211_G_8 U1252 (.X(net83452), 
	.C(n471), 
	.B(net83453), 
	.A2(net83455), 
	.A1(n478));
   SEN_INV_2 U1264 (.X(n89), 
	.A(n88));
   SEN_NR2_6 U1294 (.X(n565), 
	.A2(net90705), 
	.A1(net83740));
   SEN_NR2B_V1DG_8 U1365 (.X(n1446), 
	.B(net82962), 
	.A(n1439));
   SEN_INV_1 U1424 (.X(net84192), 
	.A(net84276));
   SEN_ND2_S_3 U1431 (.X(n1598), 
	.A2(n1597), 
	.A1(n1596));
   SEN_AO21B_2 U1440 (.X(n745), 
	.B(n1337), 
	.A2(n1334), 
	.A1(n1333));
   SEN_EO2_2 U1441 (.X(n1339), 
	.A2(n745), 
	.A1(n744));
   SEN_INV_10 U1445 (.X(net82335), 
	.A(net82333));
   SEN_ND2_T_8 U1456 (.X(net82333), 
	.A2(\bmul/neg14 ), 
	.A1(n1760));
   SEN_EO2_8 U1482 (.X(n1760), 
	.A2(n103), 
	.A1(n1759));
   SEN_OAI21B_4 U1495 (.X(n2052), 
	.B(n21), 
	.A2(n1546), 
	.A1(n1545));
   SEN_INV_S_4 U1539 (.X(n1659), 
	.A(n18));
   SEN_ND2_G_1 U1549 (.X(n1279), 
	.A2(pprow1_qual[14]), 
	.A1(pprow1_qual[16]));
   SEN_NR2_S_2 U1552 (.X(n1277), 
	.A2(n1271), 
	.A1(n94));
   SEN_ND3_2 U1575 (.X(n1271), 
	.A3(n1270), 
	.A2(n1278), 
	.A1(n1279));
   SEN_ND2_4 U1587 (.X(n959), 
	.A2(net84223), 
	.A1(n946));
   SEN_EN2_3 U1596 (.X(n946), 
	.A2(n930), 
	.A1(n727));
   SEN_NR2_T_5 U1605 (.X(n930), 
	.A2(n570), 
	.A1(net84281));
   SEN_EN2_S_2 U1612 (.X(n875), 
	.A2(n873), 
	.A1(net84405));
   SEN_NR2_G_4 U1614 (.X(n890), 
	.A2(n886), 
	.A1(n887));
   SEN_INV_4 U1615 (.X(n1324), 
	.A(n1452));
   SEN_AOAI211_8 U1620 (.X(net82857), 
	.C(n61), 
	.B(net82936), 
	.A2(n60), 
	.A1(n2053));
   SEN_ND2_8 U1657 (.X(net84002), 
	.A2(net84202), 
	.A1(net84201));
   SEN_NR2_T_5 U1705 (.X(n1057), 
	.A2(net88108), 
	.A1(n572));
   SEN_EO2_S_6 U1708 (.X(n1448), 
	.A2(net83452), 
	.A1(net83451));
   SEN_NR2_T_8 U1709 (.X(n1702), 
	.A2(n549), 
	.A1(n1698));
   SEN_INV_S_4 U1716 (.X(net87798), 
	.A(n186));
   SEN_INV_0P8 U1720 (.X(n567), 
	.A(net83634));
   SEN_ND2_T_5 U1721 (.X(n2053), 
	.A2(n66), 
	.A1(n65));
   SEN_ND2_12 U1723 (.X(n63), 
	.A2(n66), 
	.A1(n65));
   SEN_ND2B_V1_4 U1733 (.X(net84003), 
	.B(net84007), 
	.A(net84009));
   SEN_ND3_T_2 U1734 (.X(net83374), 
	.A3(n1106), 
	.A2(n1105), 
	.A1(n1104));
   SEN_ND2_S_4 U1736 (.X(n1444), 
	.A2(n1448), 
	.A1(n1324));
   SEN_EO2_4 U1738 (.X(net90868), 
	.A2(n930), 
	.A1(n727));
   SEN_NR2_T_8 U1741 (.X(net82836), 
	.A2(n302), 
	.A1(net86483));
   SEN_EO2_2 U1743 (.X(n1169), 
	.A2(n1167), 
	.A1(n1168));
   SEN_ND3_T_2 U1746 (.X(n2054), 
	.A3(n304), 
	.A2(net84186), 
	.A1(n303));
   SEN_NR3_T_6 U1747 (.X(n591), 
	.A3(net97222), 
	.A2(net90258), 
	.A1(net87990));
   SEN_INV_6 U1760 (.X(net84322), 
	.A(net84283));
   SEN_ND2_T_4 U1765 (.X(n1613), 
	.A2(n1611), 
	.A1(n1612));
   SEN_ND2_T_0P5 U1768 (.X(n393), 
	.A2(net82430), 
	.A1(net88080));
   SEN_ND2_G_4 U1769 (.X(n304), 
	.A2(n305), 
	.A1(n309));
   SEN_INV_4 U1777 (.X(n305), 
	.A(net84372));
   SEN_ND3_6 U1779 (.X(net83861), 
	.A3(n304), 
	.A2(net84186), 
	.A1(n303));
   SEN_INV_5 U1786 (.X(net88014), 
	.A(net82310));
   SEN_ND2_T_2 U1789 (.X(net87837), 
	.A2(net86446), 
	.A1(net82436));
   SEN_INV_3 U1791 (.X(n379), 
	.A(n378));
   SEN_INV_3 U1802 (.X(n378), 
	.A(n470));
   SEN_AN4B_4 U1803 (.X(n423), 
	.B3(net83565), 
	.B2(net83566), 
	.B1(net83584), 
	.A(net83585));
   SEN_ND2_2 U1834 (.X(n214), 
	.A2(net83114), 
	.A1(n232));
   SEN_ND2_S_4 U1837 (.X(n231), 
	.A2(n137), 
	.A1(n232));
   SEN_ND3_T_4 U1844 (.X(net83585), 
	.A3(net83781), 
	.A2(n1133), 
	.A1(net83577));
   SEN_ND2_T_2 U1846 (.X(n648), 
	.A2(net83299), 
	.A1(net83308));
   SEN_INV_3 U1876 (.X(n1779), 
	.A(n1775));
   SEN_INV_4 U1900 (.X(net84156), 
	.A(net84152));
   SEN_INV_3 U1909 (.X(n1206), 
	.A(n1210));
   SEN_EO2_6 U1967 (.X(net82522), 
	.A2(n643), 
	.A1(n2055));
   SEN_EN2_DG_8 U1988 (.X(n2055), 
	.A2(n661), 
	.A1(n1660));
   SEN_ND2B_V1_6 U2050 (.X(net83301), 
	.B(net83684), 
	.A(net83678));
   SEN_AN2_1 U2058 (.X(n572), 
	.A2(net83552), 
	.A1(n1056));
   SEN_ND2_4 U2063 (.X(n474), 
	.A2(net94064), 
	.A1(n477));
   SEN_INV_2P5 U2065 (.X(n1450), 
	.A(n1448));
   SEN_INV_S_4 U2069 (.X(net87836), 
	.A(net82436));
   SEN_OAOI211_8 U2099 (.X(n520), 
	.C(n1589), 
	.B(n1590), 
	.A2(pprow10_qual[3]), 
	.A1(pprow11_qual[1]));
   SEN_EO2_2 U2101 (.X(n1488), 
	.A2(net82768), 
	.A1(n86));
   SEN_ND2_T_5 U2161 (.X(net82309), 
	.A2(net82428), 
	.A1(net82429));
   SEN_EN2_6 U2184 (.X(net83096), 
	.A2(n519), 
	.A1(n684));
   SEN_AOI21B_4 U2217 (.X(n519), 
	.B(net83127), 
	.A2(n1347), 
	.A1(n1348));
   SEN_EO2_S_3 U2246 (.X(n512), 
	.A2(net84066), 
	.A1(net85880));
   SEN_ND3_T_1 U2255 (.X(n1430), 
	.A3(n1365), 
	.A2(n1366), 
	.A1(n1367));
   SEN_EN2_5 U2260 (.X(net91120), 
	.A2(net83156), 
	.A1(n2056));
   SEN_EO2_DG_8 U2266 (.X(n2056), 
	.A2(net95557), 
	.A1(net83077));
   SEN_INV_AS_10 U2282 (.X(net82962), 
	.A(net82967));
   SEN_OA21_4 U2288 (.X(n41), 
	.B(n2044), 
	.A2(n312), 
	.A1(n311));
   SEN_MUX2_6 U2303 (.X(n83), 
	.S(n272), 
	.D1(n279), 
	.D0(n278));
   SEN_EN2_S_4 U2305 (.X(n513), 
	.A2(net84059), 
	.A1(net84058));
   SEN_INV_1 U2381 (.X(net84059), 
	.A(net84057));
   SEN_ND2B_4 U2396 (.X(net83332), 
	.B(net83614), 
	.A(net83611));
   SEN_ND2_T_4 U2426 (.X(n475), 
	.A2(n472), 
	.A1(n327));
   SEN_ND2_1P5 U2546 (.X(n1629), 
	.A2(n1627), 
	.A1(n1628));
   SEN_EO2_0P5 U3210 (.X(n683), 
	.A2(n1628), 
	.A1(n1627));
   SEN_EN2_S_4 U3229 (.X(net82114), 
	.A2(n179), 
	.A1(n43));
   SEN_NR3_T_6 U3235 (.X(n2057), 
	.A3(n2060), 
	.A2(n2059), 
	.A1(n2058));
   SEN_INV_S_4 U3243 (.X(n2061), 
	.A(pprow5_qual[13]));
   SEN_INV_S_4 U3307 (.X(n2062), 
	.A(pprow4_qual[15]));
   SEN_ND2B_4 U3308 (.X(n2068), 
	.B(n2069), 
	.A(n2062));
   SEN_ND2B_4 U3309 (.X(n2064), 
	.B(n2069), 
	.A(n2061));
   SEN_ND2_4 U3310 (.X(n2070), 
	.A2(pprow4_qual[16]), 
	.A1(pprow5_qual[14]));
   SEN_NR2_T_4 U3311 (.X(n2071), 
	.A2(n2070), 
	.A1(n2072));
   SEN_ND2B_4 U3312 (.X(n2073), 
	.B(n2074), 
	.A(n2072));
   SEN_ND2_4 U3313 (.X(n2075), 
	.A2(pprow4_qual[15]), 
	.A1(pprow5_qual[13]));
   SEN_NR2_T_4 U3314 (.X(n2076), 
	.A2(n2075), 
	.A1(n2077));
   SEN_NR2_T_4 U3315 (.X(n2078), 
	.A2(n2075), 
	.A1(n2073));
   SEN_EO2_6 U3316 (.X(n747), 
	.A2(pprow4_qual[14]), 
	.A1(pprow5_qual[12]));
   SEN_NR2B_4 U3317 (.X(n2080), 
	.B(n2077), 
	.A(n2081));
   SEN_NR2B_4 U3318 (.X(n2082), 
	.B(n2077), 
	.A(n2083));
   SEN_NR2B_4 U3319 (.X(n2089), 
	.B(n2064), 
	.A(n2090));
   SEN_NR2B_4 U3320 (.X(n2091), 
	.B(n2068), 
	.A(n2090));
   SEN_ND2_4 U3321 (.X(n2092), 
	.A2(n2094), 
	.A1(n2093));
   SEN_ND2_4 U3322 (.X(n2097), 
	.A2(n2095), 
	.A1(n2096));
   SEN_INV_S_4 U3323 (.X(n1727), 
	.A(n2097));
   SEN_INV_S_4 U3324 (.X(n2094), 
	.A(n1669));
   SEN_OR2_5 U3325 (.X(n2069), 
	.A2(pprow4_qual[14]), 
	.A1(pprow5_qual[12]));
   SEN_INV_S_4 U3326 (.X(n2059), 
	.A(n2069));
   SEN_OR2_5 U3327 (.X(n2085), 
	.A2(pprow5_qual[12]), 
	.A1(n1517));
   SEN_INV_S_4 U3328 (.X(n2058), 
	.A(n2085));
   SEN_OR2_5 U3329 (.X(n2074), 
	.A2(pprow5_qual[14]), 
	.A1(pprow4_qual[16]));
   SEN_INV_S_4 U3330 (.X(n2077), 
	.A(n2074));
   SEN_INV_S_4 U3331 (.X(n2087), 
	.A(n2070));
   SEN_ND2_4 U3332 (.X(n2098), 
	.A2(n2084), 
	.A1(n2088));
   SEN_INV_S_4 U3333 (.X(n588), 
	.A(n2098));
   SEN_OR2_5 U3334 (.X(n2099), 
	.A2(pprow4_qual[17]), 
	.A1(pprow5_qual[15]));
   SEN_INV_S_4 U3335 (.X(n2072), 
	.A(n2099));
   SEN_INV_S_4 U3336 (.X(n2067), 
	.A(n2075));
   SEN_INV_S_4 U3337 (.X(n2083), 
	.A(n2068));
   SEN_INV_S_4 U3338 (.X(n2081), 
	.A(n2064));
   SEN_INV_S_4 U3339 (.X(n2093), 
	.A(n2071));
   SEN_INV_S_4 U3340 (.X(n2090), 
	.A(n2073));
   SEN_EN2_5 U3341 (.X(n2079), 
	.A2(pprow4_qual[16]), 
	.A1(pprow5_qual[14]));
   SEN_EN2_5 U3342 (.X(n2100), 
	.A2(pprow4_qual[15]), 
	.A1(pprow5_qual[13]));
   SEN_EN2_S_4 U3343 (.X(n1573), 
	.A2(n2057), 
	.A1(n2100));
   SEN_EO2_2 U3344 (.X(n1623), 
	.A2(n2065), 
	.A1(n2079));
   SEN_OR2_10 U3345 (.X(n2086), 
	.A2(pprow4_qual[14]), 
	.A1(n1517));
   SEN_BUF_1 U3346 (.X(n256), 
	.A(n1517));
   SEN_NR3_G_4 U3347 (.X(n2066), 
	.A3(n2058), 
	.A2(n2060), 
	.A1(n2068));
   SEN_NR3_T_4 U3348 (.X(n2063), 
	.A3(n2058), 
	.A2(n2060), 
	.A1(n2064));
   SEN_INV_3 U3349 (.X(n2060), 
	.A(n2086));
   SEN_AOI31_2 U3350 (.X(n2096), 
	.B(n2078), 
	.A3(n2091), 
	.A2(n2086), 
	.A1(n2085));
   SEN_AOI31_2 U3351 (.X(n2095), 
	.B(n2092), 
	.A3(n2089), 
	.A2(n2086), 
	.A1(n2085));
   SEN_AOI31_2 U3352 (.X(n2088), 
	.B(n2076), 
	.A3(n2082), 
	.A2(n2086), 
	.A1(n2085));
   SEN_AOI31_2 U3353 (.X(n2084), 
	.B(n2087), 
	.A3(n2080), 
	.A2(n2086), 
	.A1(n2085));
endmodule

