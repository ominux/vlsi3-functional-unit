.subckt minbuff  VDD GND A Y
mM0 GND 5 Y GND NMOS_VTG L=5e-08 W=2.15e-07 AD=5.2675e-14 AS=2.2575e-14
+ PD=9.2e-07 PS=6.4e-07
mM1 5 A GND GND NMOS_VTG L=5e-08 W=2.15e-07 AD=2.2575e-14 AS=5.2675e-14
+ PD=6.4e-07 PS=9.2e-07
mM2 VDD 5 Y VDD PMOS_VTG L=5e-08 W=4.4e-07 AD=1.078e-13 AS=4.62e-14 PD=1.37e-06
+ PS=1.09e-06
mM3 5 A VDD VDD PMOS_VTG L=5e-08 W=4.4e-07 AD=4.62e-14 AS=1.078e-13 PD=1.09e-06
+ PS=1.37e-06
c_4 Y 0 0.0941572f
c_8 GND 0 0.0653631f
c_12 VDD 0 0.0960324f
c_16 A 0 0.0871267f
c_21 5 0 0.204263f
cc_1 GND Y 0.0606384f
cc_2 VDD Y 0.0394141f
cc_3 5 Y 0.144025f
cc_4 A GND 0.00182271f
cc_5 5 GND 0.0781011f
cc_6 A VDD 0.0015602f
cc_7 5 VDD 0.0620091f
cc_8 5 A 0.124202f
.ends

