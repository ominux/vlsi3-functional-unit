module Alu (
	Z, 
	A, 
	B, 
	INST, 
	FLAGS);
   output [31:0] Z;
   input [31:0] A;
   input [31:0] B;
   input [3:0] INST;
   output [3:0] FLAGS;

   // Internal wires
   wire \*Logic0* ;
   wire n20;
   wire n22;
   wire n24;
   wire n26;
   wire n28;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire net3712;
   wire net3715;
   wire net3718;
   wire net3721;
   wire net3724;
   wire net3727;
   wire net3730;
   wire net3733;
   wire net3736;
   wire net3739;
   wire net3742;
   wire net3745;
   wire net3748;
   wire net3751;
   wire net3754;
   wire net3757;
   wire net15760;
   wire net15762;
   wire net15763;
   wire net15769;
   wire net15775;
   wire net15784;
   wire net15785;
   wire net15786;
   wire net15787;
   wire net15790;
   wire net15791;
   wire net15794;
   wire net15795;
   wire net15796;
   wire net15797;
   wire net15798;
   wire net15799;
   wire net15800;
   wire net15801;
   wire net15817;
   wire net15818;
   wire net15819;
   wire net15829;
   wire net15830;
   wire net15831;
   wire net15832;
   wire net15846;
   wire net15847;
   wire net15848;
   wire net15857;
   wire net15858;
   wire net15859;
   wire net15865;
   wire net15869;
   wire net15870;
   wire net15871;
   wire net15880;
   wire net15881;
   wire net15882;
   wire net15883;
   wire net15884;
   wire net15885;
   wire net15886;
   wire net15888;
   wire net15889;
   wire net15894;
   wire net15899;
   wire net15902;
   wire net15903;
   wire net15904;
   wire net15910;
   wire net15912;
   wire net15913;
   wire net15914;
   wire net15915;
   wire net15919;
   wire net15920;
   wire net15921;
   wire net15927;
   wire net15928;
   wire net15929;
   wire net15934;
   wire net15936;
   wire net15937;
   wire net15938;
   wire net15939;
   wire net15941;
   wire net15945;
   wire net15946;
   wire net15947;
   wire net15948;
   wire net15949;
   wire net15953;
   wire net15956;
   wire net15958;
   wire net15960;
   wire net15961;
   wire net15963;
   wire net15964;
   wire net15965;
   wire net15967;
   wire net15968;
   wire net15969;
   wire net15971;
   wire net15973;
   wire net15975;
   wire net15976;
   wire net15977;
   wire net15979;
   wire net15980;
   wire net15985;
   wire net15986;
   wire net15987;
   wire net15988;
   wire net15995;
   wire net15996;
   wire net15997;
   wire net16005;
   wire net16006;
   wire net16007;
   wire net16009;
   wire net16010;
   wire net16013;
   wire net16014;
   wire net16015;
   wire net16018;
   wire net16020;
   wire net16021;
   wire net16023;
   wire net16028;
   wire net16029;
   wire net16030;
   wire net16037;
   wire net16038;
   wire net16039;
   wire net16051;
   wire net16052;
   wire net16053;
   wire net16057;
   wire net16062;
   wire net16064;
   wire net16065;
   wire net16066;
   wire net16069;
   wire net16070;
   wire net16073;
   wire net16074;
   wire net16077;
   wire net16078;
   wire net16079;
   wire net16080;
   wire net16084;
   wire net16085;
   wire net16086;
   wire net16087;
   wire net16102;
   wire net16103;
   wire net16104;
   wire net16113;
   wire net16123;
   wire net16125;
   wire net16134;
   wire net16143;
   wire net16144;
   wire net16145;
   wire net16146;
   wire net16152;
   wire net16153;
   wire net16154;
   wire net16155;
   wire net16156;
   wire net16165;
   wire net16178;
   wire net16179;
   wire net16180;
   wire net16182;
   wire net16188;
   wire net16190;
   wire net16191;
   wire net16192;
   wire net16193;
   wire net16196;
   wire net16197;
   wire net16200;
   wire net16201;
   wire net16220;
   wire net16222;
   wire net16223;
   wire net16284;
   wire net16288;
   wire net16289;
   wire net16291;
   wire net16293;
   wire net16298;
   wire net16299;
   wire net16300;
   wire net16301;
   wire net16309;
   wire net16311;
   wire net16322;
   wire net16325;
   wire net16326;
   wire net16327;
   wire net16328;
   wire net16336;
   wire net16337;
   wire net16344;
   wire net16345;
   wire net16360;
   wire net16395;
   wire net16400;
   wire net16407;
   wire net16408;
   wire net16412;
   wire net16410;
   wire net16424;
   wire net16422;
   wire net16440;
   wire net16434;
   wire net16448;
   wire net16444;
   wire net16478;
   wire net16476;
   wire net16474;
   wire net16486;
   wire net16482;
   wire net16480;
   wire net16495;
   wire net16497;
   wire net16499;
   wire net16501;
   wire net16669;
   wire net16691;
   wire net16701;
   wire net16723;
   wire net16774;
   wire net16772;
   wire net16938;
   wire net16949;
   wire net16968;
   wire net16985;
   wire net16999;
   wire net17000;
   wire net17005;
   wire net17035;
   wire net17190;
   wire net17189;
   wire net17414;
   wire net17420;
   wire net17428;
   wire net17427;
   wire net17564;
   wire net17573;
   wire net17572;
   wire net17579;
   wire net17584;
   wire net17602;
   wire net17601;
   wire net17600;
   wire net17648;
   wire net17656;
   wire net17655;
   wire net17669;
   wire net17668;
   wire net17713;
   wire net17749;
   wire net17760;
   wire net17788;
   wire net17799;
   wire net17804;
   wire net17816;
   wire net17829;
   wire net17843;
   wire net18157;
   wire net18184;
   wire net18219;
   wire net18229;
   wire net18246;
   wire net16215;
   wire net16127;
   wire net17773;
   wire net17750;
   wire net17550;
   wire net16287;
   wire net16282;
   wire net16281;
   wire net15942;
   wire net15916;
   wire net15897;
   wire net17349;
   wire net16292;
   wire net15940;
   wire net16361;
   wire net16177;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire n587;
   wire n588;
   wire n589;
   wire n590;
   wire n591;
   wire n592;
   wire n593;
   wire n594;
   wire n595;
   wire n596;
   wire n597;
   wire n598;
   wire n599;
   wire n600;
   wire n601;
   wire n602;
   wire n603;
   wire n604;
   wire n605;
   wire n606;
   wire n607;
   wire n608;
   wire n609;
   wire n610;
   wire n611;
   wire n612;
   wire n613;
   wire n614;
   wire n615;
   wire n616;
   wire n617;
   wire n618;
   wire n619;
   wire n620;
   wire n621;
   wire n622;
   wire n623;
   wire n624;
   wire n625;
   wire n626;
   wire n627;
   wire n628;
   wire n629;
   wire n630;
   wire n631;
   wire n632;
   wire n633;
   wire n634;
   wire n635;
   wire n636;
   wire n637;
   wire n638;
   wire n639;
   wire n640;
   wire n641;
   wire n642;
   wire n643;
   wire n644;
   wire n645;
   wire n646;
   wire n647;
   wire n648;
   wire n649;
   wire n650;
   wire n651;
   wire n652;
   wire n653;
   wire n654;
   wire n655;
   wire n656;
   wire n657;
   wire n658;
   wire n659;
   wire n660;
   wire n661;
   wire n662;
   wire n663;
   wire n664;
   wire n665;
   wire n666;
   wire n667;
   wire n668;
   wire n669;
   wire n670;
   wire n671;
   wire n672;
   wire n673;
   wire n674;
   wire n675;
   wire n676;
   wire n677;
   wire n678;
   wire n679;
   wire n680;
   wire n681;
   wire n682;
   wire n683;
   wire n684;
   wire n685;
   wire n686;
   wire n687;
   wire n688;
   wire n689;
   wire n690;
   wire n691;
   wire n692;
   wire n693;
   wire n694;
   wire n695;
   wire n696;
   wire n697;
   wire n698;
   wire n699;
   wire n700;
   wire n701;
   wire n702;
   wire n703;
   wire n704;
   wire n705;
   wire n706;
   wire n707;
   wire n708;
   wire n709;
   wire n710;
   wire n711;
   wire n712;
   wire n713;
   wire n714;
   wire n715;
   wire n716;
   wire n717;
   wire n718;
   wire n719;
   wire n720;
   wire n721;
   wire n722;
   wire n723;
   wire n724;
   wire n725;
   wire n726;
   wire n727;
   wire n728;
   wire n729;
   wire n730;
   wire n731;
   wire n732;
   wire n733;
   wire n734;
   wire n735;
   wire n736;
   wire n737;
   wire n738;
   wire n739;
   wire n740;
   wire n741;
   wire n742;
   wire n743;
   wire n744;
   wire n745;
   wire n746;
   wire n747;
   wire n748;
   wire n749;
   wire n750;
   wire n751;
   wire n752;
   wire n753;
   wire n754;
   wire n755;
   wire n756;
   wire n757;
   wire n758;
   wire n759;
   wire n760;
   wire n761;
   wire n762;
   wire n763;
   wire n764;
   wire n765;
   wire n766;
   wire n767;
   wire n768;
   wire n769;
   wire n770;
   wire n771;
   wire n772;
   wire n773;
   wire n774;
   wire n775;
   wire n776;
   wire n777;
   wire n778;
   wire n779;
   wire n780;
   wire n781;
   wire n782;
   wire n783;
   wire n784;
   wire n785;
   wire n786;
   wire n787;
   wire n788;
   wire n789;
   wire n790;
   wire n791;
   wire n792;
   wire n793;
   wire n794;
   wire n795;
   wire n796;
   wire n797;
   wire n798;
   wire n799;
   wire n800;
   wire n801;
   wire n802;
   wire n803;
   wire n804;
   wire n805;
   wire n806;
   wire n807;
   wire n808;
   wire n809;
   wire n810;
   wire n811;
   wire n812;
   wire n813;
   wire n814;
   wire n815;
   wire n816;
   wire n817;
   wire n818;
   wire n819;
   wire n820;
   wire n821;
   wire n822;
   wire n823;
   wire n824;
   wire n825;
   wire n826;
   wire n827;
   wire n828;
   wire n829;
   wire n830;
   wire n831;
   wire n832;
   wire n833;
   wire n834;
   wire n835;
   wire n836;
   wire n837;
   wire n838;
   wire n839;
   wire n840;
   wire n841;
   wire n842;
   wire n843;
   wire n844;
   wire n845;
   wire n846;
   wire n847;
   wire n848;
   wire n849;
   wire n850;
   wire n851;
   wire n852;
   wire n853;
   wire n854;
   wire n855;
   wire n856;
   wire n857;
   wire n858;
   wire n859;
   wire n860;
   wire n861;
   wire n862;
   wire n863;
   wire n864;
   wire n865;
   wire n866;
   wire n867;
   wire n868;
   wire n869;
   wire n870;
   wire n871;
   wire n872;
   wire n873;
   wire n874;
   wire n875;
   wire n876;
   wire n877;
   wire n878;
   wire n879;
   wire n880;
   wire n881;
   wire n882;
   wire n883;
   wire n884;
   wire n885;
   wire n886;
   wire n887;
   wire n888;
   wire n889;

   assign FLAGS[3] = \*Logic0*  ;
   assign Z[6] = net3712 ;
   assign Z[7] = net3715 ;
   assign Z[8] = net3718 ;
   assign Z[9] = net3721 ;
   assign Z[31] = net3724 ;
   assign Z[3] = net3727 ;
   assign Z[4] = net3730 ;
   assign Z[5] = net3733 ;
   assign Z[28] = net3736 ;
   assign Z[29] = net3739 ;
   assign Z[2] = net3742 ;
   assign Z[30] = net3745 ;
   assign Z[24] = net3748 ;
   assign Z[25] = net3751 ;
   assign Z[26] = net3754 ;
   assign Z[27] = net3757 ;

   SEN_ND2_3 U471 (.X(n780), 
	.A2(n619), 
	.A1(net16476));
   SEN_ND2_T_1 U472 (.X(n474), 
	.A2(n473), 
	.A1(n472));
   SEN_ND2_G_1 U473 (.X(n472), 
	.A2(n471), 
	.A1(net16482));
   SEN_ND2_S_2 U474 (.X(n647), 
	.A2(n554), 
	.A1(n641));
   SEN_AOAI211_6 U475 (.X(n855), 
	.C(n848), 
	.B(n666), 
	.A2(n667), 
	.A1(n543));
   SEN_OAI21_T_4 U476 (.X(n666), 
	.B(n532), 
	.A2(n847), 
	.A1(n533));
   SEN_INV_AS_5 U477 (.X(n667), 
	.A(n838));
   SEN_INV_1 U478 (.X(n847), 
	.A(n746));
   SEN_ND2_2 U479 (.X(n746), 
	.A2(n663), 
	.A1(n662));
   SEN_NR2_T_5 U480 (.X(n610), 
	.A2(net15882), 
	.A1(n772));
   SEN_ND2_T_5 U481 (.X(n643), 
	.A2(n527), 
	.A1(n360));
   SEN_INV_S_3 U482 (.X(n818), 
	.A(n638));
   SEN_INV_4 U483 (.X(n672), 
	.A(n855));
   SEN_INV_3 U484 (.X(n843), 
	.A(n665));
   SEN_ND2_G_1 U485 (.X(n759), 
	.A2(n648), 
	.A1(n649));
   SEN_OAI21_2 U486 (.X(n559), 
	.B(n558), 
	.A2(net16400), 
	.A1(n703));
   SEN_INV_4 U487 (.X(n703), 
	.A(n557));
   SEN_INV_4 U488 (.X(n552), 
	.A(n698));
   SEN_ND2_1P5 U489 (.X(n691), 
	.A2(n885), 
	.A1(n690));
   SEN_ND2_S_6 U490 (.X(n397), 
	.A2(net15940), 
	.A1(net15941));
   SEN_OAI211_2 U491 (.X(net3721), 
	.B2(net15886), 
	.B1(net15885), 
	.A2(net16410), 
	.A1(net15884));
   SEN_EN2_S_2 U492 (.X(net15884), 
	.A2(n824), 
	.A1(n523));
   SEN_INV_S_6 U493 (.X(n358), 
	.A(n651));
   SEN_ND2_T_4 U494 (.X(n651), 
	.A2(n554), 
	.A1(n635));
   SEN_INV_S_0P5 U495 (.X(n835), 
	.A(n651));
   SEN_ND2_T_0P5 U496 (.X(n454), 
	.A2(net16152), 
	.A1(net16085));
   SEN_ND2_G_4 U497 (.X(n533), 
	.A2(n456), 
	.A1(n455));
   SEN_MUXI2_DG_2 U498 (.X(n593), 
	.S(A[17]), 
	.D1(net16669), 
	.D0(net16480));
   SEN_INV_5 U499 (.X(net16311), 
	.A(net16499));
   SEN_AN3_0P5 U500 (.X(n359), 
	.A3(net16501), 
	.A2(n703), 
	.A1(net16311));
   SEN_OAI211_3 U501 (.X(Z[23]), 
	.B2(net15787), 
	.B1(net15786), 
	.A2(net16410), 
	.A1(net15785));
   SEN_OAI211_2 U502 (.X(net3751), 
	.B2(net16146), 
	.B1(net16145), 
	.A2(net16410), 
	.A1(net16144));
   SEN_OAI21B_4 U503 (.X(net3739), 
	.B(n386), 
	.A2(net16410), 
	.A1(net16113));
   SEN_OR3_8 U504 (.X(net15916), 
	.A3(net17773), 
	.A2(net16282), 
	.A1(net16281));
   SEN_ND2_2 U505 (.X(n884), 
	.A2(n464), 
	.A1(n463));
   SEN_INV_S_2 U506 (.X(net16010), 
	.A(net16336));
   SEN_AOI31_4 U507 (.X(n738), 
	.B(n735), 
	.A3(n736), 
	.A2(n885), 
	.A1(n737));
   SEN_INV_1 U508 (.X(net15881), 
	.A(net15897));
   SEN_OAI21_G_4 U509 (.X(n871), 
	.B(n868), 
	.A2(n869), 
	.A1(n870));
   SEN_ND2_T_1 U510 (.X(n668), 
	.A2(n587), 
	.A1(n553));
   SEN_ND2_3 U511 (.X(net16289), 
	.A2(n628), 
	.A1(net16474));
   SEN_MUXI2_S_3 U512 (.X(n628), 
	.S(A[2]), 
	.D1(n549), 
	.D0(net16482));
   SEN_INV_S_3 U513 (.X(net16281), 
	.A(net16015));
   SEN_NR3_T_4 U514 (.X(net16293), 
	.A3(net16287), 
	.A2(net15985), 
	.A1(net16284));
   SEN_ND2_S_6 U515 (.X(net15985), 
	.A2(n506), 
	.A1(n505));
   SEN_INV_6 U516 (.X(n549), 
	.A(n504));
   SEN_INV_2 U517 (.X(n834), 
	.A(n758));
   SEN_NR2_G_2 U518 (.X(n653), 
	.A2(n758), 
	.A1(n534));
   SEN_AOI211_G_5 U519 (.X(n611), 
	.B2(n770), 
	.B1(n610), 
	.A2(n370), 
	.A1(n771));
   SEN_INV_4 U520 (.X(n370), 
	.A(n369));
   SEN_BUF_8 U521 (.X(net16499), 
	.A(INST[1]));
   SEN_ND2_T_1 U522 (.X(n704), 
	.A2(net16499), 
	.A1(net16501));
   SEN_INV_1P25 U523 (.X(n511), 
	.A(n512));
   SEN_ND2_2 U524 (.X(n394), 
	.A2(net16499), 
	.A1(net16495));
   SEN_INV_4 U525 (.X(n782), 
	.A(n620));
   SEN_ND2_G_3 U526 (.X(net15769), 
	.A2(n561), 
	.A1(n489));
   SEN_ND2_S_3 U527 (.X(n376), 
	.A2(n786), 
	.A1(n791));
   SEN_ND2_1P5 U528 (.X(n792), 
	.A2(n786), 
	.A1(n787));
   SEN_NR2_T_1 U529 (.X(n561), 
	.A2(net16501), 
	.A1(net16497));
   SEN_INV_S_2 U530 (.X(n428), 
	.A(net3715));
   SEN_ND2_T_2 U531 (.X(n617), 
	.A2(n614), 
	.A1(n554));
   SEN_MUXI2_S_3 U532 (.X(n396), 
	.S(A[4]), 
	.D1(net16669), 
	.D0(net16482));
   SEN_INV_6 U533 (.X(net16486), 
	.A(net16200));
   SEN_INV_3 U534 (.X(n381), 
	.A(Z[17]));
   SEN_OAI211_4 U535 (.X(net3757), 
	.B2(net15763), 
	.B1(net15762), 
	.A2(net16412), 
	.A1(net15760));
   SEN_ND3_T_2 U536 (.X(n799), 
	.A3(n796), 
	.A2(net15973), 
	.A1(n797));
   SEN_ND2_6 U537 (.X(net16292), 
	.A2(net16476), 
	.A1(n396));
   SEN_INV_5 U538 (.X(n491), 
	.A(n490));
   SEN_INV_2 U539 (.X(n518), 
	.A(n512));
   SEN_EN2_8 U540 (.X(n878), 
	.A2(n810), 
	.A1(n811));
   SEN_ND2_4 U541 (.X(net15760), 
	.A2(n547), 
	.A1(n548));
   SEN_INV_2 U542 (.X(n360), 
	.A(net15915));
   SEN_INV_4 U543 (.X(net16057), 
	.A(net15915));
   SEN_ND2_G_1 U544 (.X(net16014), 
	.A2(net16298), 
	.A1(net17648));
   SEN_INV_2 U545 (.X(n767), 
	.A(n544));
   SEN_INV_S_1P5 U546 (.X(n768), 
	.A(n632));
   SEN_ND2_S_6 U547 (.X(net15961), 
	.A2(net15946), 
	.A1(net15945));
   SEN_INV_4 U548 (.X(net15940), 
	.A(net16292));
   SEN_EN2_S_4 U549 (.X(n771), 
	.A2(net16009), 
	.A1(net16010));
   SEN_ND2_T_2 U550 (.X(n510), 
	.A2(n509), 
	.A1(n508));
   SEN_AOI222_1 U551 (.X(net16087), 
	.C2(n740), 
	.C1(n741), 
	.B2(n374), 
	.B1(net17584), 
	.A2(n742), 
	.A1(n451));
   SEN_NR2_T_5 U552 (.X(n451), 
	.A2(n499), 
	.A1(n560));
   SEN_MUXI2_S_4 U553 (.X(n603), 
	.S(A[7]), 
	.D1(net16669), 
	.D0(net16480));
   SEN_ND2_T_3 U554 (.X(net15865), 
	.A2(net16062), 
	.A1(net15916));
   SEN_INV_S_8 U555 (.X(net16480), 
	.A(net16486));
   SEN_MUXI2_S_4 U556 (.X(n602), 
	.S(B[7]), 
	.D1(n493), 
	.D0(n550));
   SEN_OAI211_3 U557 (.X(Z[11]), 
	.B2(net16030), 
	.B1(net16029), 
	.A2(net16412), 
	.A1(net16028));
   SEN_EN2_5 U558 (.X(n770), 
	.A2(net16020), 
	.A1(net16021));
   SEN_ND2_T_6 U559 (.X(n838), 
	.A2(net17669), 
	.A1(n878));
   SEN_INV_S_3 U560 (.X(net17668), 
	.A(net15784));
   SEN_ND2_3 U561 (.X(net15784), 
	.A2(n361), 
	.A1(n660));
   SEN_ND2_T_4 U562 (.X(n607), 
	.A2(n604), 
	.A1(n554));
   SEN_ND2_T_5 U563 (.X(n772), 
	.A2(net17656), 
	.A1(n804));
   SEN_ND2_S_1P5 U564 (.X(n547), 
	.A2(n885), 
	.A1(n537));
   SEN_INV_AS_10 U565 (.X(net16482), 
	.A(net16486));
   SEN_INV_3 U566 (.X(n755), 
	.A(n649));
   SEN_ND2_T_2 U567 (.X(n456), 
	.A2(n881), 
	.A1(n662));
   SEN_INV_1P25 U568 (.X(n881), 
	.A(n663));
   SEN_ND2_S_0P5 U569 (.X(n883), 
	.A2(n539), 
	.A1(net16434));
   SEN_OA21_4 U570 (.X(net17713), 
	.B(n883), 
	.A2(net16410), 
	.A1(n884));
   SEN_OAI21_2 U571 (.X(n822), 
	.B(n821), 
	.A2(net15882), 
	.A1(n521));
   SEN_NR2_S_1 U572 (.X(n823), 
	.A2(net15882), 
	.A1(net15881));
   SEN_NR3_T_0P8 U573 (.X(n826), 
	.A3(net15883), 
	.A2(net15882), 
	.A1(net15881));
   SEN_ND3_T_1 U574 (.X(n401), 
	.A3(n370), 
	.A2(net15894), 
	.A1(net15880));
   SEN_INV_5 U575 (.X(net15882), 
	.A(n370));
   SEN_ND2_T_2 U576 (.X(net16322), 
	.A2(net16337), 
	.A1(net16336));
   SEN_MUXI2_S_4 U577 (.X(n629), 
	.S(B[4]), 
	.D1(n493), 
	.D0(n551));
   SEN_INV_5 U578 (.X(n493), 
	.A(n512));
   SEN_OA21_4 U579 (.X(n652), 
	.B(n760), 
	.A2(n759), 
	.A1(n758));
   SEN_ND2_G_0P65 U580 (.X(net16153), 
	.A2(n681), 
	.A1(n680));
   SEN_INV_S_2 U581 (.X(n743), 
	.A(n680));
   SEN_ND2_G_2 U582 (.X(n488), 
	.A2(net16495), 
	.A1(net16311));
   SEN_ND2_G_1 U583 (.X(n361), 
	.A2(n597), 
	.A1(net17602));
   SEN_ND2_2 U584 (.X(n661), 
	.A2(n597), 
	.A1(net17602));
   SEN_MUXI2_S_2 U585 (.X(n597), 
	.S(A[16]), 
	.D1(net16669), 
	.D0(net16480));
   SEN_INV_2 U586 (.X(net15973), 
	.A(net15985));
   SEN_ND2_T_4 U587 (.X(n796), 
	.A2(n377), 
	.A1(n787));
   SEN_AN2_DG_2 U588 (.X(net16949), 
	.A2(net16292), 
	.A1(net16291));
   SEN_BUF_1 U589 (.X(n362), 
	.A(n847));
   SEN_INV_4 U590 (.X(n807), 
	.A(n606));
   SEN_ND2_T_4 U591 (.X(n606), 
	.A2(n605), 
	.A1(net17602));
   SEN_INV_S_6 U592 (.X(n806), 
	.A(n607));
   SEN_INV_8 U593 (.X(n683), 
	.A(n504));
   SEN_NR2B_V1_8 U594 (.X(n504), 
	.B(net17414), 
	.A(net16179));
   SEN_EO2_6 U595 (.X(net15945), 
	.A2(net15967), 
	.A1(net16300));
   SEN_ND2_S_2 U596 (.X(n459), 
	.A2(n816), 
	.A1(net16985));
   SEN_ND2_G_1 U597 (.X(net16407), 
	.A2(net16408), 
	.A1(net16311));
   SEN_INV_2 U598 (.X(n781), 
	.A(n622));
   SEN_NR2_S_4 U599 (.X(n623), 
	.A2(n781), 
	.A1(n780));
   SEN_NR3_T_6 U600 (.X(n412), 
	.A3(n414), 
	.A2(net3757), 
	.A1(n388));
   SEN_INV_3 U601 (.X(n450), 
	.A(n611));
   SEN_EN2_S_6 U602 (.X(net16113), 
	.A2(n722), 
	.A1(n737));
   SEN_OAI211_3 U603 (.X(n720), 
	.B2(n736), 
	.B1(net16125), 
	.A2(n719), 
	.A1(net16123));
   SEN_ND2_T_2 U604 (.X(n616), 
	.A2(n615), 
	.A1(net16476));
   SEN_INV_3 U605 (.X(n377), 
	.A(n376));
   SEN_ND2_2 U606 (.X(n791), 
	.A2(n616), 
	.A1(n617));
   SEN_ND2_S_4 U607 (.X(n405), 
	.A2(n410), 
	.A1(n409));
   SEN_INV_2P5 U608 (.X(n811), 
	.A(n661));
   SEN_INV_4 U609 (.X(n553), 
	.A(n556));
   SEN_ND2_S_4 U610 (.X(n662), 
	.A2(n553), 
	.A1(n592));
   SEN_ND2_T_2 U611 (.X(n664), 
	.A2(n590), 
	.A1(n553));
   SEN_ND2_S_4 U612 (.X(n414), 
	.A2(n416), 
	.A1(n415));
   SEN_MUXI2_DG_2 U613 (.X(n631), 
	.S(A[11]), 
	.D1(net16669), 
	.D0(net16482));
   SEN_OAI211_3 U614 (.X(Z[19]), 
	.B2(net15832), 
	.B1(net15831), 
	.A2(net16410), 
	.A1(net15830));
   SEN_ND2_S_3 U615 (.X(net16299), 
	.A2(n612), 
	.A1(n554));
   SEN_MUXI2_DG_3 U616 (.X(n612), 
	.S(B[5]), 
	.D1(n518), 
	.D0(n551));
   SEN_INV_S_4 U617 (.X(n499), 
	.A(n498));
   SEN_ND2B_V1_2 U618 (.X(n560), 
	.B(net16495), 
	.A(net16501));
   SEN_OAI21_5 U619 (.X(net3745), 
	.B(net16087), 
	.A2(net16410), 
	.A1(net16086));
   SEN_ND2_6 U620 (.X(n532), 
	.A2(n385), 
	.A1(n384));
   SEN_NR2_S_3 U621 (.X(n498), 
	.A2(net16497), 
	.A1(net16311));
   SEN_ND2_T_4 U622 (.X(net16301), 
	.A2(net17602), 
	.A1(n626));
   SEN_ND2_S_0P5 U623 (.X(n867), 
	.A2(n856), 
	.A1(n855));
   SEN_OAI21_S_1P5 U624 (.X(n803), 
	.B(net15946), 
	.A2(net18184), 
	.A1(n531));
   SEN_INV_4 U625 (.X(n836), 
	.A(n650));
   SEN_ND3_S_8 U626 (.X(n419), 
	.A3(n422), 
	.A2(n421), 
	.A1(n420));
   SEN_ND2_T_2 U627 (.X(n478), 
	.A2(B[18]), 
	.A1(n518));
   SEN_OAI21_G_2 U628 (.X(n876), 
	.B(net15795), 
	.A2(net15794), 
	.A1(n875));
   SEN_INV_S_1 U629 (.X(net15960), 
	.A(net15961));
   SEN_ND2_3 U630 (.X(n506), 
	.A2(net17420), 
	.A1(net16288));
   SEN_INV_4 U631 (.X(net17420), 
	.A(net15979));
   SEN_ND2_T_2 U632 (.X(n663), 
	.A2(n593), 
	.A1(net16476));
   SEN_AN3_4 U633 (.X(net18229), 
	.A3(net16501), 
	.A2(n703), 
	.A1(net17564));
   SEN_ND2_S_6 U634 (.X(n864), 
	.A2(n371), 
	.A1(n846));
   SEN_INV_AS_10 U635 (.X(n846), 
	.A(n839));
   SEN_EO2_1 U636 (.X(net15919), 
	.A2(n519), 
	.A1(n809));
   SEN_OAI21_5 U637 (.X(net16073), 
	.B(n522), 
	.A2(n747), 
	.A1(n675));
   SEN_INV_S_4 U638 (.X(net15941), 
	.A(net16291));
   SEN_EN2_S_3 U639 (.X(n865), 
	.A2(n861), 
	.A1(n860));
   SEN_INV_S_3 U640 (.X(n860), 
	.A(n670));
   SEN_INV_2 U641 (.X(n800), 
	.A(n799));
   SEN_ND2_4 U642 (.X(net16064), 
	.A2(n477), 
	.A1(n476));
   SEN_INV_S_6 U643 (.X(n413), 
	.A(net3745));
   SEN_ND2_S_4 U644 (.X(n620), 
	.A2(n554), 
	.A1(n618));
   SEN_INV_S_2 U645 (.X(n886), 
	.A(n580));
   SEN_BUF_1 U646 (.X(n363), 
	.A(n499));
   SEN_EN2_3 U647 (.X(net15799), 
	.A2(n871), 
	.A1(n522));
   SEN_NR3_T_3 U648 (.X(n433), 
	.A3(Z[1]), 
	.A2(Z[0]), 
	.A1(net3742));
   SEN_OAI211_1 U649 (.X(Z[0]), 
	.B2(net15997), 
	.B1(net15996), 
	.A2(net16412), 
	.A1(net15995));
   SEN_EO2_1 U650 (.X(n524), 
	.A2(n783), 
	.A1(n782));
   SEN_INV_1P25 U651 (.X(net16408), 
	.A(net16497));
   SEN_ND2_T_4 U652 (.X(net16179), 
	.A2(net16309), 
	.A1(net16501));
   SEN_INV_10 U653 (.X(n554), 
	.A(n556));
   SEN_INV_S_8 U654 (.X(n556), 
	.A(n700));
   SEN_INV_0P5 U655 (.X(n778), 
	.A(n771));
   SEN_ND2_4 U656 (.X(net17189), 
	.A2(n797), 
	.A1(net16293));
   SEN_AOI211_G_2 U657 (.X(n801), 
	.B2(net15958), 
	.B1(net16949), 
	.A2(net15956), 
	.A1(n800));
   SEN_AN2_S_1P5 U658 (.X(n534), 
	.A2(n752), 
	.A1(n492));
   SEN_ND2_T_1 U659 (.X(n476), 
	.A2(net17000), 
	.A1(n749));
   SEN_ND2_3 U660 (.X(net16200), 
	.A2(net16395), 
	.A1(n563));
   SEN_EO2_DG_1 U661 (.X(net15995), 
	.A2(n524), 
	.A1(n781));
   SEN_OAOI211_4 U662 (.X(n440), 
	.C(net16143), 
	.B(net17035), 
	.A2(n442), 
	.A1(n441));
   SEN_INV_1 U663 (.X(net16009), 
	.A(net16337));
   SEN_MUXI2_S_6 U664 (.X(n604), 
	.S(B[6]), 
	.D1(n493), 
	.D0(n551));
   SEN_OAI211_4 U665 (.X(Z[12]), 
	.B2(net16053), 
	.B1(net16052), 
	.A2(net16412), 
	.A1(net16051));
   SEN_INV_2P5 U666 (.X(n494), 
	.A(n512));
   SEN_ND2_T_3 U667 (.X(n441), 
	.A2(net16154), 
	.A1(net16127));
   SEN_INV_0P65 U668 (.X(n368), 
	.A(n512));
   SEN_INV_2 U669 (.X(n517), 
	.A(n512));
   SEN_NR3_T_6 U670 (.X(n420), 
	.A3(Z[14]), 
	.A2(n445), 
	.A1(Z[12]));
   SEN_ND2_S_2 U671 (.X(n820), 
	.A2(net16014), 
	.A1(net16015));
   SEN_AN2_S_1 U672 (.X(n521), 
	.A2(n375), 
	.A1(n778));
   SEN_ND2_S_1 U673 (.X(n375), 
	.A2(net17656), 
	.A1(n804));
   SEN_ND2B_V1_4 U674 (.X(net16291), 
	.B(n629), 
	.A(n556));
   SEN_INV_3 U675 (.X(net16282), 
	.A(net15897));
   SEN_ND2_2 U676 (.X(n502), 
	.A2(B[2]), 
	.A1(n494));
   SEN_ND2_T_2 U677 (.X(n503), 
	.A2(n501), 
	.A1(n502));
   SEN_AOAI211_2 U678 (.X(n824), 
	.C(net15894), 
	.B(n822), 
	.A2(n823), 
	.A1(n526));
   SEN_ND2_2 U679 (.X(net16074), 
	.A2(n674), 
	.A1(n673));
   SEN_EN2_S_4 U680 (.X(net15915), 
	.A2(n756), 
	.A1(n755));
   SEN_INV_3 U681 (.X(n654), 
	.A(n832));
   SEN_ND2_G_1 U682 (.X(net16154), 
	.A2(net16192), 
	.A1(net16191));
   SEN_ND2_T_2 U683 (.X(n689), 
	.A2(n719), 
	.A1(net16125));
   SEN_ND2_T_4 U684 (.X(n385), 
	.A2(n843), 
	.A1(n383));
   SEN_INV_S_4 U685 (.X(n842), 
	.A(n664));
   SEN_ND2_T_1 U686 (.X(n656), 
	.A2(n633), 
	.A1(n554));
   SEN_ND2_T_2 U687 (.X(n649), 
	.A2(n639), 
	.A1(n554));
   SEN_ND2_S_4 U688 (.X(net16300), 
	.A2(n554), 
	.A1(n625));
   SEN_AO21B_1 U689 (.X(n869), 
	.B(n859), 
	.A2(n866), 
	.A1(n867));
   SEN_ND2_2 U690 (.X(net17550), 
	.A2(net16292), 
	.A1(net16291));
   SEN_ND2_6 U691 (.X(net16287), 
	.A2(net17550), 
	.A1(n397));
   SEN_INV_1P25 U692 (.X(n828), 
	.A(n647));
   SEN_ND2_T_1 U693 (.X(n752), 
	.A2(n646), 
	.A1(n647));
   SEN_EN2_S_3 U694 (.X(net15785), 
	.A2(n876), 
	.A1(net17005));
   SEN_INV_S_3 U695 (.X(n788), 
	.A(n617));
   SEN_INV_4 U696 (.X(net15953), 
	.A(net16284));
   SEN_INV_S_6 U697 (.X(n410), 
	.A(net3739));
   SEN_INV_0P8 U698 (.X(n736), 
	.A(n718));
   SEN_INV_3 U699 (.X(n445), 
	.A(n444));
   SEN_INV_S_2 U700 (.X(n793), 
	.A(n785));
   SEN_OAI211_4 U701 (.X(net3712), 
	.B2(net15929), 
	.B1(net15928), 
	.A2(net16412), 
	.A1(net15927));
   SEN_ND2_S_4 U702 (.X(net3718), 
	.A2(net16018), 
	.A1(net17804));
   SEN_ND2_8 U703 (.X(n751), 
	.A2(net15880), 
	.A1(n380));
   SEN_INV_2 U704 (.X(net16020), 
	.A(net16328));
   SEN_ND2_T_2 U705 (.X(net16328), 
	.A2(net17602), 
	.A1(n609));
   SEN_MUXI2_DG_2 U706 (.X(n609), 
	.S(A[8]), 
	.D1(n683), 
	.D0(net16482));
   SEN_AO21B_2 U707 (.X(n711), 
	.B(net16153), 
	.A2(net16084), 
	.A1(n441));
   SEN_EN2_3 U708 (.X(net16152), 
	.A2(n744), 
	.A1(n743));
   SEN_INV_2P5 U709 (.X(net16084), 
	.A(net16152));
   SEN_INV_6 U710 (.X(net16361), 
	.A(net16177));
   SEN_INV_S_4 U711 (.X(n430), 
	.A(net3718));
   SEN_ND2_S_2 U712 (.X(n453), 
	.A2(net17843), 
	.A1(net16084));
   SEN_INV_S_4 U713 (.X(n817), 
	.A(n637));
   SEN_ND2_S_3 U714 (.X(n637), 
	.A2(n594), 
	.A1(n555));
   SEN_INV_6 U715 (.X(net15942), 
	.A(net16287));
   SEN_INV_S_0P5 U716 (.X(n364), 
	.A(net17668));
   SEN_INV_S_0P5 U717 (.X(n365), 
	.A(net17668));
   SEN_INV_4 U718 (.X(net17669), 
	.A(net17668));
   SEN_INV_S_3 U719 (.X(n369), 
	.A(net16322));
   SEN_NR2_T_1P5 U720 (.X(n495), 
	.A2(n765), 
	.A1(n530));
   SEN_AOAI211_G_2 U721 (.X(n827), 
	.C(net15880), 
	.B(n380), 
	.A2(n826), 
	.A1(n526));
   SEN_ND2_T_6 U722 (.X(n380), 
	.A2(n523), 
	.A1(n457));
   SEN_EO2_S_3 U723 (.X(net16086), 
	.A2(n738), 
	.A1(n742));
   SEN_ND2_T_6 U724 (.X(n885), 
	.A2(n689), 
	.A1(n514));
   SEN_NR2_T_4 U725 (.X(n514), 
	.A2(n470), 
	.A1(net17788));
   SEN_MUXI2_S_1 U726 (.X(n687), 
	.S(B[26]), 
	.D1(n367), 
	.D0(n551));
   SEN_MUX2_DG_1 U727 (.X(n635), 
	.S(n541), 
	.D1(n552), 
	.D0(n512));
   SEN_MUXI2_S_3 U728 (.X(n615), 
	.S(A[1]), 
	.D1(n683), 
	.D0(net16482));
   SEN_OAI211_3 U729 (.X(Z[21]), 
	.B2(net15801), 
	.B1(net15800), 
	.A2(net16410), 
	.A1(net15799));
   SEN_OR2_5 U730 (.X(n513), 
	.A2(n497), 
	.A1(net18229));
   SEN_INV_0P65 U731 (.X(net15913), 
	.A(net15914));
   SEN_ND2_T_8 U732 (.X(n839), 
	.A2(net16077), 
	.A1(net15796));
   SEN_ND2_8 U733 (.X(net15796), 
	.A2(net16985), 
	.A1(net15914));
   SEN_EO2_G_2 U734 (.X(net15975), 
	.A2(n794), 
	.A1(net15973));
   SEN_EN2_3 U735 (.X(n845), 
	.A2(n853), 
	.A1(n852));
   SEN_INV_S_2 U736 (.X(n852), 
	.A(n668));
   SEN_ND2_6 U737 (.X(n660), 
	.A2(n596), 
	.A1(n553));
   SEN_INV_3 U738 (.X(n407), 
	.A(net3754));
   SEN_INV_4 U739 (.X(n596), 
	.A(n510));
   SEN_EN2_6 U740 (.X(net16284), 
	.A2(net16298), 
	.A1(net17648));
   SEN_ND3_T_1P5 U741 (.X(net16395), 
	.A3(net17573), 
	.A2(net16968), 
	.A1(n389));
   SEN_MUXI2_S_3 U742 (.X(n639), 
	.S(B[12]), 
	.D1(n517), 
	.D0(n551));
   SEN_INV_0P8 U743 (.X(net17843), 
	.A(net16085));
   SEN_EO2_5 U744 (.X(n787), 
	.A2(n624), 
	.A1(n623));
   SEN_OAI21_S_3 U745 (.X(n879), 
	.B(n364), 
	.A2(n378), 
	.A1(n519));
   SEN_NR2_2 U746 (.X(n850), 
	.A2(n362), 
	.A1(net15797));
   SEN_INV_S_4 U747 (.X(n417), 
	.A(Z[22]));
   SEN_EN2_3 U748 (.X(net16051), 
	.A2(n754), 
	.A1(n360));
   SEN_OAI211_4 U749 (.X(Z[22]), 
	.B2(net16066), 
	.B1(net16065), 
	.A2(net16412), 
	.A1(net16064));
   SEN_OR2_2P5 U750 (.X(n754), 
	.A2(n496), 
	.A1(n495));
   SEN_INV_S_2 U751 (.X(n366), 
	.A(n494));
   SEN_INV_3 U752 (.X(n367), 
	.A(n366));
   SEN_ND2_1P5 U753 (.X(n786), 
	.A2(n620), 
	.A1(n780));
   SEN_ND2_S_4 U754 (.X(n624), 
	.A2(n622), 
	.A1(n782));
   SEN_AOAI211_3 U755 (.X(n851), 
	.C(n848), 
	.B(n849), 
	.A2(n850), 
	.A1(n525));
   SEN_ND3_T_1 U756 (.X(net15934), 
	.A3(net16014), 
	.A2(net16015), 
	.A1(net15897));
   SEN_OAI21_S_3 U757 (.X(n777), 
	.B(net17656), 
	.A2(n804), 
	.A1(net16013));
   SEN_INV_S_6 U758 (.X(n409), 
	.A(net3736));
   SEN_OAI211_8 U759 (.X(net3736), 
	.B2(net16104), 
	.B1(net16103), 
	.A2(n443), 
	.A1(net16102));
   SEN_EO2_G_8 U760 (.X(net16102), 
	.A2(n727), 
	.A1(n535));
   SEN_ND2_T_1 U761 (.X(net17572), 
	.A2(A[31]), 
	.A1(net16497));
   SEN_NR2_G_1 U762 (.X(n391), 
	.A2(net16495), 
	.A1(net16497));
   SEN_BUF_8 U763 (.X(net16497), 
	.A(INST[2]));
   SEN_ND2_2 U764 (.X(net15971), 
	.A2(net16289), 
	.A1(net16288));
   SEN_INV_2 U765 (.X(net16085), 
	.A(n441));
   SEN_AO21B_6 U766 (.X(n399), 
	.B(net15942), 
	.A2(net15946), 
	.A1(net15971));
   SEN_AN2_3 U767 (.X(n531), 
	.A2(n799), 
	.A1(net15971));
   SEN_INV_S_4 U768 (.X(n416), 
	.A(Z[19]));
   SEN_INV_S_4 U769 (.X(n422), 
	.A(Z[18]));
   SEN_ND2_2 U770 (.X(n505), 
	.A2(net15979), 
	.A1(net15980));
   SEN_INV_S_2 U771 (.X(net15980), 
	.A(net16288));
   SEN_INV_S_4 U772 (.X(net16062), 
	.A(net15910));
   SEN_ND2_T_3 U773 (.X(net15910), 
	.A2(n527), 
	.A1(n751));
   SEN_BUF_S_6 U774 (.X(net17648), 
	.A(net16299));
   SEN_ND2_S_1 U775 (.X(n468), 
	.A2(n777), 
	.A1(n778));
   SEN_INV_S_2 U776 (.X(net17600), 
	.A(net16180));
   SEN_MUXI2_DG_3 U777 (.X(n618), 
	.S(B[0]), 
	.D1(n511), 
	.D0(n551));
   SEN_OAI211_3 U778 (.X(net3742), 
	.B2(net15977), 
	.B1(net15976), 
	.A2(net16412), 
	.A1(net15975));
   SEN_MUXI2_S_0P5 U779 (.X(n682), 
	.S(B[25]), 
	.D1(n494), 
	.D0(n550));
   SEN_OAI21B_2 U780 (.X(n833), 
	.B(n831), 
	.A2(n832), 
	.A1(net15865));
   SEN_ND2_T_4 U781 (.X(net16215), 
	.A2(net15795), 
	.A1(net15794));
   SEN_ND2_G_1 U782 (.X(net15795), 
	.A2(net16222), 
	.A1(net16223));
   SEN_NR3B_DG_8 U783 (.X(n645), 
	.B2(n643), 
	.B1(n644), 
	.A(n813));
   SEN_ND2_S_1P5 U784 (.X(n402), 
	.A2(net17656), 
	.A1(net16014));
   SEN_EN2_8 U785 (.X(n758), 
	.A2(n836), 
	.A1(n358));
   SEN_MUXI2_S_1 U786 (.X(n594), 
	.S(B[15]), 
	.D1(n494), 
	.D0(n550));
   SEN_ND4_S_3 U787 (.X(net15798), 
	.A4(n364), 
	.A3(net16077), 
	.A2(net16345), 
	.A1(net16344));
   SEN_ND2_S_1 U788 (.X(net16023), 
	.A2(net15897), 
	.A1(net17656));
   SEN_OAI21_5 U789 (.X(net15914), 
	.B(n657), 
	.A2(n658), 
	.A1(n659));
   SEN_INV_2 U790 (.X(n442), 
	.A(net16153));
   SEN_EN2_8 U791 (.X(n804), 
	.A2(n807), 
	.A1(n806));
   SEN_ND2_S_6 U792 (.X(net17414), 
	.A2(net16360), 
	.A1(net16361));
   SEN_ND2_T_1P5 U793 (.X(net16327), 
	.A2(n608), 
	.A1(n554));
   SEN_MUXI2_S_2 U794 (.X(n608), 
	.S(B[8]), 
	.D1(n493), 
	.D0(n551));
   SEN_OAI211_3 U795 (.X(net3727), 
	.B2(net15965), 
	.B1(net15964), 
	.A2(net16412), 
	.A1(net15963));
   SEN_ND2_T_2 U796 (.X(n509), 
	.A2(B[16]), 
	.A1(n518));
   SEN_ND2B_V1_4 U797 (.X(net15912), 
	.B(net15916), 
	.A(net15915));
   SEN_NR2B_V1_2 U798 (.X(n526), 
	.B(n820), 
	.A(net17656));
   SEN_ND2_T_2 U799 (.X(n753), 
	.A2(n632), 
	.A1(n544));
   SEN_ND2_T_4 U800 (.X(n544), 
	.A2(n554), 
	.A1(n630));
   SEN_ND2_2 U801 (.X(n638), 
	.A2(n595), 
	.A1(net16476));
   SEN_MUXI2_DG_2 U802 (.X(n642), 
	.S(A[10]), 
	.D1(n683), 
	.D0(net16482));
   SEN_INV_2 U803 (.X(net16309), 
	.A(net16407));
   SEN_ND2_T_1 U804 (.X(n760), 
	.A2(n650), 
	.A1(n651));
   SEN_NR2_T_4 U805 (.X(n490), 
	.A2(n451), 
	.A1(net16691));
   SEN_EN2_S_3 U806 (.X(net15830), 
	.A2(n851), 
	.A1(n856));
   SEN_INV_S_4 U807 (.X(n415), 
	.A(Z[20]));
   SEN_OAI211_4 U808 (.X(Z[20]), 
	.B2(net15819), 
	.B1(net15818), 
	.A2(net16410), 
	.A1(net15817));
   SEN_ND2_T_1 U809 (.X(n646), 
	.A2(n642), 
	.A1(net17602));
   SEN_ND2_S_0P5 U810 (.X(net16190), 
	.A2(n685), 
	.A1(n686));
   SEN_INV_2 U811 (.X(n713), 
	.A(n685));
   SEN_ND2_G_1 U812 (.X(n685), 
	.A2(n684), 
	.A1(net17602));
   SEN_OAI21_T_4 U813 (.X(net3724), 
	.B(net16156), 
	.A2(net16155), 
	.A1(net16410));
   SEN_EN2_S_6 U814 (.X(net16155), 
	.A2(n706), 
	.A1(n710));
   SEN_OR3B_4 U815 (.X(n388), 
	.B2(Z[23]), 
	.B1(Z[21]), 
	.A(n381));
   SEN_ND2_T_2 U816 (.X(n650), 
	.A2(net17602), 
	.A1(n636));
   SEN_INV_S_2 U817 (.X(n636), 
	.A(n484));
   SEN_MUXI2_DG_0P75 U818 (.X(n562), 
	.S(B[27]), 
	.D1(n367), 
	.D0(n550));
   SEN_EO2_3 U819 (.X(net15963), 
	.A2(n531), 
	.A1(net15969));
   SEN_AOI21B_4 U820 (.X(n659), 
	.B(n652), 
	.A2(n653), 
	.A1(n654));
   SEN_EO2_1 U821 (.X(net17005), 
	.A2(net15790), 
	.A1(net15791));
   SEN_OAI21_2 U822 (.X(n735), 
	.B(n732), 
	.A2(n733), 
	.A1(n734));
   SEN_INV_3 U823 (.X(n737), 
	.A(n733));
   SEN_EO2_3 U824 (.X(n733), 
	.A2(n725), 
	.A1(n723));
   SEN_ND2_S_4 U825 (.X(net16336), 
	.A2(n602), 
	.A1(n553));
   SEN_EN2_5 U826 (.X(n785), 
	.A2(n788), 
	.A1(n789));
   SEN_INV_2 U827 (.X(n465), 
	.A(n748));
   SEN_INV_6 U828 (.X(n426), 
	.A(Z[15]));
   SEN_OAI211_8 U829 (.X(Z[15]), 
	.B2(net15904), 
	.B1(net15903), 
	.A2(net16410), 
	.A1(net15902));
   SEN_AOI21_6 U830 (.X(n675), 
	.B(n452), 
	.A2(n866), 
	.A1(n672));
   SEN_INV_S_4 U831 (.X(n810), 
	.A(n660));
   SEN_INV_0P65 U832 (.X(net16123), 
	.A(net16127));
   SEN_INV_1 U833 (.X(net16013), 
	.A(net15934));
   SEN_MUXI2_DG_3 U834 (.X(n592), 
	.S(B[17]), 
	.D1(n517), 
	.D0(n551));
   SEN_ND2_T_2 U835 (.X(net16337), 
	.A2(n603), 
	.A1(net16476));
   SEN_OR4B_4 U836 (.X(n706), 
	.B3(n692), 
	.B2(n693), 
	.B1(n694), 
	.A(n691));
   SEN_ND2_8 U837 (.X(net18157), 
	.A2(net17750), 
	.A1(net15916));
   SEN_NR2_8 U838 (.X(n512), 
	.A2(n491), 
	.A1(n513));
   SEN_EN2_S_2 U839 (.X(net15869), 
	.A2(n827), 
	.A1(n527));
   SEN_OAI211_3 U840 (.X(Z[10]), 
	.B2(net15871), 
	.B1(net15870), 
	.A2(net16410), 
	.A1(net15869));
   SEN_NR2_T_2 U841 (.X(n425), 
	.A2(Z[10]), 
	.A1(net3721));
   SEN_INV_S_6 U842 (.X(n814), 
	.A(n658));
   SEN_EN2_5 U843 (.X(n658), 
	.A2(n763), 
	.A1(n762));
   SEN_INV_1 U844 (.X(n821), 
	.A(n770));
   SEN_BUF_8 U845 (.X(net16501), 
	.A(INST[0]));
   SEN_EN2_3 U846 (.X(net16144), 
	.A2(n711), 
	.A1(net16999));
   SEN_OA21_2 U847 (.X(net17035), 
	.B(net16999), 
	.A2(net16084), 
	.A1(n442));
   SEN_EO2_G_2 U848 (.X(net16999), 
	.A2(n713), 
	.A1(n712));
   SEN_ND2_T_4 U849 (.X(net16288), 
	.A2(n554), 
	.A1(n627));
   SEN_OR3B_4 U850 (.X(n722), 
	.B2(n731), 
	.B1(n721), 
	.A(n720));
   SEN_ND2_6 U851 (.X(n398), 
	.A2(net17750), 
	.A1(net15916));
   SEN_EN2_S_1 U852 (.X(FLAGS[0]), 
	.A2(FLAGS[1]), 
	.A1(n702));
   SEN_AO2BB2_2 U853 (.X(FLAGS[1]), 
	.B2(n709), 
	.B1(n701), 
	.A2(n705), 
	.A1(n702));
   SEN_EO2_2 U854 (.X(n776), 
	.A2(n773), 
	.A1(n821));
   SEN_ND2_S_4 U855 (.X(net15902), 
	.A2(n460), 
	.A1(n459));
   SEN_ND3_T_4 U856 (.X(net16127), 
	.A3(net17005), 
	.A2(net16215), 
	.A1(n400));
   SEN_ND4B_4 U857 (.X(n400), 
	.B3(net15796), 
	.B2(net15795), 
	.B1(n398), 
	.A(net15798));
   SEN_OAOI211_2 U858 (.X(n773), 
	.C(net15882), 
	.B(n521), 
	.A2(n820), 
	.A1(net16023));
   SEN_ND2_4 U859 (.X(n813), 
	.A2(n492), 
	.A1(n765));
   SEN_ND2_4 U860 (.X(n457), 
	.A2(net17829), 
	.A1(n450));
   SEN_INV_1 U861 (.X(net17829), 
	.A(net15883));
   SEN_INV_S_1 U862 (.X(n723), 
	.A(n576));
   SEN_INV_S_1 U863 (.X(n470), 
	.A(n715));
   SEN_EO2_2 U864 (.X(n523), 
	.A2(net15888), 
	.A1(net15889));
   SEN_INV_S_1 U865 (.X(net16410), 
	.A(net16165));
   SEN_ND2_2 U866 (.X(n483), 
	.A2(A[13]), 
	.A1(n683));
   SEN_INV_2 U867 (.X(n698), 
	.A(n559));
   SEN_ND2_S_3 U868 (.X(n797), 
	.A2(n791), 
	.A1(n785));
   SEN_INV_3 U869 (.X(net17602), 
	.A(net17600));
   SEN_BUF_6 U870 (.X(net16495), 
	.A(INST[3]));
   SEN_INV_S_4 U871 (.X(net15967), 
	.A(net16301));
   SEN_INV_2 U872 (.X(n489), 
	.A(n488));
   SEN_INV_1 U873 (.X(net15889), 
	.A(net16326));
   SEN_EN2_0P5 U874 (.X(n378), 
	.A2(n811), 
	.A1(n810));
   SEN_INV_S_2 U875 (.X(n462), 
	.A(n879));
   SEN_INV_S_1 U876 (.X(n439), 
	.A(net16193));
   SEN_EO2_S_0P5 U877 (.X(n579), 
	.A2(n741), 
	.A1(n739));
   SEN_INV_S_1 U878 (.X(net16772), 
	.A(net16424));
   SEN_ND2_G_1 U879 (.X(n775), 
	.A2(n821), 
	.A1(net18219));
   SEN_EO2_G_2 U880 (.X(net17000), 
	.A2(net16069), 
	.A1(net16070));
   SEN_ND2_G_1 U881 (.X(net16134), 
	.A2(net16197), 
	.A1(net16196));
   SEN_EN2_1 U882 (.X(net16938), 
	.A2(net16134), 
	.A1(n439));
   SEN_INV_2 U883 (.X(net16412), 
	.A(net16165));
   SEN_EN2_1 U884 (.X(n535), 
	.A2(n728), 
	.A1(n730));
   SEN_ND2_S_3 U885 (.X(n406), 
	.A2(n408), 
	.A1(n407));
   SEN_ND2_G_1 U886 (.X(n473), 
	.A2(A[12]), 
	.A1(net16669));
   SEN_INV_S_1 U887 (.X(n541), 
	.A(B[13]));
   SEN_ND2_G_1 U888 (.X(n484), 
	.A2(n483), 
	.A1(n482));
   SEN_MUXI2_S_1 U889 (.X(n595), 
	.S(A[15]), 
	.D1(n683), 
	.D0(net16480));
   SEN_INV_6 U890 (.X(net16476), 
	.A(net16478));
   SEN_ND2_G_1 U891 (.X(n670), 
	.A2(n582), 
	.A1(n553));
   SEN_ND2_G_1 U892 (.X(n674), 
	.A2(n586), 
	.A1(net17602));
   SEN_INV_1 U893 (.X(net16220), 
	.A(net16074));
   SEN_ND2_G_1 U894 (.X(n681), 
	.A2(n679), 
	.A1(net17602));
   SEN_ND2_G_1 U895 (.X(n680), 
	.A2(n678), 
	.A1(n555));
   SEN_MUXI2_S_0P5 U896 (.X(n684), 
	.S(A[25]), 
	.D1(n549), 
	.D0(net16482));
   SEN_OAI21_S_2 U897 (.X(net16188), 
	.B(net16938), 
	.A2(net16143), 
	.A1(net17035));
   SEN_INV_S_3 U898 (.X(net15979), 
	.A(net16289));
   SEN_INV_S_1 U899 (.X(n546), 
	.A(B[3]));
   SEN_INV_3 U900 (.X(net16691), 
	.A(net15769));
   SEN_INV_1 U901 (.X(n861), 
	.A(n671));
   SEN_ND2_2 U902 (.X(n866), 
	.A2(n669), 
	.A1(n668));
   SEN_INV_S_1 U903 (.X(n712), 
	.A(n686));
   SEN_INV_S_1 U904 (.X(n728), 
	.A(n575));
   SEN_ND2_S_1 U905 (.X(n718), 
	.A2(n537), 
	.A1(n535));
   SEN_INV_3 U906 (.X(net16182), 
	.A(net16501));
   SEN_INV_3 U907 (.X(net16478), 
	.A(net17601));
   SEN_INV_2 U908 (.X(net17601), 
	.A(net17600));
   SEN_AOI21B_1 U909 (.X(n794), 
	.B(n791), 
	.A2(n792), 
	.A1(n793));
   SEN_ND2_T_1 U910 (.X(n469), 
	.A2(n467), 
	.A1(n771));
   SEN_INV_S_1 U911 (.X(n880), 
	.A(n662));
   SEN_ND2_G_1 U912 (.X(n463), 
	.A2(n879), 
	.A1(n539));
   SEN_ND2_G_1 U913 (.X(n464), 
	.A2(n462), 
	.A1(n461));
   SEN_ND2_T_1 U914 (.X(n840), 
	.A2(net18157), 
	.A1(n364));
   SEN_EN2_DG_1 U915 (.X(n537), 
	.A2(n889), 
	.A1(n886));
   SEN_OAI211_1 U916 (.X(Z[1]), 
	.B2(net15988), 
	.B1(net15987), 
	.A2(net16412), 
	.A1(net15986));
   SEN_EN2_1 U917 (.X(net15986), 
	.A2(n792), 
	.A1(n793));
   SEN_OAOI211_G_1 U918 (.X(net16018), 
	.C(n774), 
	.B(net16444), 
	.A2(A[8]), 
	.A1(B[8]));
   SEN_OA21_2 U919 (.X(net17804), 
	.B(n775), 
	.A2(net16412), 
	.A1(n776));
   SEN_OAI211_3 U920 (.X(net3748), 
	.B2(net16080), 
	.B1(net16079), 
	.A2(net16412), 
	.A1(net16078));
   SEN_ND2_2 U921 (.X(net16078), 
	.A2(n454), 
	.A1(n453));
   SEN_OAI211_3 U922 (.X(net3754), 
	.B2(n436), 
	.B1(n435), 
	.A2(n443), 
	.A1(n434));
   SEN_ND2B_6 U923 (.X(n395), 
	.B(n393), 
	.A(net16495));
   SEN_INV_S_2 U924 (.X(n424), 
	.A(Z[13]));
   SEN_ND3_S_0P5 U925 (.X(n815), 
	.A3(n834), 
	.A2(n813), 
	.A1(n814));
   SEN_AOAI211_8 U926 (.X(net16177), 
	.C(n390), 
	.B(net16501), 
	.A2(net16497), 
	.A1(n389));
   SEN_ND2_12 U927 (.X(net16669), 
	.A2(net17579), 
	.A1(net17349));
   SEN_OAOI211_G_1 U928 (.X(net15977), 
	.C(n795), 
	.B(net16444), 
	.A2(A[2]), 
	.A1(B[2]));
   SEN_INV_S_1 U929 (.X(n558), 
	.A(n704));
   SEN_ND2_G_4 U930 (.X(net16985), 
	.A2(n487), 
	.A1(n486));
   SEN_INV_S_3 U931 (.X(n418), 
	.A(net3748));
   SEN_ND2_S_2 U932 (.X(n449), 
	.A2(n446), 
	.A1(n440));
   SEN_ND2_2 U933 (.X(n434), 
	.A2(n449), 
	.A1(n448));
   SEN_ND2_S_0P5 U934 (.X(net16165), 
	.A2(n542), 
	.A1(n704));
   SEN_ND2_S_3 U935 (.X(n515), 
	.A2(n768), 
	.A1(n767));
   SEN_EO2_G_4 U936 (.X(net16028), 
	.A2(n530), 
	.A1(n766));
   SEN_INV_S_1 U937 (.X(net16774), 
	.A(net16691));
   SEN_ND2B_V1_3 U938 (.X(n632), 
	.B(n631), 
	.A(net16478));
   SEN_INV_S_3 U939 (.X(n550), 
	.A(n552));
   SEN_INV_S_8 U940 (.X(n551), 
	.A(n552));
   SEN_AN2_S_1 U941 (.X(n371), 
	.A2(n365), 
	.A1(n543));
   SEN_INV_S_1 U942 (.X(n555), 
	.A(n556));
   SEN_OR2_1 U943 (.X(n372), 
	.A2(B[31]), 
	.A1(A[31]));
   SEN_OR2_1 U944 (.X(n373), 
	.A2(B[29]), 
	.A1(A[29]));
   SEN_OR2_1 U945 (.X(n374), 
	.A2(B[30]), 
	.A1(A[30]));
   SEN_INV_S_1 U946 (.X(net16448), 
	.A(n359));
   SEN_NR2_0P8 U947 (.X(net15958), 
	.A2(net15960), 
	.A1(n399));
   SEN_MUXI2_S_1 U948 (.X(n584), 
	.S(A[20]), 
	.D1(n549), 
	.D0(net16480));
   SEN_NR3_T_0P5 U949 (.X(n862), 
	.A3(net16774), 
	.A2(n860), 
	.A1(n861));
   SEN_ND2B_S_4 U950 (.X(n700), 
	.B(net16400), 
	.A(net16179));
   SEN_MUXI2_DG_1 U951 (.X(n641), 
	.S(B[10]), 
	.D1(n494), 
	.D0(n551));
   SEN_ND2_T_6 U952 (.X(n392), 
	.A2(net16179), 
	.A1(net16361));
   SEN_ND2B_V1_1 U953 (.X(n695), 
	.B(net16497), 
	.A(A[31]));
   SEN_INV_0P65 U954 (.X(net15883), 
	.A(net15894));
   SEN_MUXI2_DG_1 U955 (.X(n613), 
	.S(A[5]), 
	.D1(net16669), 
	.D0(net16482));
   SEN_INV_4 U956 (.X(n393), 
	.A(net16499));
   SEN_INV_8 U957 (.X(net17656), 
	.A(net17655));
   SEN_INV_0P8 U958 (.X(n447), 
	.A(n440));
   SEN_EN2_S_3 U959 (.X(net15817), 
	.A2(n858), 
	.A1(n859));
   SEN_INV_1 U960 (.X(n853), 
	.A(n669));
   SEN_INV_S_8 U961 (.X(net17750), 
	.A(net17749));
   SEN_INV_S_3 U962 (.X(n627), 
	.A(n503));
   SEN_INV_4 U963 (.X(net16400), 
	.A(net16495));
   SEN_ND2_T_1P5 U964 (.X(n480), 
	.A2(n479), 
	.A1(n478));
   SEN_ND2_G_1 U965 (.X(n479), 
	.A2(n540), 
	.A1(n550));
   SEN_NR3_0P8 U966 (.X(net15939), 
	.A3(net16422), 
	.A2(net16723), 
	.A1(net15940));
   SEN_ND2_2 U967 (.X(net17427), 
	.A2(net15961), 
	.A1(n796));
   SEN_INV_4 U968 (.X(net17428), 
	.A(net17427));
   SEN_ND3_S_8 U969 (.X(n644), 
	.A3(net16985), 
	.A2(n834), 
	.A1(n814));
   SEN_INV_2 U970 (.X(n762), 
	.A(n656));
   SEN_NR3B_3 U971 (.X(n875), 
	.B2(net15798), 
	.B1(net15797), 
	.A(net15796));
   SEN_MUXI2_S_3 U972 (.X(n626), 
	.S(n545), 
	.D1(net16482), 
	.D0(n683));
   SEN_ND2_0P5 U973 (.X(net15996), 
	.A2(n524), 
	.A1(net18219));
   SEN_INV_S_1 U974 (.X(n859), 
	.A(n865));
   SEN_AO21_4 U975 (.X(n452), 
	.B(n865), 
	.A2(n866), 
	.A1(n845));
   SEN_ND2_S_0P5 U976 (.X(n863), 
	.A2(n848), 
	.A1(n866));
   SEN_ND2_1P5 U977 (.X(n848), 
	.A2(n665), 
	.A1(n664));
   SEN_INV_0P5 U978 (.X(n783), 
	.A(n780));
   SEN_INV_S_4 U979 (.X(n475), 
	.A(n749));
   SEN_INV_4 U980 (.X(net17190), 
	.A(net17189));
   SEN_ND2_T_2 U981 (.X(net15899), 
	.A2(n606), 
	.A1(n607));
   SEN_AN2_6 U982 (.X(net16968), 
	.A2(net16182), 
	.A1(net16400));
   SEN_NR2B_2 U983 (.X(n857), 
	.B(net15829), 
	.A(net18157));
   SEN_INV_S_0P5 U984 (.X(net15968), 
	.A(net16300));
   SEN_ND2_6 U985 (.X(n389), 
	.A2(n395), 
	.A1(n394));
   SEN_INV_2 U986 (.X(n763), 
	.A(n655));
   SEN_ND2_2 U987 (.X(n379), 
	.A2(net16182), 
	.A1(net16400));
   SEN_BUF_1 U988 (.X(n382), 
	.A(net16361));
   SEN_MUXI2_S_1 U989 (.X(n679), 
	.S(A[24]), 
	.D1(n549), 
	.D0(net16480));
   SEN_ND2_T_2 U990 (.X(n384), 
	.A2(n665), 
	.A1(n842));
   SEN_INV_S_3 U991 (.X(n383), 
	.A(n842));
   SEN_NR3B_3 U992 (.X(n870), 
	.B2(n863), 
	.B1(n864), 
	.A(net18157));
   SEN_OAI31_1 U993 (.X(n622), 
	.B(n621), 
	.A3(net16182), 
	.A2(net16309), 
	.A1(net16495));
   SEN_ND2_6 U994 (.X(net17749), 
	.A2(n751), 
	.A1(n645));
   SEN_MUXI2_DG_1 U995 (.X(n587), 
	.S(B[19]), 
	.D1(n368), 
	.D0(n550));
   SEN_INV_1 U996 (.X(n589), 
	.A(n866));
   SEN_INV_0P8 U997 (.X(net17564), 
	.A(net16499));
   SEN_ND2_4 U998 (.X(n765), 
	.A2(n516), 
	.A1(n515));
   SEN_ND2_G_1 U999 (.X(net15829), 
	.A2(n543), 
	.A1(n848));
   SEN_AO222_1 U1000 (.X(n386), 
	.C2(n724), 
	.C1(n725), 
	.B2(n373), 
	.B1(n359), 
	.A2(n737), 
	.A1(net18219));
   SEN_BUF_1 U1001 (.X(n387), 
	.A(n532));
   SEN_ND2_S_0P5 U1002 (.X(net15847), 
	.A2(n387), 
	.A1(net16434));
   SEN_OAI21_S_0P5 U1003 (.X(n849), 
	.B(n387), 
	.A2(n362), 
	.A1(n520));
   SEN_INV_S_3 U1004 (.X(n408), 
	.A(net3751));
   SEN_NR3_0P5 U1005 (.X(n808), 
	.A3(net16772), 
	.A2(n806), 
	.A1(n807));
   SEN_INV_8 U1006 (.X(net17349), 
	.A(n392));
   SEN_OR2_2 U1007 (.X(n548), 
	.A2(n537), 
	.A1(n885));
   SEN_INV_1 U1008 (.X(n458), 
	.A(n816));
   SEN_ND2_S_4 U1009 (.X(n749), 
	.A2(net16074), 
	.A1(n466));
   SEN_INV_1P5 U1010 (.X(n390), 
	.A(n391));
   SEN_INV_S_0P5 U1011 (.X(net18246), 
	.A(n382));
   SEN_ND2_S_0P5 U1012 (.X(net16201), 
	.A2(net17579), 
	.A1(net16361));
   SEN_ND2B_V1DG_2 U1013 (.X(net17579), 
	.B(net16968), 
	.A(A[31]));
   SEN_ND2_6 U1014 (.X(net16015), 
	.A2(net17428), 
	.A1(net17190));
   SEN_OAI221_4 U1015 (.X(net15897), 
	.C(net15953), 
	.B2(net16949), 
	.B1(n403), 
	.A2(net15961), 
	.A1(net16949));
   SEN_OR2_2 U1016 (.X(net17773), 
	.A2(n402), 
	.A1(n401));
   SEN_ND2_2 U1017 (.X(net15880), 
	.A2(net16325), 
	.A1(net16326));
   SEN_ND2_G_1 U1018 (.X(net15894), 
	.A2(net16327), 
	.A1(net16328));
   SEN_INV_4 U1019 (.X(n403), 
	.A(n399));
   SEN_ND2_3 U1020 (.X(net15946), 
	.A2(net16301), 
	.A1(net16300));
   SEN_NR2B_V1DG_1 U1021 (.X(net15956), 
	.B(net15960), 
	.A(net15942));
   SEN_BUF_1 U1022 (.X(net16701), 
	.A(net15942));
   SEN_NR4_3 U1023 (.X(FLAGS[2]), 
	.A4(net3724), 
	.A3(n406), 
	.A2(n405), 
	.A1(n404));
   SEN_ND3_S_4 U1024 (.X(n404), 
	.A3(n413), 
	.A2(n412), 
	.A1(n411));
   SEN_AN3B_4 U1025 (.X(n411), 
	.B2(n418), 
	.B1(n417), 
	.A(n419));
   SEN_NR2_S_4 U1026 (.X(n444), 
	.A2(Z[11]), 
	.A1(n427));
   SEN_ND3_S_4 U1027 (.X(n427), 
	.A3(n430), 
	.A2(n429), 
	.A1(n428));
   SEN_OAI211_3 U1028 (.X(net3715), 
	.B2(net16007), 
	.B1(net16006), 
	.A2(net16412), 
	.A1(net16005));
   SEN_NR4_6 U1029 (.X(n429), 
	.A4(net3733), 
	.A3(n431), 
	.A2(net3712), 
	.A1(net3730));
   SEN_OAI211_3 U1030 (.X(net3730), 
	.B2(net15938), 
	.B1(net15937), 
	.A2(net16412), 
	.A1(net15936));
   SEN_ND2_S_3 U1031 (.X(n431), 
	.A2(n433), 
	.A1(n432));
   SEN_INV_2 U1032 (.X(n432), 
	.A(net3727));
   SEN_OAI211_8 U1033 (.X(net3733), 
	.B2(net15949), 
	.B1(net15948), 
	.A2(net16412), 
	.A1(net15947));
   SEN_OAI211_4 U1034 (.X(Z[14]), 
	.B2(net16039), 
	.B1(net16038), 
	.A2(net16412), 
	.A1(net16037));
   SEN_NR2_S_4 U1035 (.X(n421), 
	.A2(Z[16]), 
	.A1(n423));
   SEN_ND3_S_4 U1036 (.X(n423), 
	.A3(n425), 
	.A2(n426), 
	.A1(n424));
   SEN_OAI211_2 U1037 (.X(Z[13]), 
	.B2(net15859), 
	.B1(net15858), 
	.A2(net16410), 
	.A1(net15857));
   SEN_OAI211_1 U1038 (.X(Z[16]), 
	.B2(net15921), 
	.B1(net15920), 
	.A2(net16410), 
	.A1(net15919));
   SEN_OAI211_3 U1039 (.X(Z[18]), 
	.B2(net15848), 
	.B1(net15847), 
	.A2(net16410), 
	.A1(net15846));
   SEN_ND2_T_6 U1040 (.X(Z[17]), 
	.A2(net15775), 
	.A1(net17713));
   SEN_ND2_2 U1041 (.X(n448), 
	.A2(net16938), 
	.A1(n447));
   SEN_INV_S_0P5 U1042 (.X(n446), 
	.A(net16938));
   SEN_INV_S_0P5 U1043 (.X(n443), 
	.A(net16165));
   SEN_ND2_S_0P5 U1044 (.X(n435), 
	.A2(net16938), 
	.A1(net18219));
   SEN_OA2BB2_0P5 U1045 (.X(n436), 
	.B2(net16448), 
	.B1(n438), 
	.A2(n437), 
	.A1(net16134));
   SEN_NR2_S_0P5 U1046 (.X(n437), 
	.A2(net16774), 
	.A1(n439));
   SEN_NR2_1 U1047 (.X(n438), 
	.A2(B[26]), 
	.A1(A[26]));
   SEN_INV_S_0P5 U1048 (.X(net16143), 
	.A(net16190));
   SEN_AO21B_6 U1049 (.X(net15794), 
	.B(net17000), 
	.A2(net16074), 
	.A1(net16073));
   SEN_NR2_T_2 U1050 (.X(net17788), 
	.A2(net16188), 
	.A1(net16127));
   SEN_ND2_6 U1051 (.X(n832), 
	.A2(n813), 
	.A1(net16057));
   SEN_AN2_3 U1052 (.X(n519), 
	.A2(n846), 
	.A1(net18157));
   SEN_INV_S_2 U1053 (.X(n467), 
	.A(n777));
   SEN_NR3_T_3 U1054 (.X(net16344), 
	.A3(n589), 
	.A2(net16220), 
	.A1(n747));
   SEN_INV_2 U1055 (.X(n747), 
	.A(n868));
   SEN_ND2_0P8 U1056 (.X(n508), 
	.A2(n507), 
	.A1(n551));
   SEN_INV_S_4 U1057 (.X(net17655), 
	.A(net15899));
   SEN_ND2B_4 U1058 (.X(n557), 
	.B(net16495), 
	.A(net16497));
   SEN_INV_S_6 U1059 (.X(net15797), 
	.A(net18157));
   SEN_ND2_2 U1060 (.X(n466), 
	.A2(net17799), 
	.A1(n465));
   SEN_INV_S_2 U1061 (.X(n829), 
	.A(n646));
   SEN_EO2_2 U1062 (.X(net15846), 
	.A2(n841), 
	.A1(n387));
   SEN_OAOI211_3 U1063 (.X(n841), 
	.C(n362), 
	.B(n520), 
	.A2(n839), 
	.A1(n840));
   SEN_ND2_2 U1064 (.X(n516), 
	.A2(n632), 
	.A1(n544));
   SEN_INV_2 U1065 (.X(n485), 
	.A(n818));
   SEN_ND2_S_2 U1066 (.X(n487), 
	.A2(n818), 
	.A1(n637));
   SEN_NR3_0P5 U1067 (.X(n819), 
	.A3(n817), 
	.A2(n818), 
	.A1(net16774));
   SEN_ND3_T_0P8 U1068 (.X(n583), 
	.A3(net16501), 
	.A2(net16497), 
	.A1(net16495));
   SEN_ND2_S_1P5 U1069 (.X(n655), 
	.A2(n634), 
	.A1(net17602));
   SEN_NR2_T_3 U1070 (.X(n497), 
	.A2(n379), 
	.A1(net17564));
   SEN_AN2_3 U1071 (.X(n525), 
	.A2(n846), 
	.A1(n365));
   SEN_INV_1 U1072 (.X(n856), 
	.A(n845));
   SEN_MUXI2_S_1 U1073 (.X(n582), 
	.S(B[20]), 
	.D1(n517), 
	.D0(n550));
   SEN_ND2B_V1_1 U1074 (.X(net16180), 
	.B(net16499), 
	.A(n583));
   SEN_MUXI2_S_2 U1075 (.X(n591), 
	.S(A[18]), 
	.D1(n683), 
	.D0(net16480));
   SEN_EN2_DG_4 U1076 (.X(net15927), 
	.A2(net15934), 
	.A1(n805));
   SEN_AOI21B_4 U1077 (.X(n727), 
	.B(n726), 
	.A2(n537), 
	.A1(n885));
   SEN_ND2_1P5 U1078 (.X(n669), 
	.A2(n588), 
	.A1(net16476));
   SEN_NR3_T_0P5 U1079 (.X(n798), 
	.A3(net15769), 
	.A2(net15968), 
	.A1(net15967));
   SEN_ND2_T_1P5 U1080 (.X(net16325), 
	.A2(n601), 
	.A1(net16476));
   SEN_INV_2 U1081 (.X(net15888), 
	.A(net16325));
   SEN_MUXI2_S_2 U1082 (.X(n601), 
	.S(A[9]), 
	.D1(n683), 
	.D0(net16480));
   SEN_MUX2_1 U1083 (.X(n625), 
	.S(n546), 
	.D1(n552), 
	.D0(n512));
   SEN_INV_S_1 U1084 (.X(net18219), 
	.A(net16440));
   SEN_OR2_DG_1 U1085 (.X(net16440), 
	.A2(n363), 
	.A1(n560));
   SEN_MUXI2_S_3 U1086 (.X(n614), 
	.S(B[1]), 
	.D1(n494), 
	.D0(n551));
   SEN_MUXI2_S_1 U1087 (.X(n600), 
	.S(B[9]), 
	.D1(n494), 
	.D0(n550));
   SEN_OAI21_S_0P5 U1088 (.X(n831), 
	.B(n759), 
	.A2(n832), 
	.A1(n534));
   SEN_MUXI2_DG_3 U1089 (.X(n630), 
	.S(B[11]), 
	.D1(n517), 
	.D0(n551));
   SEN_INV_1 U1090 (.X(net18184), 
	.A(net15969));
   SEN_INV_S_0P5 U1091 (.X(n805), 
	.A(n804));
   SEN_EO2_G_4 U1092 (.X(net15947), 
	.A2(n801), 
	.A1(net15953));
   SEN_INV_S_0P5 U1093 (.X(net15969), 
	.A(net15945));
   SEN_OAOI211_G_1 U1094 (.X(net15965), 
	.C(n798), 
	.B(net16444), 
	.A2(A[3]), 
	.A1(B[3]));
   SEN_EN2_S_2 U1095 (.X(net15936), 
	.A2(n803), 
	.A1(net16701));
   SEN_INV_S_0P5 U1096 (.X(net17799), 
	.A(net16073));
   SEN_MUXI2_S_1 U1097 (.X(n633), 
	.S(B[14]), 
	.D1(n518), 
	.D0(n551));
   SEN_ND2_T_1 U1098 (.X(net16326), 
	.A2(n600), 
	.A1(n553));
   SEN_EO2_S_3 U1099 (.X(n522), 
	.A2(n873), 
	.A1(n872));
   SEN_MUXI2_S_2 U1100 (.X(n588), 
	.S(A[19]), 
	.D1(n549), 
	.D0(net16480));
   SEN_ND2_3 U1101 (.X(n648), 
	.A2(n640), 
	.A1(net16476));
   SEN_ND3B_V1DG_1 U1102 (.X(n563), 
	.B2(net16497), 
	.B1(net16501), 
	.A(net16499));
   SEN_INV_1 U1103 (.X(net17573), 
	.A(net17572));
   SEN_NR3_T_0P5 U1104 (.X(n779), 
	.A3(net16772), 
	.A2(net16010), 
	.A1(net16009));
   SEN_ND2B_V1DG_2 U1105 (.X(net16360), 
	.B(net16968), 
	.A(A[31]));
   SEN_INV_2 U1106 (.X(n756), 
	.A(n648));
   SEN_ND2_S_3 U1107 (.X(net16298), 
	.A2(n613), 
	.A1(net16476));
   SEN_MUXI2_S_4 U1108 (.X(n619), 
	.S(A[0]), 
	.D1(n683), 
	.D0(net16482));
   SEN_INV_S_0P5 U1109 (.X(n766), 
	.A(n765));
   SEN_BUF_S_4 U1110 (.X(n492), 
	.A(n753));
   SEN_ND2_2 U1111 (.X(n665), 
	.A2(n591), 
	.A1(net16476));
   SEN_EO2_G_4 U1112 (.X(n527), 
	.A2(n829), 
	.A1(n828));
   SEN_EO2_G_2 U1113 (.X(net16037), 
	.A2(n761), 
	.A1(n814));
   SEN_INV_S_2 U1114 (.X(n789), 
	.A(n616));
   SEN_AN2_2 U1115 (.X(n530), 
	.A2(net15865), 
	.A1(n752));
   SEN_INV_0P65 U1116 (.X(n702), 
	.A(n706));
   SEN_MUXI2_S_3 U1117 (.X(n605), 
	.S(A[6]), 
	.D1(net16669), 
	.D0(net16482));
   SEN_ND2_2 U1118 (.X(net16077), 
	.A2(n638), 
	.A1(n637));
   SEN_ND2_T_3 U1119 (.X(n486), 
	.A2(n485), 
	.A1(n817));
   SEN_NR3_0P5 U1120 (.X(n697), 
	.A3(net16182), 
	.A2(n695), 
	.A1(net16499));
   SEN_INV_2 U1121 (.X(net16021), 
	.A(net16327));
   SEN_NR4B_4 U1122 (.X(n748), 
	.B3(n863), 
	.B2(n747), 
	.B1(n864), 
	.A(net18157));
   SEN_BUF_3 U1123 (.X(n543), 
	.A(n746));
   SEN_ND2_2 U1124 (.X(n455), 
	.A2(n663), 
	.A1(n880));
   SEN_ND2_2 U1125 (.X(n460), 
	.A2(net17816), 
	.A1(n458));
   SEN_INV_S_0P5 U1126 (.X(net17816), 
	.A(net16985));
   SEN_OAI31_3 U1127 (.X(n816), 
	.B(net15913), 
	.A3(net15912), 
	.A2(n815), 
	.A1(net15910));
   SEN_INV_S_1 U1128 (.X(n461), 
	.A(n539));
   SEN_ND2_2 U1129 (.X(net16005), 
	.A2(n469), 
	.A1(n468));
   SEN_INV_S_1 U1130 (.X(n471), 
	.A(A[12]));
   SEN_INV_S_3 U1131 (.X(n640), 
	.A(n474));
   SEN_ND2_S_4 U1132 (.X(n477), 
	.A2(n475), 
	.A1(net17760));
   SEN_INV_S_1 U1133 (.X(net17760), 
	.A(net17000));
   SEN_INV_2 U1134 (.X(n590), 
	.A(n480));
   SEN_ND2_G_1 U1135 (.X(n482), 
	.A2(n481), 
	.A1(net16482));
   SEN_INV_1 U1136 (.X(n481), 
	.A(A[13]));
   SEN_ND2_S_0P5 U1137 (.X(net15904), 
	.A2(net16985), 
	.A1(net16434));
   SEN_OAOI211_8 U1138 (.X(net15775), 
	.C(n882), 
	.B(net16444), 
	.A2(A[17]), 
	.A1(B[17]));
   SEN_AOAI211_3 U1139 (.X(n858), 
	.C(n866), 
	.B(n867), 
	.A2(n857), 
	.A1(n525));
   SEN_ND2_G_1 U1140 (.X(net15858), 
	.A2(n834), 
	.A1(net16434));
   SEN_INV_S_0P5 U1141 (.X(n809), 
	.A(n378));
   SEN_INV_0P8 U1142 (.X(net16474), 
	.A(net16478));
   SEN_INV_S_0P5 U1143 (.X(net17584), 
	.A(net16448));
   SEN_OAOI211_2 U1144 (.X(net15949), 
	.C(n802), 
	.B(net16444), 
	.A2(A[5]), 
	.A1(B[5]));
   SEN_OAOI211_2 U1145 (.X(net15929), 
	.C(n808), 
	.B(net16444), 
	.A2(A[6]), 
	.A1(B[6]));
   SEN_OAOI211_1 U1146 (.X(net15938), 
	.C(net15939), 
	.B(net16444), 
	.A2(A[4]), 
	.A1(B[4]));
   SEN_INV_S_0P5 U1147 (.X(n496), 
	.A(n492));
   SEN_ND2_G_1 U1148 (.X(n501), 
	.A2(n500), 
	.A1(n551));
   SEN_INV_1 U1149 (.X(n500), 
	.A(B[2]));
   SEN_INV_1 U1150 (.X(net16125), 
	.A(net16188));
   SEN_INV_1 U1151 (.X(n873), 
	.A(n674));
   SEN_INV_0P8 U1152 (.X(n744), 
	.A(n681));
   SEN_INV_S_1 U1153 (.X(n507), 
	.A(B[16]));
   SEN_OAOI211_1 U1154 (.X(net16146), 
	.C(n714), 
	.B(n359), 
	.A2(A[25]), 
	.A1(B[25]));
   SEN_NR2_S_0P5 U1155 (.X(n690), 
	.A2(n581), 
	.A1(n718));
   SEN_ND2B_1 U1156 (.X(n716), 
	.B(n535), 
	.A(n726));
   SEN_OAOI211_1 U1157 (.X(net16065), 
	.C(n750), 
	.B(net17584), 
	.A2(A[22]), 
	.A1(B[22]));
   SEN_NR3_0P5 U1158 (.X(n844), 
	.A3(net16774), 
	.A2(n842), 
	.A1(n843));
   SEN_NR3_0P5 U1159 (.X(n830), 
	.A3(net16772), 
	.A2(n828), 
	.A1(n829));
   SEN_MUXI2_S_0P5 U1160 (.X(n634), 
	.S(A[14]), 
	.D1(net16669), 
	.D0(net16482));
   SEN_NR3_T_0P5 U1161 (.X(n825), 
	.A3(net16772), 
	.A2(net15889), 
	.A1(net15888));
   SEN_INV_1 U1162 (.X(n710), 
	.A(n705));
   SEN_ND2_S_0P5 U1163 (.X(n657), 
	.A2(n655), 
	.A1(n656));
   SEN_ND2_S_0P5 U1164 (.X(n726), 
	.A2(n889), 
	.A1(n580));
   SEN_ND2_S_0P5 U1165 (.X(n701), 
	.A2(n699), 
	.A1(n555));
   SEN_OAOI211_0P5 U1166 (.X(net15859), 
	.C(n837), 
	.B(net16444), 
	.A2(A[13]), 
	.A1(B[13]));
   SEN_OAOI211_1 U1167 (.X(net16039), 
	.C(n764), 
	.B(net16444), 
	.A2(A[14]), 
	.A1(B[14]));
   SEN_INV_1 U1168 (.X(net16444), 
	.A(net16448));
   SEN_ND2_G_1 U1169 (.X(n581), 
	.A2(n742), 
	.A1(n737));
   SEN_NR3_0P5 U1170 (.X(n882), 
	.A3(net16774), 
	.A2(n880), 
	.A1(n881));
   SEN_NR3_0P5 U1171 (.X(n745), 
	.A3(net16772), 
	.A2(n743), 
	.A1(n744));
   SEN_ND3_S_0P5 U1172 (.X(n719), 
	.A3(net16190), 
	.A2(net16154), 
	.A1(net16153));
   SEN_AOI222_1 U1173 (.X(net16156), 
	.C2(n708), 
	.C1(n709), 
	.B2(n372), 
	.B1(net17584), 
	.A2(n710), 
	.A1(net16434));
   SEN_INV_S_1 U1174 (.X(net15791), 
	.A(net16191));
   SEN_OAOI211_1 U1175 (.X(net15800), 
	.C(n874), 
	.B(net17584), 
	.A2(A[21]), 
	.A1(B[21]));
   SEN_ND2_S_0P5 U1176 (.X(net15801), 
	.A2(n522), 
	.A1(net16434));
   SEN_OAOI211_1 U1177 (.X(net15832), 
	.C(n854), 
	.B(net17584), 
	.A2(A[19]), 
	.A1(B[19]));
   SEN_ND2_G_1 U1178 (.X(n741), 
	.A2(n573), 
	.A1(n574));
   SEN_OAOI211_1 U1179 (.X(net15819), 
	.C(n862), 
	.B(net17584), 
	.A2(A[20]), 
	.A1(B[20]));
   SEN_OAOI211_1 U1180 (.X(net16080), 
	.C(n745), 
	.B(n359), 
	.A2(A[24]), 
	.A1(B[24]));
   SEN_MUXI2_S_0P5 U1181 (.X(n676), 
	.S(B[23]), 
	.D1(n368), 
	.D0(n551));
   SEN_AN2_S_0P5 U1182 (.X(n520), 
	.A2(n838), 
	.A1(n533));
   SEN_INV_S_0P5 U1183 (.X(net16434), 
	.A(net16440));
   SEN_NR3_0P5 U1184 (.X(n877), 
	.A3(net15791), 
	.A2(net15790), 
	.A1(net16774));
   SEN_NR3_0P5 U1185 (.X(n874), 
	.A3(n872), 
	.A2(n873), 
	.A1(net16774));
   SEN_NR3_0P5 U1186 (.X(n750), 
	.A3(net16070), 
	.A2(net16069), 
	.A1(net16774));
   SEN_OA21B_1 U1187 (.X(n761), 
	.B(n529), 
	.A2(n528), 
	.A1(net15865));
   SEN_NR3_T_0P5 U1188 (.X(n714), 
	.A3(net16772), 
	.A2(n712), 
	.A1(n713));
   SEN_INV_1 U1189 (.X(n742), 
	.A(n579));
   SEN_INV_1 U1190 (.X(n734), 
	.A(n731));
   SEN_NR2_S_0P5 U1191 (.X(n724), 
	.A2(net16774), 
	.A1(n723));
   SEN_NR2_S_0P5 U1192 (.X(n740), 
	.A2(net16774), 
	.A1(n739));
   SEN_NR2_S_0P5 U1193 (.X(n708), 
	.A2(net16774), 
	.A1(n707));
   SEN_NR2_S_0P5 U1194 (.X(n888), 
	.A2(net16774), 
	.A1(n886));
   SEN_OAI21_S_0P5 U1195 (.X(n692), 
	.B(n578), 
	.A2(n579), 
	.A1(n732));
   SEN_NR2_S_0P5 U1196 (.X(n694), 
	.A2(n581), 
	.A1(n716));
   SEN_NR2_G_0P5 U1197 (.X(n693), 
	.A2(n581), 
	.A1(n717));
   SEN_NR2_S_0P5 U1198 (.X(n721), 
	.A2(n718), 
	.A1(n715));
   SEN_NR2_S_0P5 U1199 (.X(n729), 
	.A2(net16422), 
	.A1(n728));
   SEN_ND2_S_0P5 U1200 (.X(net16103), 
	.A2(n729), 
	.A1(n730));
   SEN_AOI22_0P5 U1201 (.X(net16104), 
	.B2(n538), 
	.B1(n359), 
	.A2(n535), 
	.A1(net18219));
   SEN_ND2_G_1 U1202 (.X(n868), 
	.A2(n671), 
	.A1(n670));
   SEN_ND2_S_0P5 U1203 (.X(net15762), 
	.A2(n537), 
	.A1(net18219));
   SEN_AN2_S_0P5 U1204 (.X(n536), 
	.A2(n542), 
	.A1(net16501));
   SEN_AN3B_0P5 U1205 (.X(n802), 
	.B2(net17648), 
	.B1(net16298), 
	.A(net16772));
   SEN_ND2_S_0P5 U1206 (.X(n732), 
	.A2(n725), 
	.A1(n576));
   SEN_ND2_S_0P5 U1207 (.X(n717), 
	.A2(n730), 
	.A1(n575));
   SEN_ND2_S_0P5 U1208 (.X(n578), 
	.A2(n741), 
	.A1(n577));
   SEN_INV_S_1 U1209 (.X(n872), 
	.A(n673));
   SEN_ND2_S_0P5 U1210 (.X(n715), 
	.A2(net16134), 
	.A1(net16193));
   SEN_OAOI211_1 U1211 (.X(net15997), 
	.C(n784), 
	.B(n359), 
	.A2(A[0]), 
	.A1(B[0]));
   SEN_OAOI211_1 U1212 (.X(net16007), 
	.C(n779), 
	.B(net16444), 
	.A2(A[7]), 
	.A1(B[7]));
   SEN_ND2_S_0P5 U1213 (.X(net16006), 
	.A2(n778), 
	.A1(net18219));
   SEN_OR3B_0P5 U1214 (.X(n709), 
	.B2(net16478), 
	.B1(n697), 
	.A(n696));
   SEN_ND2_S_0P5 U1215 (.X(net16066), 
	.A2(net17000), 
	.A1(net18219));
   SEN_ND2_S_0P5 U1216 (.X(net15818), 
	.A2(n859), 
	.A1(net16434));
   SEN_OAOI211_0P5 U1217 (.X(net15848), 
	.C(n844), 
	.B(net17584), 
	.A2(A[18]), 
	.A1(B[18]));
   SEN_ND2_S_0P5 U1218 (.X(net16145), 
	.A2(net16999), 
	.A1(n451));
   SEN_ND2_S_0P5 U1219 (.X(net15831), 
	.A2(n856), 
	.A1(net16434));
   SEN_OAOI211_1 U1220 (.X(net15786), 
	.C(n877), 
	.B(n359), 
	.A2(A[23]), 
	.A1(B[23]));
   SEN_ND2_S_0P5 U1221 (.X(net15787), 
	.A2(net17005), 
	.A1(net16434));
   SEN_OAOI211_1 U1222 (.X(net15988), 
	.C(n790), 
	.B(net17584), 
	.A2(A[1]), 
	.A1(B[1]));
   SEN_ND2_S_0P5 U1223 (.X(net15987), 
	.A2(n793), 
	.A1(net18219));
   SEN_ND2_S_0P5 U1224 (.X(net16079), 
	.A2(net16084), 
	.A1(net18219));
   SEN_ND2_S_0P5 U1225 (.X(net15976), 
	.A2(net15973), 
	.A1(net18219));
   SEN_OAOI211_0P5 U1226 (.X(net16030), 
	.C(n769), 
	.B(net16444), 
	.A2(A[11]), 
	.A1(B[11]));
   SEN_ND2_S_0P5 U1227 (.X(net16029), 
	.A2(n766), 
	.A1(net18219));
   SEN_ND2_S_0P5 U1228 (.X(net15920), 
	.A2(n809), 
	.A1(net16434));
   SEN_OAOI211_0P5 U1229 (.X(net15921), 
	.C(n812), 
	.B(net16444), 
	.A2(A[16]), 
	.A1(B[16]));
   SEN_ND2_S_0P5 U1230 (.X(net15870), 
	.A2(n527), 
	.A1(net16434));
   SEN_ND2_S_0P5 U1231 (.X(net15928), 
	.A2(n805), 
	.A1(net16434));
   SEN_MUXI2_S_0P5 U1232 (.X(n678), 
	.S(B[24]), 
	.D1(n511), 
	.D0(n550));
   SEN_INV_1 U1233 (.X(n545), 
	.A(A[3]));
   SEN_MUXI2_S_0P5 U1234 (.X(n565), 
	.S(A[27]), 
	.D1(net16201), 
	.D0(net16480));
   SEN_MUXI2_S_0P5 U1235 (.X(net16196), 
	.S(A[26]), 
	.D1(net16201), 
	.D0(net16482));
   SEN_INV_1 U1236 (.X(n540), 
	.A(B[18]));
   SEN_MUXI2_S_0P5 U1237 (.X(n586), 
	.S(A[21]), 
	.D1(n549), 
	.D0(net16480));
   SEN_MUXI2_S_0P5 U1238 (.X(n699), 
	.S(B[31]), 
	.D1(n367), 
	.D0(n550));
   SEN_INV_S_1 U1239 (.X(net16345), 
	.A(net15829));
   SEN_NR3_0P5 U1240 (.X(n790), 
	.A3(net16422), 
	.A2(n788), 
	.A1(n789));
   SEN_NR3_0P5 U1241 (.X(n757), 
	.A3(net16772), 
	.A2(n755), 
	.A1(n756));
   SEN_NR3_0P5 U1242 (.X(n795), 
	.A3(net16772), 
	.A2(net15980), 
	.A1(net15979));
   SEN_NR3_0P5 U1243 (.X(n774), 
	.A3(net16772), 
	.A2(net16021), 
	.A1(net16020));
   SEN_NR3_T_0P5 U1244 (.X(n854), 
	.A3(net16774), 
	.A2(n852), 
	.A1(n853));
   SEN_NR3_0P5 U1245 (.X(n764), 
	.A3(net16772), 
	.A2(n762), 
	.A1(n763));
   SEN_NR3_0P5 U1246 (.X(n837), 
	.A3(net16774), 
	.A2(n835), 
	.A1(n836));
   SEN_NR3_0P5 U1247 (.X(n769), 
	.A3(net16772), 
	.A2(n767), 
	.A1(n768));
   SEN_OR2_DG_1 U1248 (.X(n528), 
	.A2(n758), 
	.A1(n832));
   SEN_AO21B_1 U1249 (.X(n529), 
	.B(n760), 
	.A2(n831), 
	.A1(n834));
   SEN_ND2_G_1 U1250 (.X(n731), 
	.A2(n716), 
	.A1(n717));
   SEN_EO2_S_0P5 U1251 (.X(n705), 
	.A2(n707), 
	.A1(n709));
   SEN_OA2BB2_0P5 U1252 (.X(net15763), 
	.B2(net16448), 
	.B1(n887), 
	.A2(n888), 
	.A1(n889));
   SEN_INV_S_1 U1253 (.X(net15790), 
	.A(net16192));
   SEN_INV_S_1 U1254 (.X(net16069), 
	.A(net16222));
   SEN_INV_S_1 U1255 (.X(net16070), 
	.A(net16223));
   SEN_INV_S_1 U1256 (.X(n707), 
	.A(n701));
   SEN_INV_S_1 U1257 (.X(n739), 
	.A(n577));
   SEN_ND2_G_1 U1258 (.X(n889), 
	.A2(n564), 
	.A1(n565));
   SEN_INV_S_1 U1259 (.X(n26), 
	.A(n353));
   SEN_OAOI211_G_1 U1260 (.X(net15886), 
	.C(n825), 
	.B(net16444), 
	.A2(A[9]), 
	.A1(B[9]));
   SEN_ND2_S_0P5 U1261 (.X(net15885), 
	.A2(n523), 
	.A1(net16434));
   SEN_OAOI211_G_1 U1262 (.X(net15871), 
	.C(n830), 
	.B(net16444), 
	.A2(A[10]), 
	.A1(B[10]));
   SEN_ND2_G_1 U1263 (.X(net15964), 
	.A2(net15969), 
	.A1(net18219));
   SEN_OAOI211_G_1 U1264 (.X(net15903), 
	.C(n819), 
	.B(net16444), 
	.A2(A[15]), 
	.A1(B[15]));
   SEN_EN2_S_1 U1265 (.X(net15857), 
	.A2(n833), 
	.A1(n834));
   SEN_ND2_G_1 U1266 (.X(net16192), 
	.A2(n677), 
	.A1(net17602));
   SEN_INV_S_1 U1267 (.X(n28), 
	.A(n352));
   SEN_ND2_G_1 U1268 (.X(n730), 
	.A2(n567), 
	.A1(n568));
   SEN_MUXI2_S_0P5 U1269 (.X(n568), 
	.S(A[28]), 
	.D1(net16201), 
	.D0(net16480));
   SEN_INV_S_1 U1270 (.X(n24), 
	.A(n354));
   SEN_ND2_S_0P5 U1271 (.X(net16038), 
	.A2(n814), 
	.A1(net18219));
   SEN_OAOI211_G_1 U1272 (.X(net16053), 
	.C(n757), 
	.B(net17584), 
	.A2(A[12]), 
	.A1(B[12]));
   SEN_ND2_S_0P5 U1273 (.X(net16052), 
	.A2(n360), 
	.A1(net18219));
   SEN_ND2_G_1 U1274 (.X(n725), 
	.A2(n570), 
	.A1(n571));
   SEN_MUXI2_S_0P5 U1275 (.X(n571), 
	.S(A[29]), 
	.D1(net16201), 
	.D0(net16480));
   SEN_INV_S_1 U1276 (.X(n22), 
	.A(n355));
   SEN_MUXI2_S_0P5 U1277 (.X(n574), 
	.S(A[30]), 
	.D1(net16201), 
	.D0(net16480));
   SEN_INV_S_1 U1278 (.X(n20), 
	.A(n356));
   SEN_OR2_1 U1279 (.X(n538), 
	.A2(B[28]), 
	.A1(A[28]));
   SEN_NR2_1 U1280 (.X(n887), 
	.A2(B[27]), 
	.A1(A[27]));
   SEN_ND2_G_1 U1281 (.X(n671), 
	.A2(n584), 
	.A1(net17602));
   SEN_ND2_G_1 U1282 (.X(net16222), 
	.A2(n599), 
	.A1(net17602));
   SEN_MUXI2_S_0P5 U1283 (.X(n599), 
	.S(A[22]), 
	.D1(n549), 
	.D0(net16480));
   SEN_ND2_G_1 U1284 (.X(net16193), 
	.A2(n687), 
	.A1(n555));
   SEN_ND2_G_1 U1285 (.X(n576), 
	.A2(n569), 
	.A1(n553));
   SEN_MUXI2_S_0P5 U1286 (.X(n569), 
	.S(B[29]), 
	.D1(n367), 
	.D0(n550));
   SEN_ND2_G_1 U1287 (.X(n575), 
	.A2(n566), 
	.A1(n555));
   SEN_MUXI2_S_0P5 U1288 (.X(n566), 
	.S(B[28]), 
	.D1(n367), 
	.D0(n550));
   SEN_ND2_G_1 U1289 (.X(n577), 
	.A2(n572), 
	.A1(n553));
   SEN_MUXI2_S_0P5 U1290 (.X(n572), 
	.S(B[30]), 
	.D1(n367), 
	.D0(n550));
   SEN_ND2_G_1 U1291 (.X(n580), 
	.A2(n562), 
	.A1(n553));
   SEN_ND2_G_1 U1292 (.X(n686), 
	.A2(n682), 
	.A1(n555));
   SEN_ND2_G_1 U1293 (.X(n673), 
	.A2(n585), 
	.A1(n553));
   SEN_MUXI2_S_0P5 U1294 (.X(n585), 
	.S(B[21]), 
	.D1(n368), 
	.D0(n550));
   SEN_ND2_S_0P5 U1295 (.X(net16191), 
	.A2(n676), 
	.A1(n554));
   SEN_ND2_G_1 U1296 (.X(net16223), 
	.A2(n598), 
	.A1(n553));
   SEN_MUXI2_S_0P5 U1297 (.X(n598), 
	.S(B[22]), 
	.D1(n367), 
	.D0(n550));
   SEN_ND2B_S_0P5 U1298 (.X(n352), 
	.B(A[26]), 
	.A(net16499));
   SEN_ND2B_S_0P5 U1299 (.X(n353), 
	.B(A[27]), 
	.A(net16499));
   SEN_ND2B_S_0P5 U1300 (.X(n354), 
	.B(A[28]), 
	.A(net16499));
   SEN_ND2B_S_0P5 U1301 (.X(n355), 
	.B(A[29]), 
	.A(net16499));
   SEN_ND2B_S_0P5 U1302 (.X(n356), 
	.B(A[30]), 
	.A(net16499));
   SEN_NR3_0P5 U1303 (.X(n812), 
	.A3(net16772), 
	.A2(n810), 
	.A1(n811));
   SEN_MUXI2_S_1 U1304 (.X(net16197), 
	.S(n28), 
	.D1(n536), 
	.D0(n688));
   SEN_MUXI2_S_1 U1305 (.X(n573), 
	.S(n20), 
	.D1(n536), 
	.D0(n688));
   SEN_MUXI2_S_1 U1306 (.X(n570), 
	.S(n22), 
	.D1(n536), 
	.D0(n688));
   SEN_MUXI2_S_1 U1307 (.X(n567), 
	.S(n24), 
	.D1(n536), 
	.D0(n688));
   SEN_MUXI2_S_1 U1308 (.X(n564), 
	.S(n26), 
	.D1(n536), 
	.D0(n688));
   SEN_TIE0_1 U1309 (.X(\*Logic0* ));
   SEN_BUF_1 U1310 (.X(n539), 
	.A(n533));
   SEN_BUF_1 U1311 (.X(n542), 
	.A(n703));
   SEN_INV_S_0P5 U1312 (.X(net16178), 
	.A(net16179));
   SEN_BUF_1 U1313 (.X(net16723), 
	.A(net15941));
   SEN_MUXI2_S_0P5 U1314 (.X(n677), 
	.S(A[23]), 
	.D1(n549), 
	.D0(net16200));
   SEN_INV_S_0P5 U1315 (.X(n688), 
	.A(n583));
   SEN_ND3_S_0P5 U1316 (.X(n621), 
	.A3(n695), 
	.A2(net16968), 
	.A1(net16311));
   SEN_INV_S_1 U1317 (.X(net16424), 
	.A(net16774));
   SEN_OAI21_S_0P5 U1318 (.X(n696), 
	.B(A[31]), 
	.A2(net16178), 
	.A1(net18246));
   SEN_ND2_G_1 U1319 (.X(net15948), 
	.A2(net15953), 
	.A1(net16434));
   SEN_ND2_S_0P65 U1320 (.X(net15937), 
	.A2(net16701), 
	.A1(net16434));
   SEN_NR3_0P5 U1321 (.X(n784), 
	.A3(net15769), 
	.A2(n782), 
	.A1(n783));
   SEN_INV_S_1 U1322 (.X(net16422), 
	.A(net16424));
endmodule

