
module Alu ( Z, A, B, INST, FLAGS );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  output [3:0] FLAGS;
  wire   \*Logic0* , n20, n22, n24, n26, n28, n352, n353, n354, n355, n356,
         net3712, net3715, net3718, net3721, net3724, net3727, net3730,
         net3733, net3736, net3739, net3742, net3745, net3748, net3751,
         net3754, net3757, net15760, net15762, net15763, net15769, net15775,
         net15784, net15785, net15786, net15787, net15790, net15791, net15794,
         net15795, net15796, net15797, net15798, net15799, net15800, net15801,
         net15817, net15818, net15819, net15829, net15830, net15831, net15832,
         net15846, net15847, net15848, net15857, net15858, net15859, net15865,
         net15869, net15870, net15871, net15880, net15881, net15882, net15883,
         net15884, net15885, net15886, net15888, net15889, net15894, net15899,
         net15902, net15903, net15904, net15910, net15912, net15913, net15914,
         net15915, net15919, net15920, net15921, net15927, net15928, net15929,
         net15934, net15936, net15937, net15938, net15939, net15941, net15945,
         net15946, net15947, net15948, net15949, net15953, net15956, net15958,
         net15960, net15961, net15963, net15964, net15965, net15967, net15968,
         net15969, net15971, net15973, net15975, net15976, net15977, net15979,
         net15980, net15985, net15986, net15987, net15988, net15995, net15996,
         net15997, net16005, net16006, net16007, net16009, net16010, net16013,
         net16014, net16015, net16018, net16020, net16021, net16023, net16028,
         net16029, net16030, net16037, net16038, net16039, net16051, net16052,
         net16053, net16057, net16062, net16064, net16065, net16066, net16069,
         net16070, net16073, net16074, net16077, net16078, net16079, net16080,
         net16084, net16085, net16086, net16087, net16102, net16103, net16104,
         net16113, net16123, net16125, net16134, net16143, net16144, net16145,
         net16146, net16152, net16153, net16154, net16155, net16156, net16165,
         net16178, net16179, net16180, net16182, net16188, net16190, net16191,
         net16192, net16193, net16196, net16197, net16200, net16201, net16220,
         net16222, net16223, net16284, net16288, net16289, net16291, net16293,
         net16298, net16299, net16300, net16301, net16309, net16311, net16322,
         net16325, net16326, net16327, net16328, net16336, net16337, net16344,
         net16345, net16360, net16395, net16400, net16407, net16408, net16412,
         net16410, net16424, net16422, net16440, net16434, net16448, net16444,
         net16478, net16476, net16474, net16486, net16482, net16480, net16495,
         net16497, net16499, net16501, net16669, net16691, net16701, net16723,
         net16774, net16772, net16938, net16949, net16968, net16985, net16999,
         net17000, net17005, net17035, net17190, net17189, net17414, net17420,
         net17428, net17427, net17564, net17573, net17572, net17579, net17584,
         net17602, net17601, net17600, net17648, net17656, net17655, net17669,
         net17668, net17713, net17749, net17760, net17788, net17799, net17804,
         net17816, net17829, net17843, net18157, net18184, net18219, net18229,
         net18246, net16215, net16127, net17773, net17750, net17550, net16287,
         net16282, net16281, net15942, net15916, net15897, net17349, net16292,
         net15940, net16361, net16177, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889;
  assign FLAGS[3] = \*Logic0* ;
  assign Z[6] = net3712;
  assign Z[7] = net3715;
  assign Z[8] = net3718;
  assign Z[9] = net3721;
  assign Z[31] = net3724;
  assign Z[3] = net3727;
  assign Z[4] = net3730;
  assign Z[5] = net3733;
  assign Z[28] = net3736;
  assign Z[29] = net3739;
  assign Z[2] = net3742;
  assign Z[30] = net3745;
  assign Z[24] = net3748;
  assign Z[25] = net3751;
  assign Z[26] = net3754;
  assign Z[27] = net3757;

  SEN_ND2_3 U471 ( .A1(net16476), .A2(n619), .X(n780) );
  SEN_ND2_T_1 U472 ( .A1(n472), .A2(n473), .X(n474) );
  SEN_ND2_G_1 U473 ( .A1(net16482), .A2(n471), .X(n472) );
  SEN_ND2_S_2 U474 ( .A1(n641), .A2(n554), .X(n647) );
  SEN_AOAI211_6 U475 ( .A1(n543), .A2(n667), .B(n666), .C(n848), .X(n855) );
  SEN_OAI21_T_4 U476 ( .A1(n533), .A2(n847), .B(n532), .X(n666) );
  SEN_INV_AS_5 U477 ( .A(n838), .X(n667) );
  SEN_INV_1 U478 ( .A(n746), .X(n847) );
  SEN_ND2_2 U479 ( .A1(n662), .A2(n663), .X(n746) );
  SEN_NR2_T_5 U480 ( .A1(n772), .A2(net15882), .X(n610) );
  SEN_ND2_T_5 U481 ( .A1(n360), .A2(n527), .X(n643) );
  SEN_INV_S_3 U482 ( .A(n638), .X(n818) );
  SEN_INV_4 U483 ( .A(n855), .X(n672) );
  SEN_INV_3 U484 ( .A(n665), .X(n843) );
  SEN_ND2_G_1 U485 ( .A1(n649), .A2(n648), .X(n759) );
  SEN_OAI21_2 U486 ( .A1(n703), .A2(net16400), .B(n558), .X(n559) );
  SEN_INV_4 U487 ( .A(n557), .X(n703) );
  SEN_INV_4 U488 ( .A(n698), .X(n552) );
  SEN_ND2_1P5 U489 ( .A1(n690), .A2(n885), .X(n691) );
  SEN_ND2_S_6 U490 ( .A1(net15941), .A2(net15940), .X(n397) );
  SEN_OAI211_2 U491 ( .A1(net15884), .A2(net16410), .B1(net15885), .B2(
        net15886), .X(net3721) );
  SEN_EN2_S_2 U492 ( .A1(n523), .A2(n824), .X(net15884) );
  SEN_INV_S_6 U493 ( .A(n651), .X(n358) );
  SEN_ND2_T_4 U494 ( .A1(n635), .A2(n554), .X(n651) );
  SEN_INV_S_0P5 U495 ( .A(n651), .X(n835) );
  SEN_ND2_T_0P5 U496 ( .A1(net16085), .A2(net16152), .X(n454) );
  SEN_ND2_G_4 U497 ( .A1(n455), .A2(n456), .X(n533) );
  SEN_MUXI2_DG_2 U498 ( .D0(net16480), .D1(net16669), .S(A[17]), .X(n593) );
  SEN_INV_5 U499 ( .A(net16499), .X(net16311) );
  SEN_AN3_0P5 U500 ( .A1(net16311), .A2(n703), .A3(net16501), .X(n359) );
  SEN_OAI211_3 U501 ( .A1(net15785), .A2(net16410), .B1(net15786), .B2(
        net15787), .X(Z[23]) );
  SEN_OAI211_2 U502 ( .A1(net16144), .A2(net16410), .B1(net16145), .B2(
        net16146), .X(net3751) );
  SEN_OAI21B_4 U503 ( .A1(net16113), .A2(net16410), .B(n386), .X(net3739) );
  SEN_OR3_8 U504 ( .A1(net16281), .A2(net16282), .A3(net17773), .X(net15916)
         );
  SEN_ND2_2 U505 ( .A1(n463), .A2(n464), .X(n884) );
  SEN_INV_S_2 U506 ( .A(net16336), .X(net16010) );
  SEN_AOI31_4 U507 ( .A1(n737), .A2(n885), .A3(n736), .B(n735), .X(n738) );
  SEN_INV_1 U508 ( .A(net15897), .X(net15881) );
  SEN_OAI21_G_4 U509 ( .A1(n870), .A2(n869), .B(n868), .X(n871) );
  SEN_ND2_T_1 U510 ( .A1(n553), .A2(n587), .X(n668) );
  SEN_ND2_3 U511 ( .A1(net16474), .A2(n628), .X(net16289) );
  SEN_MUXI2_S_3 U512 ( .D0(net16482), .D1(n549), .S(A[2]), .X(n628) );
  SEN_INV_S_3 U513 ( .A(net16015), .X(net16281) );
  SEN_NR3_T_4 U514 ( .A1(net16284), .A2(net15985), .A3(net16287), .X(net16293)
         );
  SEN_ND2_S_6 U515 ( .A1(n505), .A2(n506), .X(net15985) );
  SEN_INV_6 U516 ( .A(n504), .X(n549) );
  SEN_INV_2 U517 ( .A(n758), .X(n834) );
  SEN_NR2_G_2 U518 ( .A1(n534), .A2(n758), .X(n653) );
  SEN_AOI211_G_5 U519 ( .A1(n771), .A2(n370), .B1(n610), .B2(n770), .X(n611)
         );
  SEN_INV_4 U520 ( .A(n369), .X(n370) );
  SEN_BUF_8 U521 ( .A(INST[1]), .X(net16499) );
  SEN_ND2_T_1 U522 ( .A1(net16501), .A2(net16499), .X(n704) );
  SEN_INV_1P25 U523 ( .A(n512), .X(n511) );
  SEN_ND2_2 U524 ( .A1(net16495), .A2(net16499), .X(n394) );
  SEN_INV_4 U525 ( .A(n620), .X(n782) );
  SEN_ND2_G_3 U526 ( .A1(n489), .A2(n561), .X(net15769) );
  SEN_ND2_S_3 U527 ( .A1(n791), .A2(n786), .X(n376) );
  SEN_ND2_1P5 U528 ( .A1(n787), .A2(n786), .X(n792) );
  SEN_NR2_T_1 U529 ( .A1(net16497), .A2(net16501), .X(n561) );
  SEN_INV_S_2 U530 ( .A(net3715), .X(n428) );
  SEN_ND2_T_2 U531 ( .A1(n554), .A2(n614), .X(n617) );
  SEN_MUXI2_S_3 U532 ( .D0(net16482), .D1(net16669), .S(A[4]), .X(n396) );
  SEN_INV_6 U533 ( .A(net16200), .X(net16486) );
  SEN_INV_3 U534 ( .A(Z[17]), .X(n381) );
  SEN_OAI211_4 U535 ( .A1(net15760), .A2(net16412), .B1(net15762), .B2(
        net15763), .X(net3757) );
  SEN_ND3_T_2 U536 ( .A1(n797), .A2(net15973), .A3(n796), .X(n799) );
  SEN_ND2_6 U537 ( .A1(n396), .A2(net16476), .X(net16292) );
  SEN_INV_5 U538 ( .A(n490), .X(n491) );
  SEN_INV_2 U539 ( .A(n512), .X(n518) );
  SEN_EN2_8 U540 ( .A1(n811), .A2(n810), .X(n878) );
  SEN_ND2_4 U541 ( .A1(n548), .A2(n547), .X(net15760) );
  SEN_INV_2 U542 ( .A(net15915), .X(n360) );
  SEN_INV_4 U543 ( .A(net15915), .X(net16057) );
  SEN_ND2_G_1 U544 ( .A1(net17648), .A2(net16298), .X(net16014) );
  SEN_INV_2 U545 ( .A(n544), .X(n767) );
  SEN_INV_S_1P5 U546 ( .A(n632), .X(n768) );
  SEN_ND2_S_6 U547 ( .A1(net15945), .A2(net15946), .X(net15961) );
  SEN_INV_4 U548 ( .A(net16292), .X(net15940) );
  SEN_EN2_S_4 U549 ( .A1(net16010), .A2(net16009), .X(n771) );
  SEN_ND2_T_2 U550 ( .A1(n508), .A2(n509), .X(n510) );
  SEN_AOI222_1 U551 ( .A1(n451), .A2(n742), .B1(net17584), .B2(n374), .C1(n741), .C2(n740), .X(net16087) );
  SEN_NR2_T_5 U552 ( .A1(n560), .A2(n499), .X(n451) );
  SEN_MUXI2_S_4 U553 ( .D0(net16480), .D1(net16669), .S(A[7]), .X(n603) );
  SEN_ND2_T_3 U554 ( .A1(net15916), .A2(net16062), .X(net15865) );
  SEN_INV_S_8 U555 ( .A(net16486), .X(net16480) );
  SEN_MUXI2_S_4 U556 ( .D0(n550), .D1(n493), .S(B[7]), .X(n602) );
  SEN_OAI211_3 U557 ( .A1(net16028), .A2(net16412), .B1(net16029), .B2(
        net16030), .X(Z[11]) );
  SEN_EN2_5 U558 ( .A1(net16021), .A2(net16020), .X(n770) );
  SEN_ND2_T_6 U559 ( .A1(n878), .A2(net17669), .X(n838) );
  SEN_INV_S_3 U560 ( .A(net15784), .X(net17668) );
  SEN_ND2_3 U561 ( .A1(n660), .A2(n361), .X(net15784) );
  SEN_ND2_T_4 U562 ( .A1(n554), .A2(n604), .X(n607) );
  SEN_ND2_T_5 U563 ( .A1(n804), .A2(net17656), .X(n772) );
  SEN_ND2_S_1P5 U564 ( .A1(n537), .A2(n885), .X(n547) );
  SEN_INV_AS_10 U565 ( .A(net16486), .X(net16482) );
  SEN_INV_3 U566 ( .A(n649), .X(n755) );
  SEN_ND2_T_2 U567 ( .A1(n662), .A2(n881), .X(n456) );
  SEN_INV_1P25 U568 ( .A(n663), .X(n881) );
  SEN_ND2_S_0P5 U569 ( .A1(net16434), .A2(n539), .X(n883) );
  SEN_OA21_4 U570 ( .A1(n884), .A2(net16410), .B(n883), .X(net17713) );
  SEN_OAI21_2 U571 ( .A1(n521), .A2(net15882), .B(n821), .X(n822) );
  SEN_NR2_S_1 U572 ( .A1(net15881), .A2(net15882), .X(n823) );
  SEN_NR3_T_0P8 U573 ( .A1(net15881), .A2(net15882), .A3(net15883), .X(n826)
         );
  SEN_ND3_T_1 U574 ( .A1(net15880), .A2(net15894), .A3(n370), .X(n401) );
  SEN_INV_5 U575 ( .A(n370), .X(net15882) );
  SEN_ND2_T_2 U576 ( .A1(net16336), .A2(net16337), .X(net16322) );
  SEN_MUXI2_S_4 U577 ( .D0(n551), .D1(n493), .S(B[4]), .X(n629) );
  SEN_INV_5 U578 ( .A(n512), .X(n493) );
  SEN_OA21_4 U579 ( .A1(n758), .A2(n759), .B(n760), .X(n652) );
  SEN_ND2_G_0P65 U580 ( .A1(n680), .A2(n681), .X(net16153) );
  SEN_INV_S_2 U581 ( .A(n680), .X(n743) );
  SEN_ND2_G_2 U582 ( .A1(net16311), .A2(net16495), .X(n488) );
  SEN_ND2_G_1 U583 ( .A1(net17602), .A2(n597), .X(n361) );
  SEN_ND2_2 U584 ( .A1(net17602), .A2(n597), .X(n661) );
  SEN_MUXI2_S_2 U585 ( .D0(net16480), .D1(net16669), .S(A[16]), .X(n597) );
  SEN_INV_2 U586 ( .A(net15985), .X(net15973) );
  SEN_ND2_T_4 U587 ( .A1(n787), .A2(n377), .X(n796) );
  SEN_AN2_DG_2 U588 ( .A1(net16291), .A2(net16292), .X(net16949) );
  SEN_BUF_1 U589 ( .A(n847), .X(n362) );
  SEN_INV_4 U590 ( .A(n606), .X(n807) );
  SEN_ND2_T_4 U591 ( .A1(net17602), .A2(n605), .X(n606) );
  SEN_INV_S_6 U592 ( .A(n607), .X(n806) );
  SEN_INV_8 U593 ( .A(n504), .X(n683) );
  SEN_NR2B_V1_8 U594 ( .A(net16179), .B(net17414), .X(n504) );
  SEN_EO2_6 U595 ( .A1(net16300), .A2(net15967), .X(net15945) );
  SEN_ND2_S_2 U596 ( .A1(net16985), .A2(n816), .X(n459) );
  SEN_ND2_G_1 U597 ( .A1(net16311), .A2(net16408), .X(net16407) );
  SEN_INV_2 U598 ( .A(n622), .X(n781) );
  SEN_NR2_S_4 U599 ( .A1(n780), .A2(n781), .X(n623) );
  SEN_NR3_T_6 U600 ( .A1(n388), .A2(net3757), .A3(n414), .X(n412) );
  SEN_INV_3 U601 ( .A(n611), .X(n450) );
  SEN_EN2_S_6 U602 ( .A1(n737), .A2(n722), .X(net16113) );
  SEN_OAI211_3 U603 ( .A1(net16123), .A2(n719), .B1(net16125), .B2(n736), .X(
        n720) );
  SEN_ND2_T_2 U604 ( .A1(net16476), .A2(n615), .X(n616) );
  SEN_INV_3 U605 ( .A(n376), .X(n377) );
  SEN_ND2_2 U606 ( .A1(n617), .A2(n616), .X(n791) );
  SEN_ND2_S_4 U607 ( .A1(n409), .A2(n410), .X(n405) );
  SEN_INV_2P5 U608 ( .A(n661), .X(n811) );
  SEN_INV_4 U609 ( .A(n556), .X(n553) );
  SEN_ND2_S_4 U610 ( .A1(n592), .A2(n553), .X(n662) );
  SEN_ND2_T_2 U611 ( .A1(n553), .A2(n590), .X(n664) );
  SEN_ND2_S_4 U612 ( .A1(n415), .A2(n416), .X(n414) );
  SEN_MUXI2_DG_2 U613 ( .D0(net16482), .D1(net16669), .S(A[11]), .X(n631) );
  SEN_OAI211_3 U614 ( .A1(net15830), .A2(net16410), .B1(net15831), .B2(
        net15832), .X(Z[19]) );
  SEN_ND2_S_3 U615 ( .A1(n554), .A2(n612), .X(net16299) );
  SEN_MUXI2_DG_3 U616 ( .D0(n551), .D1(n518), .S(B[5]), .X(n612) );
  SEN_INV_S_4 U617 ( .A(n498), .X(n499) );
  SEN_ND2B_V1_2 U618 ( .A(net16501), .B(net16495), .X(n560) );
  SEN_OAI21_5 U619 ( .A1(net16086), .A2(net16410), .B(net16087), .X(net3745)
         );
  SEN_ND2_6 U620 ( .A1(n384), .A2(n385), .X(n532) );
  SEN_NR2_S_3 U621 ( .A1(net16311), .A2(net16497), .X(n498) );
  SEN_ND2_T_4 U622 ( .A1(n626), .A2(net17602), .X(net16301) );
  SEN_ND2_S_0P5 U623 ( .A1(n855), .A2(n856), .X(n867) );
  SEN_OAI21_S_1P5 U624 ( .A1(n531), .A2(net18184), .B(net15946), .X(n803) );
  SEN_INV_4 U625 ( .A(n650), .X(n836) );
  SEN_ND3_S_8 U626 ( .A1(n420), .A2(n421), .A3(n422), .X(n419) );
  SEN_ND2_T_2 U627 ( .A1(n518), .A2(B[18]), .X(n478) );
  SEN_OAI21_G_2 U628 ( .A1(n875), .A2(net15794), .B(net15795), .X(n876) );
  SEN_INV_S_1 U629 ( .A(net15961), .X(net15960) );
  SEN_ND2_3 U630 ( .A1(net16288), .A2(net17420), .X(n506) );
  SEN_INV_4 U631 ( .A(net15979), .X(net17420) );
  SEN_ND2_T_2 U632 ( .A1(net16476), .A2(n593), .X(n663) );
  SEN_AN3_4 U633 ( .A1(net17564), .A2(n703), .A3(net16501), .X(net18229) );
  SEN_ND2_S_6 U634 ( .A1(n846), .A2(n371), .X(n864) );
  SEN_INV_AS_10 U635 ( .A(n839), .X(n846) );
  SEN_EO2_1 U636 ( .A1(n809), .A2(n519), .X(net15919) );
  SEN_OAI21_5 U637 ( .A1(n675), .A2(n747), .B(n522), .X(net16073) );
  SEN_INV_S_4 U638 ( .A(net16291), .X(net15941) );
  SEN_EN2_S_3 U639 ( .A1(n860), .A2(n861), .X(n865) );
  SEN_INV_S_3 U640 ( .A(n670), .X(n860) );
  SEN_INV_2 U641 ( .A(n799), .X(n800) );
  SEN_ND2_4 U642 ( .A1(n476), .A2(n477), .X(net16064) );
  SEN_INV_S_6 U643 ( .A(net3745), .X(n413) );
  SEN_ND2_S_4 U644 ( .A1(n618), .A2(n554), .X(n620) );
  SEN_INV_S_2 U645 ( .A(n580), .X(n886) );
  SEN_BUF_1 U646 ( .A(n499), .X(n363) );
  SEN_EN2_3 U647 ( .A1(n522), .A2(n871), .X(net15799) );
  SEN_NR3_T_3 U648 ( .A1(net3742), .A2(Z[0]), .A3(Z[1]), .X(n433) );
  SEN_OAI211_1 U649 ( .A1(net15995), .A2(net16412), .B1(net15996), .B2(
        net15997), .X(Z[0]) );
  SEN_EO2_1 U650 ( .A1(n782), .A2(n783), .X(n524) );
  SEN_INV_1P25 U651 ( .A(net16497), .X(net16408) );
  SEN_ND2_T_4 U652 ( .A1(net16501), .A2(net16309), .X(net16179) );
  SEN_INV_10 U653 ( .A(n556), .X(n554) );
  SEN_INV_S_8 U654 ( .A(n700), .X(n556) );
  SEN_INV_0P5 U655 ( .A(n771), .X(n778) );
  SEN_ND2_4 U656 ( .A1(net16293), .A2(n797), .X(net17189) );
  SEN_AOI211_G_2 U657 ( .A1(n800), .A2(net15956), .B1(net16949), .B2(net15958), 
        .X(n801) );
  SEN_AN2_S_1P5 U658 ( .A1(n492), .A2(n752), .X(n534) );
  SEN_ND2_T_1 U659 ( .A1(n749), .A2(net17000), .X(n476) );
  SEN_ND2_3 U660 ( .A1(n563), .A2(net16395), .X(net16200) );
  SEN_EO2_DG_1 U661 ( .A1(n781), .A2(n524), .X(net15995) );
  SEN_OAOI211_4 U662 ( .A1(n441), .A2(n442), .B(net17035), .C(net16143), .X(
        n440) );
  SEN_INV_1 U663 ( .A(net16337), .X(net16009) );
  SEN_MUXI2_S_6 U664 ( .D0(n551), .D1(n493), .S(B[6]), .X(n604) );
  SEN_OAI211_4 U665 ( .A1(net16051), .A2(net16412), .B1(net16052), .B2(
        net16053), .X(Z[12]) );
  SEN_INV_2P5 U666 ( .A(n512), .X(n494) );
  SEN_ND2_T_3 U667 ( .A1(net16127), .A2(net16154), .X(n441) );
  SEN_INV_0P65 U668 ( .A(n512), .X(n368) );
  SEN_INV_2 U669 ( .A(n512), .X(n517) );
  SEN_NR3_T_6 U670 ( .A1(Z[12]), .A2(n445), .A3(Z[14]), .X(n420) );
  SEN_ND2_S_2 U671 ( .A1(net16015), .A2(net16014), .X(n820) );
  SEN_AN2_S_1 U672 ( .A1(n778), .A2(n375), .X(n521) );
  SEN_ND2_S_1 U673 ( .A1(n804), .A2(net17656), .X(n375) );
  SEN_ND2B_V1_4 U674 ( .A(n556), .B(n629), .X(net16291) );
  SEN_INV_3 U675 ( .A(net15897), .X(net16282) );
  SEN_ND2_2 U676 ( .A1(n494), .A2(B[2]), .X(n502) );
  SEN_ND2_T_2 U677 ( .A1(n502), .A2(n501), .X(n503) );
  SEN_AOAI211_2 U678 ( .A1(n526), .A2(n823), .B(n822), .C(net15894), .X(n824)
         );
  SEN_ND2_2 U679 ( .A1(n673), .A2(n674), .X(net16074) );
  SEN_EN2_S_4 U680 ( .A1(n755), .A2(n756), .X(net15915) );
  SEN_INV_3 U681 ( .A(n832), .X(n654) );
  SEN_ND2_G_1 U682 ( .A1(net16191), .A2(net16192), .X(net16154) );
  SEN_ND2_T_2 U683 ( .A1(net16125), .A2(n719), .X(n689) );
  SEN_ND2_T_4 U684 ( .A1(n383), .A2(n843), .X(n385) );
  SEN_INV_S_4 U685 ( .A(n664), .X(n842) );
  SEN_ND2_T_1 U686 ( .A1(n554), .A2(n633), .X(n656) );
  SEN_ND2_T_2 U687 ( .A1(n554), .A2(n639), .X(n649) );
  SEN_ND2_S_4 U688 ( .A1(n625), .A2(n554), .X(net16300) );
  SEN_AO21B_1 U689 ( .A1(n867), .A2(n866), .B(n859), .X(n869) );
  SEN_ND2_2 U690 ( .A1(net16291), .A2(net16292), .X(net17550) );
  SEN_ND2_6 U691 ( .A1(n397), .A2(net17550), .X(net16287) );
  SEN_INV_1P25 U692 ( .A(n647), .X(n828) );
  SEN_ND2_T_1 U693 ( .A1(n647), .A2(n646), .X(n752) );
  SEN_EN2_S_3 U694 ( .A1(net17005), .A2(n876), .X(net15785) );
  SEN_INV_S_3 U695 ( .A(n617), .X(n788) );
  SEN_INV_4 U696 ( .A(net16284), .X(net15953) );
  SEN_INV_S_6 U697 ( .A(net3739), .X(n410) );
  SEN_INV_0P8 U698 ( .A(n718), .X(n736) );
  SEN_INV_3 U699 ( .A(n444), .X(n445) );
  SEN_INV_S_2 U700 ( .A(n785), .X(n793) );
  SEN_OAI211_4 U701 ( .A1(net15927), .A2(net16412), .B1(net15928), .B2(
        net15929), .X(net3712) );
  SEN_ND2_S_4 U702 ( .A1(net17804), .A2(net16018), .X(net3718) );
  SEN_ND2_8 U703 ( .A1(n380), .A2(net15880), .X(n751) );
  SEN_INV_2 U704 ( .A(net16328), .X(net16020) );
  SEN_ND2_T_2 U705 ( .A1(n609), .A2(net17602), .X(net16328) );
  SEN_MUXI2_DG_2 U706 ( .D0(net16482), .D1(n683), .S(A[8]), .X(n609) );
  SEN_AO21B_2 U707 ( .A1(n441), .A2(net16084), .B(net16153), .X(n711) );
  SEN_EN2_3 U708 ( .A1(n743), .A2(n744), .X(net16152) );
  SEN_INV_2P5 U709 ( .A(net16152), .X(net16084) );
  SEN_INV_6 U710 ( .A(net16177), .X(net16361) );
  SEN_INV_S_4 U711 ( .A(net3718), .X(n430) );
  SEN_ND2_S_2 U712 ( .A1(net16084), .A2(net17843), .X(n453) );
  SEN_INV_S_4 U713 ( .A(n637), .X(n817) );
  SEN_ND2_S_3 U714 ( .A1(n555), .A2(n594), .X(n637) );
  SEN_INV_6 U715 ( .A(net16287), .X(net15942) );
  SEN_INV_S_0P5 U716 ( .A(net17668), .X(n364) );
  SEN_INV_S_0P5 U717 ( .A(net17668), .X(n365) );
  SEN_INV_4 U718 ( .A(net17668), .X(net17669) );
  SEN_INV_S_3 U719 ( .A(net16322), .X(n369) );
  SEN_NR2_T_1P5 U720 ( .A1(n530), .A2(n765), .X(n495) );
  SEN_AOAI211_G_2 U721 ( .A1(n526), .A2(n826), .B(n380), .C(net15880), .X(n827) );
  SEN_ND2_T_6 U722 ( .A1(n457), .A2(n523), .X(n380) );
  SEN_EO2_S_3 U723 ( .A1(n742), .A2(n738), .X(net16086) );
  SEN_ND2_T_6 U724 ( .A1(n514), .A2(n689), .X(n885) );
  SEN_NR2_T_4 U725 ( .A1(net17788), .A2(n470), .X(n514) );
  SEN_MUXI2_S_1 U726 ( .D0(n551), .D1(n367), .S(B[26]), .X(n687) );
  SEN_MUX2_DG_1 U727 ( .D0(n512), .D1(n552), .S(n541), .X(n635) );
  SEN_MUXI2_S_3 U728 ( .D0(net16482), .D1(n683), .S(A[1]), .X(n615) );
  SEN_OAI211_3 U729 ( .A1(net15799), .A2(net16410), .B1(net15800), .B2(
        net15801), .X(Z[21]) );
  SEN_OR2_5 U730 ( .A1(net18229), .A2(n497), .X(n513) );
  SEN_INV_0P65 U731 ( .A(net15914), .X(net15913) );
  SEN_ND2_T_8 U732 ( .A1(net15796), .A2(net16077), .X(n839) );
  SEN_ND2_8 U733 ( .A1(net15914), .A2(net16985), .X(net15796) );
  SEN_EO2_G_2 U734 ( .A1(net15973), .A2(n794), .X(net15975) );
  SEN_EN2_3 U735 ( .A1(n852), .A2(n853), .X(n845) );
  SEN_INV_S_2 U736 ( .A(n668), .X(n852) );
  SEN_ND2_6 U737 ( .A1(n553), .A2(n596), .X(n660) );
  SEN_INV_3 U738 ( .A(net3754), .X(n407) );
  SEN_INV_4 U739 ( .A(n510), .X(n596) );
  SEN_EN2_6 U740 ( .A1(net17648), .A2(net16298), .X(net16284) );
  SEN_ND3_T_1P5 U741 ( .A1(n389), .A2(net16968), .A3(net17573), .X(net16395)
         );
  SEN_MUXI2_S_3 U742 ( .D0(n551), .D1(n517), .S(B[12]), .X(n639) );
  SEN_INV_0P8 U743 ( .A(net16085), .X(net17843) );
  SEN_EO2_5 U744 ( .A1(n623), .A2(n624), .X(n787) );
  SEN_OAI21_S_3 U745 ( .A1(n519), .A2(n378), .B(n364), .X(n879) );
  SEN_NR2_2 U746 ( .A1(net15797), .A2(n362), .X(n850) );
  SEN_INV_S_4 U747 ( .A(Z[22]), .X(n417) );
  SEN_EN2_3 U748 ( .A1(n360), .A2(n754), .X(net16051) );
  SEN_OAI211_4 U749 ( .A1(net16064), .A2(net16412), .B1(net16065), .B2(
        net16066), .X(Z[22]) );
  SEN_OR2_2P5 U750 ( .A1(n495), .A2(n496), .X(n754) );
  SEN_INV_S_2 U751 ( .A(n494), .X(n366) );
  SEN_INV_3 U752 ( .A(n366), .X(n367) );
  SEN_ND2_1P5 U753 ( .A1(n780), .A2(n620), .X(n786) );
  SEN_ND2_S_4 U754 ( .A1(n782), .A2(n622), .X(n624) );
  SEN_AOAI211_3 U755 ( .A1(n525), .A2(n850), .B(n849), .C(n848), .X(n851) );
  SEN_ND3_T_1 U756 ( .A1(net15897), .A2(net16015), .A3(net16014), .X(net15934)
         );
  SEN_OAI21_S_3 U757 ( .A1(net16013), .A2(n804), .B(net17656), .X(n777) );
  SEN_INV_S_6 U758 ( .A(net3736), .X(n409) );
  SEN_OAI211_8 U759 ( .A1(net16102), .A2(n443), .B1(net16103), .B2(net16104), 
        .X(net3736) );
  SEN_EO2_G_8 U760 ( .A1(n535), .A2(n727), .X(net16102) );
  SEN_ND2_T_1 U761 ( .A1(net16497), .A2(A[31]), .X(net17572) );
  SEN_NR2_G_1 U762 ( .A1(net16497), .A2(net16495), .X(n391) );
  SEN_BUF_8 U763 ( .A(INST[2]), .X(net16497) );
  SEN_ND2_2 U764 ( .A1(net16288), .A2(net16289), .X(net15971) );
  SEN_INV_2 U765 ( .A(n441), .X(net16085) );
  SEN_AO21B_6 U766 ( .A1(net15971), .A2(net15946), .B(net15942), .X(n399) );
  SEN_AN2_3 U767 ( .A1(net15971), .A2(n799), .X(n531) );
  SEN_INV_S_4 U768 ( .A(Z[19]), .X(n416) );
  SEN_INV_S_4 U769 ( .A(Z[18]), .X(n422) );
  SEN_ND2_2 U770 ( .A1(net15980), .A2(net15979), .X(n505) );
  SEN_INV_S_2 U771 ( .A(net16288), .X(net15980) );
  SEN_INV_S_4 U772 ( .A(net15910), .X(net16062) );
  SEN_ND2_T_3 U773 ( .A1(n751), .A2(n527), .X(net15910) );
  SEN_BUF_S_6 U774 ( .A(net16299), .X(net17648) );
  SEN_ND2_S_1 U775 ( .A1(n778), .A2(n777), .X(n468) );
  SEN_INV_S_2 U776 ( .A(net16180), .X(net17600) );
  SEN_MUXI2_DG_3 U777 ( .D0(n551), .D1(n511), .S(B[0]), .X(n618) );
  SEN_OAI211_3 U778 ( .A1(net15975), .A2(net16412), .B1(net15976), .B2(
        net15977), .X(net3742) );
  SEN_MUXI2_S_0P5 U779 ( .D0(n550), .D1(n494), .S(B[25]), .X(n682) );
  SEN_OAI21B_2 U780 ( .A1(net15865), .A2(n832), .B(n831), .X(n833) );
  SEN_ND2_T_4 U781 ( .A1(net15794), .A2(net15795), .X(net16215) );
  SEN_ND2_G_1 U782 ( .A1(net16223), .A2(net16222), .X(net15795) );
  SEN_NR3B_DG_8 U783 ( .A(n813), .B1(n644), .B2(n643), .X(n645) );
  SEN_ND2_S_1P5 U784 ( .A1(net16014), .A2(net17656), .X(n402) );
  SEN_EN2_8 U785 ( .A1(n358), .A2(n836), .X(n758) );
  SEN_MUXI2_S_1 U786 ( .D0(n550), .D1(n494), .S(B[15]), .X(n594) );
  SEN_ND4_S_3 U787 ( .A1(net16344), .A2(net16345), .A3(net16077), .A4(n364), 
        .X(net15798) );
  SEN_ND2_S_1 U788 ( .A1(net17656), .A2(net15897), .X(net16023) );
  SEN_OAI21_5 U789 ( .A1(n659), .A2(n658), .B(n657), .X(net15914) );
  SEN_INV_2 U790 ( .A(net16153), .X(n442) );
  SEN_EN2_8 U791 ( .A1(n806), .A2(n807), .X(n804) );
  SEN_ND2_S_6 U792 ( .A1(net16361), .A2(net16360), .X(net17414) );
  SEN_ND2_T_1P5 U793 ( .A1(n554), .A2(n608), .X(net16327) );
  SEN_MUXI2_S_2 U794 ( .D0(n551), .D1(n493), .S(B[8]), .X(n608) );
  SEN_OAI211_3 U795 ( .A1(net15963), .A2(net16412), .B1(net15964), .B2(
        net15965), .X(net3727) );
  SEN_ND2_T_2 U796 ( .A1(n518), .A2(B[16]), .X(n509) );
  SEN_ND2B_V1_4 U797 ( .A(net15915), .B(net15916), .X(net15912) );
  SEN_NR2B_V1_2 U798 ( .A(net17656), .B(n820), .X(n526) );
  SEN_ND2_T_2 U799 ( .A1(n544), .A2(n632), .X(n753) );
  SEN_ND2_T_4 U800 ( .A1(n630), .A2(n554), .X(n544) );
  SEN_ND2_2 U801 ( .A1(net16476), .A2(n595), .X(n638) );
  SEN_MUXI2_DG_2 U802 ( .D0(net16482), .D1(n683), .S(A[10]), .X(n642) );
  SEN_INV_2 U803 ( .A(net16407), .X(net16309) );
  SEN_ND2_T_1 U804 ( .A1(n651), .A2(n650), .X(n760) );
  SEN_NR2_T_4 U805 ( .A1(net16691), .A2(n451), .X(n490) );
  SEN_EN2_S_3 U806 ( .A1(n856), .A2(n851), .X(net15830) );
  SEN_INV_S_4 U807 ( .A(Z[20]), .X(n415) );
  SEN_OAI211_4 U808 ( .A1(net15817), .A2(net16410), .B1(net15818), .B2(
        net15819), .X(Z[20]) );
  SEN_ND2_T_1 U809 ( .A1(net17602), .A2(n642), .X(n646) );
  SEN_ND2_S_0P5 U810 ( .A1(n686), .A2(n685), .X(net16190) );
  SEN_INV_2 U811 ( .A(n685), .X(n713) );
  SEN_ND2_G_1 U812 ( .A1(net17602), .A2(n684), .X(n685) );
  SEN_OAI21_T_4 U813 ( .A1(net16410), .A2(net16155), .B(net16156), .X(net3724)
         );
  SEN_EN2_S_6 U814 ( .A1(n710), .A2(n706), .X(net16155) );
  SEN_OR3B_4 U815 ( .B1(Z[21]), .B2(Z[23]), .A(n381), .X(n388) );
  SEN_ND2_T_2 U816 ( .A1(n636), .A2(net17602), .X(n650) );
  SEN_INV_S_2 U817 ( .A(n484), .X(n636) );
  SEN_MUXI2_DG_0P75 U818 ( .D0(n550), .D1(n367), .S(B[27]), .X(n562) );
  SEN_EO2_3 U819 ( .A1(net15969), .A2(n531), .X(net15963) );
  SEN_AOI21B_4 U820 ( .A1(n654), .A2(n653), .B(n652), .X(n659) );
  SEN_EO2_1 U821 ( .A1(net15791), .A2(net15790), .X(net17005) );
  SEN_OAI21_2 U822 ( .A1(n734), .A2(n733), .B(n732), .X(n735) );
  SEN_INV_3 U823 ( .A(n733), .X(n737) );
  SEN_EO2_3 U824 ( .A1(n723), .A2(n725), .X(n733) );
  SEN_ND2_S_4 U825 ( .A1(n553), .A2(n602), .X(net16336) );
  SEN_EN2_5 U826 ( .A1(n789), .A2(n788), .X(n785) );
  SEN_INV_2 U827 ( .A(n748), .X(n465) );
  SEN_INV_6 U828 ( .A(Z[15]), .X(n426) );
  SEN_OAI211_8 U829 ( .A1(net15902), .A2(net16410), .B1(net15903), .B2(
        net15904), .X(Z[15]) );
  SEN_AOI21_6 U830 ( .A1(n672), .A2(n866), .B(n452), .X(n675) );
  SEN_INV_S_4 U831 ( .A(n660), .X(n810) );
  SEN_INV_0P65 U832 ( .A(net16127), .X(net16123) );
  SEN_INV_1 U833 ( .A(net15934), .X(net16013) );
  SEN_MUXI2_DG_3 U834 ( .D0(n551), .D1(n517), .S(B[17]), .X(n592) );
  SEN_ND2_T_2 U835 ( .A1(net16476), .A2(n603), .X(net16337) );
  SEN_OR4B_4 U836 ( .B1(n694), .B2(n693), .B3(n692), .A(n691), .X(n706) );
  SEN_ND2_8 U837 ( .A1(net15916), .A2(net17750), .X(net18157) );
  SEN_NR2_8 U838 ( .A1(n513), .A2(n491), .X(n512) );
  SEN_EN2_S_2 U839 ( .A1(n527), .A2(n827), .X(net15869) );
  SEN_OAI211_3 U840 ( .A1(net15869), .A2(net16410), .B1(net15870), .B2(
        net15871), .X(Z[10]) );
  SEN_NR2_T_2 U841 ( .A1(net3721), .A2(Z[10]), .X(n425) );
  SEN_INV_S_6 U842 ( .A(n658), .X(n814) );
  SEN_EN2_5 U843 ( .A1(n762), .A2(n763), .X(n658) );
  SEN_INV_1 U844 ( .A(n770), .X(n821) );
  SEN_BUF_8 U845 ( .A(INST[0]), .X(net16501) );
  SEN_EN2_3 U846 ( .A1(net16999), .A2(n711), .X(net16144) );
  SEN_OA21_2 U847 ( .A1(n442), .A2(net16084), .B(net16999), .X(net17035) );
  SEN_EO2_G_2 U848 ( .A1(n712), .A2(n713), .X(net16999) );
  SEN_ND2_T_4 U849 ( .A1(n627), .A2(n554), .X(net16288) );
  SEN_OR3B_4 U850 ( .B1(n721), .B2(n731), .A(n720), .X(n722) );
  SEN_ND2_6 U851 ( .A1(net15916), .A2(net17750), .X(n398) );
  SEN_EN2_S_1 U852 ( .A1(n702), .A2(FLAGS[1]), .X(FLAGS[0]) );
  SEN_AO2BB2_2 U853 ( .A1(n702), .A2(n705), .B1(n701), .B2(n709), .X(FLAGS[1])
         );
  SEN_EO2_2 U854 ( .A1(n821), .A2(n773), .X(n776) );
  SEN_ND2_S_4 U855 ( .A1(n459), .A2(n460), .X(net15902) );
  SEN_ND3_T_4 U856 ( .A1(n400), .A2(net16215), .A3(net17005), .X(net16127) );
  SEN_ND4B_4 U857 ( .A(net15798), .B1(n398), .B2(net15795), .B3(net15796), .X(
        n400) );
  SEN_OAOI211_2 U858 ( .A1(net16023), .A2(n820), .B(n521), .C(net15882), .X(
        n773) );
  SEN_ND2_4 U859 ( .A1(n765), .A2(n492), .X(n813) );
  SEN_ND2_4 U860 ( .A1(n450), .A2(net17829), .X(n457) );
  SEN_INV_1 U861 ( .A(net15883), .X(net17829) );
  SEN_INV_S_1 U862 ( .A(n576), .X(n723) );
  SEN_INV_S_1 U863 ( .A(n715), .X(n470) );
  SEN_EO2_2 U864 ( .A1(net15889), .A2(net15888), .X(n523) );
  SEN_INV_S_1 U865 ( .A(net16165), .X(net16410) );
  SEN_ND2_2 U866 ( .A1(n683), .A2(A[13]), .X(n483) );
  SEN_INV_2 U867 ( .A(n559), .X(n698) );
  SEN_ND2_S_3 U868 ( .A1(n785), .A2(n791), .X(n797) );
  SEN_INV_3 U869 ( .A(net17600), .X(net17602) );
  SEN_BUF_6 U870 ( .A(INST[3]), .X(net16495) );
  SEN_INV_S_4 U871 ( .A(net16301), .X(net15967) );
  SEN_INV_2 U872 ( .A(n488), .X(n489) );
  SEN_INV_1 U873 ( .A(net16326), .X(net15889) );
  SEN_EN2_0P5 U874 ( .A1(n810), .A2(n811), .X(n378) );
  SEN_INV_S_2 U875 ( .A(n879), .X(n462) );
  SEN_INV_S_1 U876 ( .A(net16193), .X(n439) );
  SEN_EO2_S_0P5 U877 ( .A1(n739), .A2(n741), .X(n579) );
  SEN_INV_S_1 U878 ( .A(net16424), .X(net16772) );
  SEN_ND2_G_1 U879 ( .A1(net18219), .A2(n821), .X(n775) );
  SEN_EO2_G_2 U880 ( .A1(net16070), .A2(net16069), .X(net17000) );
  SEN_ND2_G_1 U881 ( .A1(net16196), .A2(net16197), .X(net16134) );
  SEN_EN2_1 U882 ( .A1(n439), .A2(net16134), .X(net16938) );
  SEN_INV_2 U883 ( .A(net16165), .X(net16412) );
  SEN_EN2_1 U884 ( .A1(n730), .A2(n728), .X(n535) );
  SEN_ND2_S_3 U885 ( .A1(n407), .A2(n408), .X(n406) );
  SEN_ND2_G_1 U886 ( .A1(net16669), .A2(A[12]), .X(n473) );
  SEN_INV_S_1 U887 ( .A(B[13]), .X(n541) );
  SEN_ND2_G_1 U888 ( .A1(n482), .A2(n483), .X(n484) );
  SEN_MUXI2_S_1 U889 ( .D0(net16480), .D1(n683), .S(A[15]), .X(n595) );
  SEN_INV_6 U890 ( .A(net16478), .X(net16476) );
  SEN_ND2_G_1 U891 ( .A1(n553), .A2(n582), .X(n670) );
  SEN_ND2_G_1 U892 ( .A1(net17602), .A2(n586), .X(n674) );
  SEN_INV_1 U893 ( .A(net16074), .X(net16220) );
  SEN_ND2_G_1 U894 ( .A1(net17602), .A2(n679), .X(n681) );
  SEN_ND2_G_1 U895 ( .A1(n555), .A2(n678), .X(n680) );
  SEN_MUXI2_S_0P5 U896 ( .D0(net16482), .D1(n549), .S(A[25]), .X(n684) );
  SEN_OAI21_S_2 U897 ( .A1(net17035), .A2(net16143), .B(net16938), .X(net16188) );
  SEN_INV_S_3 U898 ( .A(net16289), .X(net15979) );
  SEN_INV_S_1 U899 ( .A(B[3]), .X(n546) );
  SEN_INV_3 U900 ( .A(net15769), .X(net16691) );
  SEN_INV_1 U901 ( .A(n671), .X(n861) );
  SEN_ND2_2 U902 ( .A1(n668), .A2(n669), .X(n866) );
  SEN_INV_S_1 U903 ( .A(n686), .X(n712) );
  SEN_INV_S_1 U904 ( .A(n575), .X(n728) );
  SEN_ND2_S_1 U905 ( .A1(n535), .A2(n537), .X(n718) );
  SEN_INV_3 U906 ( .A(net16501), .X(net16182) );
  SEN_INV_3 U907 ( .A(net17601), .X(net16478) );
  SEN_INV_2 U908 ( .A(net17600), .X(net17601) );
  SEN_AOI21B_1 U909 ( .A1(n793), .A2(n792), .B(n791), .X(n794) );
  SEN_ND2_T_1 U910 ( .A1(n771), .A2(n467), .X(n469) );
  SEN_INV_S_1 U911 ( .A(n662), .X(n880) );
  SEN_ND2_G_1 U912 ( .A1(n539), .A2(n879), .X(n463) );
  SEN_ND2_G_1 U913 ( .A1(n461), .A2(n462), .X(n464) );
  SEN_ND2_T_1 U914 ( .A1(n364), .A2(net18157), .X(n840) );
  SEN_EN2_DG_1 U915 ( .A1(n886), .A2(n889), .X(n537) );
  SEN_OAI211_1 U916 ( .A1(net15986), .A2(net16412), .B1(net15987), .B2(
        net15988), .X(Z[1]) );
  SEN_EN2_1 U917 ( .A1(n793), .A2(n792), .X(net15986) );
  SEN_OAOI211_G_1 U918 ( .A1(B[8]), .A2(A[8]), .B(net16444), .C(n774), .X(
        net16018) );
  SEN_OA21_2 U919 ( .A1(n776), .A2(net16412), .B(n775), .X(net17804) );
  SEN_OAI211_3 U920 ( .A1(net16078), .A2(net16412), .B1(net16079), .B2(
        net16080), .X(net3748) );
  SEN_ND2_2 U921 ( .A1(n453), .A2(n454), .X(net16078) );
  SEN_OAI211_3 U922 ( .A1(n434), .A2(n443), .B1(n435), .B2(n436), .X(net3754)
         );
  SEN_ND2B_6 U923 ( .A(net16495), .B(n393), .X(n395) );
  SEN_INV_S_2 U924 ( .A(Z[13]), .X(n424) );
  SEN_ND3_S_0P5 U925 ( .A1(n814), .A2(n813), .A3(n834), .X(n815) );
  SEN_AOAI211_8 U926 ( .A1(n389), .A2(net16497), .B(net16501), .C(n390), .X(
        net16177) );
  SEN_ND2_12 U927 ( .A1(net17349), .A2(net17579), .X(net16669) );
  SEN_OAOI211_G_1 U928 ( .A1(B[2]), .A2(A[2]), .B(net16444), .C(n795), .X(
        net15977) );
  SEN_INV_S_1 U929 ( .A(n704), .X(n558) );
  SEN_ND2_G_4 U930 ( .A1(n486), .A2(n487), .X(net16985) );
  SEN_INV_S_3 U931 ( .A(net3748), .X(n418) );
  SEN_ND2_S_2 U932 ( .A1(n440), .A2(n446), .X(n449) );
  SEN_ND2_2 U933 ( .A1(n448), .A2(n449), .X(n434) );
  SEN_ND2_S_0P5 U934 ( .A1(n704), .A2(n542), .X(net16165) );
  SEN_ND2_S_3 U935 ( .A1(n767), .A2(n768), .X(n515) );
  SEN_EO2_G_4 U936 ( .A1(n766), .A2(n530), .X(net16028) );
  SEN_INV_S_1 U937 ( .A(net16691), .X(net16774) );
  SEN_ND2B_V1_3 U938 ( .A(net16478), .B(n631), .X(n632) );
  SEN_INV_S_3 U939 ( .A(n552), .X(n550) );
  SEN_INV_S_8 U940 ( .A(n552), .X(n551) );
  SEN_AN2_S_1 U941 ( .A1(n543), .A2(n365), .X(n371) );
  SEN_INV_S_1 U942 ( .A(n556), .X(n555) );
  SEN_OR2_1 U943 ( .A1(A[31]), .A2(B[31]), .X(n372) );
  SEN_OR2_1 U944 ( .A1(A[29]), .A2(B[29]), .X(n373) );
  SEN_OR2_1 U945 ( .A1(A[30]), .A2(B[30]), .X(n374) );
  SEN_INV_S_1 U946 ( .A(n359), .X(net16448) );
  SEN_NR2_0P8 U947 ( .A1(n399), .A2(net15960), .X(net15958) );
  SEN_MUXI2_S_1 U948 ( .D0(net16480), .D1(n549), .S(A[20]), .X(n584) );
  SEN_NR3_T_0P5 U949 ( .A1(n861), .A2(n860), .A3(net16774), .X(n862) );
  SEN_ND2B_S_4 U950 ( .A(net16179), .B(net16400), .X(n700) );
  SEN_MUXI2_DG_1 U951 ( .D0(n551), .D1(n494), .S(B[10]), .X(n641) );
  SEN_ND2_T_6 U952 ( .A1(net16361), .A2(net16179), .X(n392) );
  SEN_ND2B_V1_1 U953 ( .A(A[31]), .B(net16497), .X(n695) );
  SEN_INV_0P65 U954 ( .A(net15894), .X(net15883) );
  SEN_MUXI2_DG_1 U955 ( .D0(net16482), .D1(net16669), .S(A[5]), .X(n613) );
  SEN_INV_4 U956 ( .A(net16499), .X(n393) );
  SEN_INV_8 U957 ( .A(net17655), .X(net17656) );
  SEN_INV_0P8 U958 ( .A(n440), .X(n447) );
  SEN_EN2_S_3 U959 ( .A1(n859), .A2(n858), .X(net15817) );
  SEN_INV_1 U960 ( .A(n669), .X(n853) );
  SEN_INV_S_8 U961 ( .A(net17749), .X(net17750) );
  SEN_INV_S_3 U962 ( .A(n503), .X(n627) );
  SEN_INV_4 U963 ( .A(net16495), .X(net16400) );
  SEN_ND2_T_1P5 U964 ( .A1(n478), .A2(n479), .X(n480) );
  SEN_ND2_G_1 U965 ( .A1(n550), .A2(n540), .X(n479) );
  SEN_NR3_0P8 U966 ( .A1(net15940), .A2(net16723), .A3(net16422), .X(net15939)
         );
  SEN_ND2_2 U967 ( .A1(n796), .A2(net15961), .X(net17427) );
  SEN_INV_4 U968 ( .A(net17427), .X(net17428) );
  SEN_ND3_S_8 U969 ( .A1(n814), .A2(n834), .A3(net16985), .X(n644) );
  SEN_INV_2 U970 ( .A(n656), .X(n762) );
  SEN_NR3B_3 U971 ( .A(net15796), .B1(net15797), .B2(net15798), .X(n875) );
  SEN_MUXI2_S_3 U972 ( .D0(n683), .D1(net16482), .S(n545), .X(n626) );
  SEN_ND2_0P5 U973 ( .A1(net18219), .A2(n524), .X(net15996) );
  SEN_INV_S_1 U974 ( .A(n865), .X(n859) );
  SEN_AO21_4 U975 ( .A1(n845), .A2(n866), .B(n865), .X(n452) );
  SEN_ND2_S_0P5 U976 ( .A1(n866), .A2(n848), .X(n863) );
  SEN_ND2_1P5 U977 ( .A1(n664), .A2(n665), .X(n848) );
  SEN_INV_0P5 U978 ( .A(n780), .X(n783) );
  SEN_INV_S_4 U979 ( .A(n749), .X(n475) );
  SEN_INV_4 U980 ( .A(net17189), .X(net17190) );
  SEN_ND2_T_2 U981 ( .A1(n607), .A2(n606), .X(net15899) );
  SEN_AN2_6 U982 ( .A1(net16400), .A2(net16182), .X(net16968) );
  SEN_NR2B_2 U983 ( .A(net18157), .B(net15829), .X(n857) );
  SEN_INV_S_0P5 U984 ( .A(net16300), .X(net15968) );
  SEN_ND2_6 U985 ( .A1(n394), .A2(n395), .X(n389) );
  SEN_INV_2 U986 ( .A(n655), .X(n763) );
  SEN_ND2_2 U987 ( .A1(net16400), .A2(net16182), .X(n379) );
  SEN_BUF_1 U988 ( .A(net16361), .X(n382) );
  SEN_MUXI2_S_1 U989 ( .D0(net16480), .D1(n549), .S(A[24]), .X(n679) );
  SEN_ND2_T_2 U990 ( .A1(n842), .A2(n665), .X(n384) );
  SEN_INV_S_3 U991 ( .A(n842), .X(n383) );
  SEN_NR3B_3 U992 ( .A(net18157), .B1(n864), .B2(n863), .X(n870) );
  SEN_OAI31_1 U993 ( .A1(net16495), .A2(net16309), .A3(net16182), .B(n621), 
        .X(n622) );
  SEN_ND2_6 U994 ( .A1(n645), .A2(n751), .X(net17749) );
  SEN_MUXI2_DG_1 U995 ( .D0(n550), .D1(n368), .S(B[19]), .X(n587) );
  SEN_INV_1 U996 ( .A(n866), .X(n589) );
  SEN_INV_0P8 U997 ( .A(net16499), .X(net17564) );
  SEN_ND2_4 U998 ( .A1(n515), .A2(n516), .X(n765) );
  SEN_ND2_G_1 U999 ( .A1(n848), .A2(n543), .X(net15829) );
  SEN_AO222_1 U1000 ( .A1(net18219), .A2(n737), .B1(n359), .B2(n373), .C1(n725), .C2(n724), .X(n386) );
  SEN_BUF_1 U1001 ( .A(n532), .X(n387) );
  SEN_ND2_S_0P5 U1002 ( .A1(net16434), .A2(n387), .X(net15847) );
  SEN_OAI21_S_0P5 U1003 ( .A1(n520), .A2(n362), .B(n387), .X(n849) );
  SEN_INV_S_3 U1004 ( .A(net3751), .X(n408) );
  SEN_NR3_0P5 U1005 ( .A1(n807), .A2(n806), .A3(net16772), .X(n808) );
  SEN_INV_8 U1006 ( .A(n392), .X(net17349) );
  SEN_OR2_2 U1007 ( .A1(n885), .A2(n537), .X(n548) );
  SEN_INV_1 U1008 ( .A(n816), .X(n458) );
  SEN_ND2_S_4 U1009 ( .A1(n466), .A2(net16074), .X(n749) );
  SEN_INV_1P5 U1010 ( .A(n391), .X(n390) );
  SEN_INV_S_0P5 U1011 ( .A(n382), .X(net18246) );
  SEN_ND2_S_0P5 U1012 ( .A1(net16361), .A2(net17579), .X(net16201) );
  SEN_ND2B_V1DG_2 U1013 ( .A(A[31]), .B(net16968), .X(net17579) );
  SEN_ND2_6 U1014 ( .A1(net17190), .A2(net17428), .X(net16015) );
  SEN_OAI221_4 U1015 ( .A1(net16949), .A2(net15961), .B1(n403), .B2(net16949), 
        .C(net15953), .X(net15897) );
  SEN_OR2_2 U1016 ( .A1(n401), .A2(n402), .X(net17773) );
  SEN_ND2_2 U1017 ( .A1(net16326), .A2(net16325), .X(net15880) );
  SEN_ND2_G_1 U1018 ( .A1(net16328), .A2(net16327), .X(net15894) );
  SEN_INV_4 U1019 ( .A(n399), .X(n403) );
  SEN_ND2_3 U1020 ( .A1(net16300), .A2(net16301), .X(net15946) );
  SEN_NR2B_V1DG_1 U1021 ( .A(net15942), .B(net15960), .X(net15956) );
  SEN_BUF_1 U1022 ( .A(net15942), .X(net16701) );
  SEN_NR4_3 U1023 ( .A1(n404), .A2(n405), .A3(n406), .A4(net3724), .X(FLAGS[2]) );
  SEN_ND3_S_4 U1024 ( .A1(n411), .A2(n412), .A3(n413), .X(n404) );
  SEN_AN3B_4 U1025 ( .B1(n417), .B2(n418), .A(n419), .X(n411) );
  SEN_NR2_S_4 U1026 ( .A1(n427), .A2(Z[11]), .X(n444) );
  SEN_ND3_S_4 U1027 ( .A1(n428), .A2(n429), .A3(n430), .X(n427) );
  SEN_OAI211_3 U1028 ( .A1(net16005), .A2(net16412), .B1(net16006), .B2(
        net16007), .X(net3715) );
  SEN_NR4_6 U1029 ( .A1(net3730), .A2(net3712), .A3(n431), .A4(net3733), .X(
        n429) );
  SEN_OAI211_3 U1030 ( .A1(net15936), .A2(net16412), .B1(net15937), .B2(
        net15938), .X(net3730) );
  SEN_ND2_S_3 U1031 ( .A1(n432), .A2(n433), .X(n431) );
  SEN_INV_2 U1032 ( .A(net3727), .X(n432) );
  SEN_OAI211_8 U1033 ( .A1(net15947), .A2(net16412), .B1(net15948), .B2(
        net15949), .X(net3733) );
  SEN_OAI211_4 U1034 ( .A1(net16037), .A2(net16412), .B1(net16038), .B2(
        net16039), .X(Z[14]) );
  SEN_NR2_S_4 U1035 ( .A1(n423), .A2(Z[16]), .X(n421) );
  SEN_ND3_S_4 U1036 ( .A1(n424), .A2(n426), .A3(n425), .X(n423) );
  SEN_OAI211_2 U1037 ( .A1(net15857), .A2(net16410), .B1(net15858), .B2(
        net15859), .X(Z[13]) );
  SEN_OAI211_1 U1038 ( .A1(net15919), .A2(net16410), .B1(net15920), .B2(
        net15921), .X(Z[16]) );
  SEN_OAI211_3 U1039 ( .A1(net15846), .A2(net16410), .B1(net15847), .B2(
        net15848), .X(Z[18]) );
  SEN_ND2_T_6 U1040 ( .A1(net17713), .A2(net15775), .X(Z[17]) );
  SEN_ND2_2 U1041 ( .A1(n447), .A2(net16938), .X(n448) );
  SEN_INV_S_0P5 U1042 ( .A(net16938), .X(n446) );
  SEN_INV_S_0P5 U1043 ( .A(net16165), .X(n443) );
  SEN_ND2_S_0P5 U1044 ( .A1(net18219), .A2(net16938), .X(n435) );
  SEN_OA2BB2_0P5 U1045 ( .A1(net16134), .A2(n437), .B1(n438), .B2(net16448), 
        .X(n436) );
  SEN_NR2_S_0P5 U1046 ( .A1(n439), .A2(net16774), .X(n437) );
  SEN_NR2_1 U1047 ( .A1(A[26]), .A2(B[26]), .X(n438) );
  SEN_INV_S_0P5 U1048 ( .A(net16190), .X(net16143) );
  SEN_AO21B_6 U1049 ( .A1(net16073), .A2(net16074), .B(net17000), .X(net15794)
         );
  SEN_NR2_T_2 U1050 ( .A1(net16127), .A2(net16188), .X(net17788) );
  SEN_ND2_6 U1051 ( .A1(net16057), .A2(n813), .X(n832) );
  SEN_AN2_3 U1052 ( .A1(net18157), .A2(n846), .X(n519) );
  SEN_INV_S_2 U1053 ( .A(n777), .X(n467) );
  SEN_NR3_T_3 U1054 ( .A1(n747), .A2(net16220), .A3(n589), .X(net16344) );
  SEN_INV_2 U1055 ( .A(n868), .X(n747) );
  SEN_ND2_0P8 U1056 ( .A1(n551), .A2(n507), .X(n508) );
  SEN_INV_S_4 U1057 ( .A(net15899), .X(net17655) );
  SEN_ND2B_4 U1058 ( .A(net16497), .B(net16495), .X(n557) );
  SEN_INV_S_6 U1059 ( .A(net18157), .X(net15797) );
  SEN_ND2_2 U1060 ( .A1(n465), .A2(net17799), .X(n466) );
  SEN_INV_S_2 U1061 ( .A(n646), .X(n829) );
  SEN_EO2_2 U1062 ( .A1(n387), .A2(n841), .X(net15846) );
  SEN_OAOI211_3 U1063 ( .A1(n840), .A2(n839), .B(n520), .C(n362), .X(n841) );
  SEN_ND2_2 U1064 ( .A1(n544), .A2(n632), .X(n516) );
  SEN_INV_2 U1065 ( .A(n818), .X(n485) );
  SEN_ND2_S_2 U1066 ( .A1(n637), .A2(n818), .X(n487) );
  SEN_NR3_0P5 U1067 ( .A1(net16774), .A2(n818), .A3(n817), .X(n819) );
  SEN_ND3_T_0P8 U1068 ( .A1(net16495), .A2(net16497), .A3(net16501), .X(n583)
         );
  SEN_ND2_S_1P5 U1069 ( .A1(net17602), .A2(n634), .X(n655) );
  SEN_NR2_T_3 U1070 ( .A1(net17564), .A2(n379), .X(n497) );
  SEN_AN2_3 U1071 ( .A1(n365), .A2(n846), .X(n525) );
  SEN_INV_1 U1072 ( .A(n845), .X(n856) );
  SEN_MUXI2_S_1 U1073 ( .D0(n550), .D1(n517), .S(B[20]), .X(n582) );
  SEN_ND2B_V1_1 U1074 ( .A(n583), .B(net16499), .X(net16180) );
  SEN_MUXI2_S_2 U1075 ( .D0(net16480), .D1(n683), .S(A[18]), .X(n591) );
  SEN_EN2_DG_4 U1076 ( .A1(n805), .A2(net15934), .X(net15927) );
  SEN_AOI21B_4 U1077 ( .A1(n885), .A2(n537), .B(n726), .X(n727) );
  SEN_ND2_1P5 U1078 ( .A1(net16476), .A2(n588), .X(n669) );
  SEN_NR3_T_0P5 U1079 ( .A1(net15967), .A2(net15968), .A3(net15769), .X(n798)
         );
  SEN_ND2_T_1P5 U1080 ( .A1(net16476), .A2(n601), .X(net16325) );
  SEN_INV_2 U1081 ( .A(net16325), .X(net15888) );
  SEN_MUXI2_S_2 U1082 ( .D0(net16480), .D1(n683), .S(A[9]), .X(n601) );
  SEN_MUX2_1 U1083 ( .D0(n512), .D1(n552), .S(n546), .X(n625) );
  SEN_INV_S_1 U1084 ( .A(net16440), .X(net18219) );
  SEN_OR2_DG_1 U1085 ( .A1(n560), .A2(n363), .X(net16440) );
  SEN_MUXI2_S_3 U1086 ( .D0(n551), .D1(n494), .S(B[1]), .X(n614) );
  SEN_MUXI2_S_1 U1087 ( .D0(n550), .D1(n494), .S(B[9]), .X(n600) );
  SEN_OAI21_S_0P5 U1088 ( .A1(n534), .A2(n832), .B(n759), .X(n831) );
  SEN_MUXI2_DG_3 U1089 ( .D0(n551), .D1(n517), .S(B[11]), .X(n630) );
  SEN_INV_1 U1090 ( .A(net15969), .X(net18184) );
  SEN_INV_S_0P5 U1091 ( .A(n804), .X(n805) );
  SEN_EO2_G_4 U1092 ( .A1(net15953), .A2(n801), .X(net15947) );
  SEN_INV_S_0P5 U1093 ( .A(net15945), .X(net15969) );
  SEN_OAOI211_G_1 U1094 ( .A1(B[3]), .A2(A[3]), .B(net16444), .C(n798), .X(
        net15965) );
  SEN_EN2_S_2 U1095 ( .A1(net16701), .A2(n803), .X(net15936) );
  SEN_INV_S_0P5 U1096 ( .A(net16073), .X(net17799) );
  SEN_MUXI2_S_1 U1097 ( .D0(n551), .D1(n518), .S(B[14]), .X(n633) );
  SEN_ND2_T_1 U1098 ( .A1(n553), .A2(n600), .X(net16326) );
  SEN_EO2_S_3 U1099 ( .A1(n872), .A2(n873), .X(n522) );
  SEN_MUXI2_S_2 U1100 ( .D0(net16480), .D1(n549), .S(A[19]), .X(n588) );
  SEN_ND2_3 U1101 ( .A1(net16476), .A2(n640), .X(n648) );
  SEN_ND3B_V1DG_1 U1102 ( .A(net16499), .B1(net16501), .B2(net16497), .X(n563)
         );
  SEN_INV_1 U1103 ( .A(net17572), .X(net17573) );
  SEN_NR3_T_0P5 U1104 ( .A1(net16009), .A2(net16010), .A3(net16772), .X(n779)
         );
  SEN_ND2B_V1DG_2 U1105 ( .A(A[31]), .B(net16968), .X(net16360) );
  SEN_INV_2 U1106 ( .A(n648), .X(n756) );
  SEN_ND2_S_3 U1107 ( .A1(net16476), .A2(n613), .X(net16298) );
  SEN_MUXI2_S_4 U1108 ( .D0(net16482), .D1(n683), .S(A[0]), .X(n619) );
  SEN_INV_S_0P5 U1109 ( .A(n765), .X(n766) );
  SEN_BUF_S_4 U1110 ( .A(n753), .X(n492) );
  SEN_ND2_2 U1111 ( .A1(net16476), .A2(n591), .X(n665) );
  SEN_EO2_G_4 U1112 ( .A1(n828), .A2(n829), .X(n527) );
  SEN_EO2_G_2 U1113 ( .A1(n814), .A2(n761), .X(net16037) );
  SEN_INV_S_2 U1114 ( .A(n616), .X(n789) );
  SEN_AN2_2 U1115 ( .A1(n752), .A2(net15865), .X(n530) );
  SEN_INV_0P65 U1116 ( .A(n706), .X(n702) );
  SEN_MUXI2_S_3 U1117 ( .D0(net16482), .D1(net16669), .S(A[6]), .X(n605) );
  SEN_ND2_2 U1118 ( .A1(n637), .A2(n638), .X(net16077) );
  SEN_ND2_T_3 U1119 ( .A1(n817), .A2(n485), .X(n486) );
  SEN_NR3_0P5 U1120 ( .A1(net16499), .A2(n695), .A3(net16182), .X(n697) );
  SEN_INV_2 U1121 ( .A(net16327), .X(net16021) );
  SEN_NR4B_4 U1122 ( .A(net18157), .B1(n864), .B2(n747), .B3(n863), .X(n748)
         );
  SEN_BUF_3 U1123 ( .A(n746), .X(n543) );
  SEN_ND2_2 U1124 ( .A1(n880), .A2(n663), .X(n455) );
  SEN_ND2_2 U1125 ( .A1(n458), .A2(net17816), .X(n460) );
  SEN_INV_S_0P5 U1126 ( .A(net16985), .X(net17816) );
  SEN_OAI31_3 U1127 ( .A1(net15910), .A2(n815), .A3(net15912), .B(net15913), 
        .X(n816) );
  SEN_INV_S_1 U1128 ( .A(n539), .X(n461) );
  SEN_ND2_2 U1129 ( .A1(n468), .A2(n469), .X(net16005) );
  SEN_INV_S_1 U1130 ( .A(A[12]), .X(n471) );
  SEN_INV_S_3 U1131 ( .A(n474), .X(n640) );
  SEN_ND2_S_4 U1132 ( .A1(net17760), .A2(n475), .X(n477) );
  SEN_INV_S_1 U1133 ( .A(net17000), .X(net17760) );
  SEN_INV_2 U1134 ( .A(n480), .X(n590) );
  SEN_ND2_G_1 U1135 ( .A1(net16482), .A2(n481), .X(n482) );
  SEN_INV_1 U1136 ( .A(A[13]), .X(n481) );
  SEN_ND2_S_0P5 U1137 ( .A1(net16434), .A2(net16985), .X(net15904) );
  SEN_OAOI211_8 U1138 ( .A1(B[17]), .A2(A[17]), .B(net16444), .C(n882), .X(
        net15775) );
  SEN_AOAI211_3 U1139 ( .A1(n525), .A2(n857), .B(n867), .C(n866), .X(n858) );
  SEN_ND2_G_1 U1140 ( .A1(net16434), .A2(n834), .X(net15858) );
  SEN_INV_S_0P5 U1141 ( .A(n378), .X(n809) );
  SEN_INV_0P8 U1142 ( .A(net16478), .X(net16474) );
  SEN_INV_S_0P5 U1143 ( .A(net16448), .X(net17584) );
  SEN_OAOI211_2 U1144 ( .A1(B[5]), .A2(A[5]), .B(net16444), .C(n802), .X(
        net15949) );
  SEN_OAOI211_2 U1145 ( .A1(B[6]), .A2(A[6]), .B(net16444), .C(n808), .X(
        net15929) );
  SEN_OAOI211_1 U1146 ( .A1(B[4]), .A2(A[4]), .B(net16444), .C(net15939), .X(
        net15938) );
  SEN_INV_S_0P5 U1147 ( .A(n492), .X(n496) );
  SEN_ND2_G_1 U1148 ( .A1(n551), .A2(n500), .X(n501) );
  SEN_INV_1 U1149 ( .A(B[2]), .X(n500) );
  SEN_INV_1 U1150 ( .A(net16188), .X(net16125) );
  SEN_INV_1 U1151 ( .A(n674), .X(n873) );
  SEN_INV_0P8 U1152 ( .A(n681), .X(n744) );
  SEN_INV_S_1 U1153 ( .A(B[16]), .X(n507) );
  SEN_OAOI211_1 U1154 ( .A1(B[25]), .A2(A[25]), .B(n359), .C(n714), .X(
        net16146) );
  SEN_NR2_S_0P5 U1155 ( .A1(n718), .A2(n581), .X(n690) );
  SEN_ND2B_1 U1156 ( .A(n726), .B(n535), .X(n716) );
  SEN_OAOI211_1 U1157 ( .A1(B[22]), .A2(A[22]), .B(net17584), .C(n750), .X(
        net16065) );
  SEN_NR3_0P5 U1158 ( .A1(n843), .A2(n842), .A3(net16774), .X(n844) );
  SEN_NR3_0P5 U1159 ( .A1(n829), .A2(n828), .A3(net16772), .X(n830) );
  SEN_MUXI2_S_0P5 U1160 ( .D0(net16482), .D1(net16669), .S(A[14]), .X(n634) );
  SEN_NR3_T_0P5 U1161 ( .A1(net15888), .A2(net15889), .A3(net16772), .X(n825)
         );
  SEN_INV_1 U1162 ( .A(n705), .X(n710) );
  SEN_ND2_S_0P5 U1163 ( .A1(n656), .A2(n655), .X(n657) );
  SEN_ND2_S_0P5 U1164 ( .A1(n580), .A2(n889), .X(n726) );
  SEN_ND2_S_0P5 U1165 ( .A1(n555), .A2(n699), .X(n701) );
  SEN_OAOI211_0P5 U1166 ( .A1(B[13]), .A2(A[13]), .B(net16444), .C(n837), .X(
        net15859) );
  SEN_OAOI211_1 U1167 ( .A1(B[14]), .A2(A[14]), .B(net16444), .C(n764), .X(
        net16039) );
  SEN_INV_1 U1168 ( .A(net16448), .X(net16444) );
  SEN_ND2_G_1 U1169 ( .A1(n737), .A2(n742), .X(n581) );
  SEN_NR3_0P5 U1170 ( .A1(n881), .A2(n880), .A3(net16774), .X(n882) );
  SEN_NR3_0P5 U1171 ( .A1(n744), .A2(n743), .A3(net16772), .X(n745) );
  SEN_ND3_S_0P5 U1172 ( .A1(net16153), .A2(net16154), .A3(net16190), .X(n719)
         );
  SEN_AOI222_1 U1173 ( .A1(net16434), .A2(n710), .B1(net17584), .B2(n372), 
        .C1(n709), .C2(n708), .X(net16156) );
  SEN_INV_S_1 U1174 ( .A(net16191), .X(net15791) );
  SEN_OAOI211_1 U1175 ( .A1(B[21]), .A2(A[21]), .B(net17584), .C(n874), .X(
        net15800) );
  SEN_ND2_S_0P5 U1176 ( .A1(net16434), .A2(n522), .X(net15801) );
  SEN_OAOI211_1 U1177 ( .A1(B[19]), .A2(A[19]), .B(net17584), .C(n854), .X(
        net15832) );
  SEN_ND2_G_1 U1178 ( .A1(n574), .A2(n573), .X(n741) );
  SEN_OAOI211_1 U1179 ( .A1(B[20]), .A2(A[20]), .B(net17584), .C(n862), .X(
        net15819) );
  SEN_OAOI211_1 U1180 ( .A1(B[24]), .A2(A[24]), .B(n359), .C(n745), .X(
        net16080) );
  SEN_MUXI2_S_0P5 U1181 ( .D0(n551), .D1(n368), .S(B[23]), .X(n676) );
  SEN_AN2_S_0P5 U1182 ( .A1(n533), .A2(n838), .X(n520) );
  SEN_INV_S_0P5 U1183 ( .A(net16440), .X(net16434) );
  SEN_NR3_0P5 U1184 ( .A1(net16774), .A2(net15790), .A3(net15791), .X(n877) );
  SEN_NR3_0P5 U1185 ( .A1(net16774), .A2(n873), .A3(n872), .X(n874) );
  SEN_NR3_0P5 U1186 ( .A1(net16774), .A2(net16069), .A3(net16070), .X(n750) );
  SEN_OA21B_1 U1187 ( .A1(net15865), .A2(n528), .B(n529), .X(n761) );
  SEN_NR3_T_0P5 U1188 ( .A1(n713), .A2(n712), .A3(net16772), .X(n714) );
  SEN_INV_1 U1189 ( .A(n579), .X(n742) );
  SEN_INV_1 U1190 ( .A(n731), .X(n734) );
  SEN_NR2_S_0P5 U1191 ( .A1(n723), .A2(net16774), .X(n724) );
  SEN_NR2_S_0P5 U1192 ( .A1(n739), .A2(net16774), .X(n740) );
  SEN_NR2_S_0P5 U1193 ( .A1(n707), .A2(net16774), .X(n708) );
  SEN_NR2_S_0P5 U1194 ( .A1(n886), .A2(net16774), .X(n888) );
  SEN_OAI21_S_0P5 U1195 ( .A1(n732), .A2(n579), .B(n578), .X(n692) );
  SEN_NR2_S_0P5 U1196 ( .A1(n716), .A2(n581), .X(n694) );
  SEN_NR2_G_0P5 U1197 ( .A1(n717), .A2(n581), .X(n693) );
  SEN_NR2_S_0P5 U1198 ( .A1(n715), .A2(n718), .X(n721) );
  SEN_NR2_S_0P5 U1199 ( .A1(n728), .A2(net16422), .X(n729) );
  SEN_ND2_S_0P5 U1200 ( .A1(n730), .A2(n729), .X(net16103) );
  SEN_AOI22_0P5 U1201 ( .A1(net18219), .A2(n535), .B1(n359), .B2(n538), .X(
        net16104) );
  SEN_ND2_G_1 U1202 ( .A1(n670), .A2(n671), .X(n868) );
  SEN_ND2_S_0P5 U1203 ( .A1(net18219), .A2(n537), .X(net15762) );
  SEN_AN2_S_0P5 U1204 ( .A1(net16501), .A2(n542), .X(n536) );
  SEN_AN3B_0P5 U1205 ( .B1(net16298), .B2(net17648), .A(net16772), .X(n802) );
  SEN_ND2_S_0P5 U1206 ( .A1(n576), .A2(n725), .X(n732) );
  SEN_ND2_S_0P5 U1207 ( .A1(n575), .A2(n730), .X(n717) );
  SEN_ND2_S_0P5 U1208 ( .A1(n577), .A2(n741), .X(n578) );
  SEN_INV_S_1 U1209 ( .A(n673), .X(n872) );
  SEN_ND2_S_0P5 U1210 ( .A1(net16193), .A2(net16134), .X(n715) );
  SEN_OAOI211_1 U1211 ( .A1(B[0]), .A2(A[0]), .B(n359), .C(n784), .X(net15997)
         );
  SEN_OAOI211_1 U1212 ( .A1(B[7]), .A2(A[7]), .B(net16444), .C(n779), .X(
        net16007) );
  SEN_ND2_S_0P5 U1213 ( .A1(net18219), .A2(n778), .X(net16006) );
  SEN_OR3B_0P5 U1214 ( .B1(n697), .B2(net16478), .A(n696), .X(n709) );
  SEN_ND2_S_0P5 U1215 ( .A1(net18219), .A2(net17000), .X(net16066) );
  SEN_ND2_S_0P5 U1216 ( .A1(net16434), .A2(n859), .X(net15818) );
  SEN_OAOI211_0P5 U1217 ( .A1(B[18]), .A2(A[18]), .B(net17584), .C(n844), .X(
        net15848) );
  SEN_ND2_S_0P5 U1218 ( .A1(n451), .A2(net16999), .X(net16145) );
  SEN_ND2_S_0P5 U1219 ( .A1(net16434), .A2(n856), .X(net15831) );
  SEN_OAOI211_1 U1220 ( .A1(B[23]), .A2(A[23]), .B(n359), .C(n877), .X(
        net15786) );
  SEN_ND2_S_0P5 U1221 ( .A1(net16434), .A2(net17005), .X(net15787) );
  SEN_OAOI211_1 U1222 ( .A1(B[1]), .A2(A[1]), .B(net17584), .C(n790), .X(
        net15988) );
  SEN_ND2_S_0P5 U1223 ( .A1(net18219), .A2(n793), .X(net15987) );
  SEN_ND2_S_0P5 U1224 ( .A1(net18219), .A2(net16084), .X(net16079) );
  SEN_ND2_S_0P5 U1225 ( .A1(net18219), .A2(net15973), .X(net15976) );
  SEN_OAOI211_0P5 U1226 ( .A1(B[11]), .A2(A[11]), .B(net16444), .C(n769), .X(
        net16030) );
  SEN_ND2_S_0P5 U1227 ( .A1(net18219), .A2(n766), .X(net16029) );
  SEN_ND2_S_0P5 U1228 ( .A1(net16434), .A2(n809), .X(net15920) );
  SEN_OAOI211_0P5 U1229 ( .A1(B[16]), .A2(A[16]), .B(net16444), .C(n812), .X(
        net15921) );
  SEN_ND2_S_0P5 U1230 ( .A1(net16434), .A2(n527), .X(net15870) );
  SEN_ND2_S_0P5 U1231 ( .A1(net16434), .A2(n805), .X(net15928) );
  SEN_MUXI2_S_0P5 U1232 ( .D0(n550), .D1(n511), .S(B[24]), .X(n678) );
  SEN_INV_1 U1233 ( .A(A[3]), .X(n545) );
  SEN_MUXI2_S_0P5 U1234 ( .D0(net16480), .D1(net16201), .S(A[27]), .X(n565) );
  SEN_MUXI2_S_0P5 U1235 ( .D0(net16482), .D1(net16201), .S(A[26]), .X(net16196) );
  SEN_INV_1 U1236 ( .A(B[18]), .X(n540) );
  SEN_MUXI2_S_0P5 U1237 ( .D0(net16480), .D1(n549), .S(A[21]), .X(n586) );
  SEN_MUXI2_S_0P5 U1238 ( .D0(n550), .D1(n367), .S(B[31]), .X(n699) );
  SEN_INV_S_1 U1239 ( .A(net15829), .X(net16345) );
  SEN_NR3_0P5 U1240 ( .A1(n789), .A2(n788), .A3(net16422), .X(n790) );
  SEN_NR3_0P5 U1241 ( .A1(n756), .A2(n755), .A3(net16772), .X(n757) );
  SEN_NR3_0P5 U1242 ( .A1(net15979), .A2(net15980), .A3(net16772), .X(n795) );
  SEN_NR3_0P5 U1243 ( .A1(net16020), .A2(net16021), .A3(net16772), .X(n774) );
  SEN_NR3_T_0P5 U1244 ( .A1(n853), .A2(n852), .A3(net16774), .X(n854) );
  SEN_NR3_0P5 U1245 ( .A1(n763), .A2(n762), .A3(net16772), .X(n764) );
  SEN_NR3_0P5 U1246 ( .A1(n836), .A2(n835), .A3(net16774), .X(n837) );
  SEN_NR3_0P5 U1247 ( .A1(n768), .A2(n767), .A3(net16772), .X(n769) );
  SEN_OR2_DG_1 U1248 ( .A1(n832), .A2(n758), .X(n528) );
  SEN_AO21B_1 U1249 ( .A1(n834), .A2(n831), .B(n760), .X(n529) );
  SEN_ND2_G_1 U1250 ( .A1(n717), .A2(n716), .X(n731) );
  SEN_EO2_S_0P5 U1251 ( .A1(n709), .A2(n707), .X(n705) );
  SEN_OA2BB2_0P5 U1252 ( .A1(n889), .A2(n888), .B1(n887), .B2(net16448), .X(
        net15763) );
  SEN_INV_S_1 U1253 ( .A(net16192), .X(net15790) );
  SEN_INV_S_1 U1254 ( .A(net16222), .X(net16069) );
  SEN_INV_S_1 U1255 ( .A(net16223), .X(net16070) );
  SEN_INV_S_1 U1256 ( .A(n701), .X(n707) );
  SEN_INV_S_1 U1257 ( .A(n577), .X(n739) );
  SEN_ND2_G_1 U1258 ( .A1(n565), .A2(n564), .X(n889) );
  SEN_INV_S_1 U1259 ( .A(n353), .X(n26) );
  SEN_OAOI211_G_1 U1260 ( .A1(B[9]), .A2(A[9]), .B(net16444), .C(n825), .X(
        net15886) );
  SEN_ND2_S_0P5 U1261 ( .A1(net16434), .A2(n523), .X(net15885) );
  SEN_OAOI211_G_1 U1262 ( .A1(B[10]), .A2(A[10]), .B(net16444), .C(n830), .X(
        net15871) );
  SEN_ND2_G_1 U1263 ( .A1(net18219), .A2(net15969), .X(net15964) );
  SEN_OAOI211_G_1 U1264 ( .A1(B[15]), .A2(A[15]), .B(net16444), .C(n819), .X(
        net15903) );
  SEN_EN2_S_1 U1265 ( .A1(n834), .A2(n833), .X(net15857) );
  SEN_ND2_G_1 U1266 ( .A1(net17602), .A2(n677), .X(net16192) );
  SEN_INV_S_1 U1267 ( .A(n352), .X(n28) );
  SEN_ND2_G_1 U1268 ( .A1(n568), .A2(n567), .X(n730) );
  SEN_MUXI2_S_0P5 U1269 ( .D0(net16480), .D1(net16201), .S(A[28]), .X(n568) );
  SEN_INV_S_1 U1270 ( .A(n354), .X(n24) );
  SEN_ND2_S_0P5 U1271 ( .A1(net18219), .A2(n814), .X(net16038) );
  SEN_OAOI211_G_1 U1272 ( .A1(B[12]), .A2(A[12]), .B(net17584), .C(n757), .X(
        net16053) );
  SEN_ND2_S_0P5 U1273 ( .A1(net18219), .A2(n360), .X(net16052) );
  SEN_ND2_G_1 U1274 ( .A1(n571), .A2(n570), .X(n725) );
  SEN_MUXI2_S_0P5 U1275 ( .D0(net16480), .D1(net16201), .S(A[29]), .X(n571) );
  SEN_INV_S_1 U1276 ( .A(n355), .X(n22) );
  SEN_MUXI2_S_0P5 U1277 ( .D0(net16480), .D1(net16201), .S(A[30]), .X(n574) );
  SEN_INV_S_1 U1278 ( .A(n356), .X(n20) );
  SEN_OR2_1 U1279 ( .A1(A[28]), .A2(B[28]), .X(n538) );
  SEN_NR2_1 U1280 ( .A1(A[27]), .A2(B[27]), .X(n887) );
  SEN_ND2_G_1 U1281 ( .A1(net17602), .A2(n584), .X(n671) );
  SEN_ND2_G_1 U1282 ( .A1(net17602), .A2(n599), .X(net16222) );
  SEN_MUXI2_S_0P5 U1283 ( .D0(net16480), .D1(n549), .S(A[22]), .X(n599) );
  SEN_ND2_G_1 U1284 ( .A1(n555), .A2(n687), .X(net16193) );
  SEN_ND2_G_1 U1285 ( .A1(n553), .A2(n569), .X(n576) );
  SEN_MUXI2_S_0P5 U1286 ( .D0(n550), .D1(n367), .S(B[29]), .X(n569) );
  SEN_ND2_G_1 U1287 ( .A1(n555), .A2(n566), .X(n575) );
  SEN_MUXI2_S_0P5 U1288 ( .D0(n550), .D1(n367), .S(B[28]), .X(n566) );
  SEN_ND2_G_1 U1289 ( .A1(n553), .A2(n572), .X(n577) );
  SEN_MUXI2_S_0P5 U1290 ( .D0(n550), .D1(n367), .S(B[30]), .X(n572) );
  SEN_ND2_G_1 U1291 ( .A1(n553), .A2(n562), .X(n580) );
  SEN_ND2_G_1 U1292 ( .A1(n555), .A2(n682), .X(n686) );
  SEN_ND2_G_1 U1293 ( .A1(n553), .A2(n585), .X(n673) );
  SEN_MUXI2_S_0P5 U1294 ( .D0(n550), .D1(n368), .S(B[21]), .X(n585) );
  SEN_ND2_S_0P5 U1295 ( .A1(n554), .A2(n676), .X(net16191) );
  SEN_ND2_G_1 U1296 ( .A1(n553), .A2(n598), .X(net16223) );
  SEN_MUXI2_S_0P5 U1297 ( .D0(n550), .D1(n367), .S(B[22]), .X(n598) );
  SEN_ND2B_S_0P5 U1298 ( .A(net16499), .B(A[26]), .X(n352) );
  SEN_ND2B_S_0P5 U1299 ( .A(net16499), .B(A[27]), .X(n353) );
  SEN_ND2B_S_0P5 U1300 ( .A(net16499), .B(A[28]), .X(n354) );
  SEN_ND2B_S_0P5 U1301 ( .A(net16499), .B(A[29]), .X(n355) );
  SEN_ND2B_S_0P5 U1302 ( .A(net16499), .B(A[30]), .X(n356) );
  SEN_NR3_0P5 U1303 ( .A1(n811), .A2(n810), .A3(net16772), .X(n812) );
  SEN_MUXI2_S_1 U1304 ( .D0(n688), .D1(n536), .S(n28), .X(net16197) );
  SEN_MUXI2_S_1 U1305 ( .D0(n688), .D1(n536), .S(n20), .X(n573) );
  SEN_MUXI2_S_1 U1306 ( .D0(n688), .D1(n536), .S(n22), .X(n570) );
  SEN_MUXI2_S_1 U1307 ( .D0(n688), .D1(n536), .S(n24), .X(n567) );
  SEN_MUXI2_S_1 U1308 ( .D0(n688), .D1(n536), .S(n26), .X(n564) );
  SEN_TIE0_1 U1309 ( .X(\*Logic0* ) );
  SEN_BUF_1 U1310 ( .A(n533), .X(n539) );
  SEN_BUF_1 U1311 ( .A(n703), .X(n542) );
  SEN_INV_S_0P5 U1312 ( .A(net16179), .X(net16178) );
  SEN_BUF_1 U1313 ( .A(net15941), .X(net16723) );
  SEN_MUXI2_S_0P5 U1314 ( .D0(net16200), .D1(n549), .S(A[23]), .X(n677) );
  SEN_INV_S_0P5 U1315 ( .A(n583), .X(n688) );
  SEN_ND3_S_0P5 U1316 ( .A1(net16311), .A2(net16968), .A3(n695), .X(n621) );
  SEN_INV_S_1 U1317 ( .A(net16774), .X(net16424) );
  SEN_OAI21_S_0P5 U1318 ( .A1(net18246), .A2(net16178), .B(A[31]), .X(n696) );
  SEN_ND2_G_1 U1319 ( .A1(net16434), .A2(net15953), .X(net15948) );
  SEN_ND2_S_0P65 U1320 ( .A1(net16434), .A2(net16701), .X(net15937) );
  SEN_NR3_0P5 U1321 ( .A1(n783), .A2(n782), .A3(net15769), .X(n784) );
  SEN_INV_S_1 U1322 ( .A(net16424), .X(net16422) );
endmodule

