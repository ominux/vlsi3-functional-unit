
module Alu ( Z, A, B, INST, FLAGS, CLOCK );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  output [3:0] FLAGS;
  input CLOCK;
  wire   \*Logic0* , n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882;
  wire   [31:0] A_qual;
  wire   [31:0] B_qual;
  wire   [3:0] INST_qual;
  assign FLAGS[3] = \*Logic0* ;

  SEN_FDPQ_4 \INST_qual_reg[3]  ( .D(INST[3]), .CK(CLOCK), .Q(INST_qual[3]) );
  SEN_FDPQ_4 \INST_qual_reg[2]  ( .D(INST[2]), .CK(CLOCK), .Q(INST_qual[2]) );
  SEN_FDPQ_4 \INST_qual_reg[1]  ( .D(INST[1]), .CK(CLOCK), .Q(INST_qual[1]) );
  SEN_FDPQ_4 \INST_qual_reg[0]  ( .D(INST[0]), .CK(CLOCK), .Q(INST_qual[0]) );
  SEN_FDPQ_D_1 \A_qual_reg[13]  ( .D(A[13]), .CK(CLOCK), .Q(A_qual[13]) );
  SEN_FDPQ_D_1 \A_qual_reg[26]  ( .D(A[26]), .CK(CLOCK), .Q(A_qual[26]) );
  SEN_FDPQ_D_1 \A_qual_reg[24]  ( .D(A[24]), .CK(CLOCK), .Q(A_qual[24]) );
  SEN_FDPQ_D_1 \A_qual_reg[23]  ( .D(A[23]), .CK(CLOCK), .Q(A_qual[23]) );
  SEN_FDPQ_D_1 \A_qual_reg[22]  ( .D(A[22]), .CK(CLOCK), .Q(A_qual[22]) );
  SEN_FDPQ_D_1 \A_qual_reg[21]  ( .D(A[21]), .CK(CLOCK), .Q(A_qual[21]) );
  SEN_FDPQ_D_1 \A_qual_reg[20]  ( .D(A[20]), .CK(CLOCK), .Q(A_qual[20]) );
  SEN_FDPQ_D_1 \A_qual_reg[19]  ( .D(A[19]), .CK(CLOCK), .Q(A_qual[19]) );
  SEN_FDPQ_D_1 \A_qual_reg[18]  ( .D(A[18]), .CK(CLOCK), .Q(A_qual[18]) );
  SEN_FDPQ_D_1 \A_qual_reg[17]  ( .D(A[17]), .CK(CLOCK), .Q(A_qual[17]) );
  SEN_FDPQ_D_1 \A_qual_reg[14]  ( .D(A[14]), .CK(CLOCK), .Q(A_qual[14]) );
  SEN_FDPQ_D_1 \A_qual_reg[3]  ( .D(A[3]), .CK(CLOCK), .Q(A_qual[3]) );
  SEN_FDPQ_D_1 \B_qual_reg[26]  ( .D(B[26]), .CK(CLOCK), .Q(B_qual[26]) );
  SEN_FDPQ_D_1 \B_qual_reg[24]  ( .D(B[24]), .CK(CLOCK), .Q(B_qual[24]) );
  SEN_FDPQ_D_1 \B_qual_reg[23]  ( .D(B[23]), .CK(CLOCK), .Q(B_qual[23]) );
  SEN_FDPQ_D_1 \B_qual_reg[22]  ( .D(B[22]), .CK(CLOCK), .Q(B_qual[22]) );
  SEN_FDPQ_D_1 \B_qual_reg[21]  ( .D(B[21]), .CK(CLOCK), .Q(B_qual[21]) );
  SEN_FDPQ_D_1 \B_qual_reg[20]  ( .D(B[20]), .CK(CLOCK), .Q(B_qual[20]) );
  SEN_FDPQ_D_1 \B_qual_reg[19]  ( .D(B[19]), .CK(CLOCK), .Q(B_qual[19]) );
  SEN_FDPQ_D_1 \B_qual_reg[18]  ( .D(B[18]), .CK(CLOCK), .Q(B_qual[18]) );
  SEN_FDPQ_D_1 \B_qual_reg[17]  ( .D(B[17]), .CK(CLOCK), .Q(B_qual[17]) );
  SEN_FDPQ_D_1 \B_qual_reg[14]  ( .D(B[14]), .CK(CLOCK), .Q(B_qual[14]) );
  SEN_FDPQ_D_1 \B_qual_reg[0]  ( .D(B[0]), .CK(CLOCK), .Q(B_qual[0]) );
  SEN_FDPQ_D_1 \A_qual_reg[8]  ( .D(A[8]), .CK(CLOCK), .Q(A_qual[8]) );
  SEN_FDPQ_D_1 \B_qual_reg[8]  ( .D(B[8]), .CK(CLOCK), .Q(B_qual[8]) );
  SEN_FDPQ_D_1 \B_qual_reg[13]  ( .D(B[13]), .CK(CLOCK), .Q(B_qual[13]) );
  SEN_FDPQ_D_1 \B_qual_reg[31]  ( .D(B[31]), .CK(CLOCK), .Q(B_qual[31]) );
  SEN_FDPQ_D_1 \B_qual_reg[30]  ( .D(B[30]), .CK(CLOCK), .Q(B_qual[30]) );
  SEN_FDPQ_D_1 \B_qual_reg[29]  ( .D(B[29]), .CK(CLOCK), .Q(B_qual[29]) );
  SEN_FDPQ_D_1 \B_qual_reg[28]  ( .D(B[28]), .CK(CLOCK), .Q(B_qual[28]) );
  SEN_FDPQ_D_1 \B_qual_reg[27]  ( .D(B[27]), .CK(CLOCK), .Q(B_qual[27]) );
  SEN_FDPQ_D_1 \B_qual_reg[25]  ( .D(B[25]), .CK(CLOCK), .Q(B_qual[25]) );
  SEN_FDPQ_D_1 \B_qual_reg[16]  ( .D(B[16]), .CK(CLOCK), .Q(B_qual[16]) );
  SEN_FDPQ_D_1 \B_qual_reg[15]  ( .D(B[15]), .CK(CLOCK), .Q(B_qual[15]) );
  SEN_FDPQ_D_1 \B_qual_reg[2]  ( .D(B[2]), .CK(CLOCK), .Q(B_qual[2]) );
  SEN_FDPQ_D_1 \B_qual_reg[5]  ( .D(B[5]), .CK(CLOCK), .Q(B_qual[5]) );
  SEN_FDPQ_D_1 \A_qual_reg[30]  ( .D(A[30]), .CK(CLOCK), .Q(A_qual[30]) );
  SEN_FDPQ_D_1 \A_qual_reg[29]  ( .D(A[29]), .CK(CLOCK), .Q(A_qual[29]) );
  SEN_FDPQ_D_1 \A_qual_reg[28]  ( .D(A[28]), .CK(CLOCK), .Q(A_qual[28]) );
  SEN_FDPQ_D_1 \A_qual_reg[27]  ( .D(A[27]), .CK(CLOCK), .Q(A_qual[27]) );
  SEN_FDPQ_D_1 \A_qual_reg[25]  ( .D(A[25]), .CK(CLOCK), .Q(A_qual[25]) );
  SEN_FDPQ_D_1 \A_qual_reg[16]  ( .D(A[16]), .CK(CLOCK), .Q(A_qual[16]) );
  SEN_FDPQ_D_1 \A_qual_reg[15]  ( .D(A[15]), .CK(CLOCK), .Q(A_qual[15]) );
  SEN_FDPQ_D_1 \A_qual_reg[2]  ( .D(A[2]), .CK(CLOCK), .Q(A_qual[2]) );
  SEN_FDPQ_D_1 \A_qual_reg[5]  ( .D(A[5]), .CK(CLOCK), .Q(A_qual[5]) );
  SEN_FDPQ_D_1 \A_qual_reg[1]  ( .D(A[1]), .CK(CLOCK), .Q(A_qual[1]) );
  SEN_FDPQ_D_1 \B_qual_reg[1]  ( .D(B[1]), .CK(CLOCK), .Q(B_qual[1]) );
  SEN_FDPQ_1 \A_qual_reg[9]  ( .D(A[9]), .CK(CLOCK), .Q(A_qual[9]) );
  SEN_FDPQ_1 \A_qual_reg[12]  ( .D(A[12]), .CK(CLOCK), .Q(A_qual[12]) );
  SEN_FDPQ_1 \B_qual_reg[12]  ( .D(B[12]), .CK(CLOCK), .Q(B_qual[12]) );
  SEN_FDPQ_4 \A_qual_reg[31]  ( .D(A[31]), .CK(CLOCK), .Q(A_qual[31]) );
  SEN_FDPQ_D_1 \A_qual_reg[0]  ( .D(A[0]), .CK(CLOCK), .Q(A_qual[0]) );
  SEN_FDPQ_1 \A_qual_reg[10]  ( .D(A[10]), .CK(CLOCK), .Q(A_qual[10]) );
  SEN_FDPQ_D_2 \B_qual_reg[10]  ( .D(B[10]), .CK(CLOCK), .Q(B_qual[10]) );
  SEN_FDPQ_D_1 \A_qual_reg[4]  ( .D(A[4]), .CK(CLOCK), .Q(A_qual[4]) );
  SEN_FDPQ_D_1 \B_qual_reg[11]  ( .D(B[11]), .CK(CLOCK), .Q(B_qual[11]) );
  SEN_FDPQ_D_1 \A_qual_reg[11]  ( .D(A[11]), .CK(CLOCK), .Q(A_qual[11]) );
  SEN_FDPQ_D_1 \B_qual_reg[7]  ( .D(B[7]), .CK(CLOCK), .Q(B_qual[7]) );
  SEN_FDPQ_D_1 \A_qual_reg[7]  ( .D(A[7]), .CK(CLOCK), .Q(A_qual[7]) );
  SEN_FDPQ_D_1 \B_qual_reg[9]  ( .D(B[9]), .CK(CLOCK), .Q(B_qual[9]) );
  SEN_FDPQ_D_1 \B_qual_reg[6]  ( .D(B[6]), .CK(CLOCK), .Q(B_qual[6]) );
  SEN_FDPQ_D_1 \A_qual_reg[6]  ( .D(A[6]), .CK(CLOCK), .Q(A_qual[6]) );
  SEN_FDPQ_D_1 \B_qual_reg[4]  ( .D(B[4]), .CK(CLOCK), .Q(B_qual[4]) );
  SEN_FDPQ_D_1 \B_qual_reg[3]  ( .D(B[3]), .CK(CLOCK), .Q(B_qual[3]) );
  SEN_ND2_S_6 U278 ( .A1(n799), .A2(n745), .X(n750) );
  SEN_ND2_T_1 U279 ( .A1(n321), .A2(A_qual[1]), .X(n268) );
  SEN_INV_6 U280 ( .A(n843), .X(n842) );
  SEN_EN2_8 U281 ( .A1(n846), .A2(n847), .X(n843) );
  SEN_ND3_1 U282 ( .A1(n873), .A2(n872), .A3(n871), .X(n874) );
  SEN_INV_S_6 U283 ( .A(n593), .X(n447) );
  SEN_EN2_DG_2 U284 ( .A1(n310), .A2(n559), .X(n566) );
  SEN_OAI211_2 U285 ( .A1(n566), .A2(n339), .B1(n565), .B2(n564), .X(Z[25]) );
  SEN_NR2_S_3 U286 ( .A1(Z[24]), .A2(Z[25]), .X(n861) );
  SEN_ND2_S_6 U287 ( .A1(n731), .A2(n732), .X(n405) );
  SEN_OAI22_3 U288 ( .A1(n647), .A2(n666), .B1(n646), .B2(n666), .X(n385) );
  SEN_ND2_T_2 U289 ( .A1(n710), .A2(n714), .X(n647) );
  SEN_ND2_T_4 U290 ( .A1(n559), .A2(n310), .X(n494) );
  SEN_ND2_2 U291 ( .A1(n854), .A2(n853), .X(n840) );
  SEN_ND2_T_3 U292 ( .A1(n325), .A2(n429), .X(n853) );
  SEN_ND2_T_4 U293 ( .A1(n255), .A2(n399), .X(n762) );
  SEN_ND2_2 U294 ( .A1(n240), .A2(n241), .X(n242) );
  SEN_ND2_T_1P5 U295 ( .A1(n203), .A2(n239), .X(n240) );
  SEN_NR2_T_1 U296 ( .A1(n727), .A2(n648), .X(n382) );
  SEN_ND2_2 U297 ( .A1(n279), .A2(n280), .X(n648) );
  SEN_ND2_T_1 U298 ( .A1(n786), .A2(n785), .X(n773) );
  SEN_ND2_T_2 U299 ( .A1(n290), .A2(n396), .X(n785) );
  SEN_ND2_S_0P5 U300 ( .A1(n744), .A2(n815), .X(n795) );
  SEN_NR2_G_1 U301 ( .A1(n744), .A2(n415), .X(n417) );
  SEN_ND2_2 U302 ( .A1(n810), .A2(n808), .X(n744) );
  SEN_ND2_T_5 U303 ( .A1(n494), .A2(n495), .X(n513) );
  SEN_NR2_T_3 U304 ( .A1(n494), .A2(n492), .X(n303) );
  SEN_ND2_T_1 U305 ( .A1(n321), .A2(A_qual[3]), .X(n232) );
  SEN_EN2_S_3 U306 ( .A1(n690), .A2(n689), .X(n666) );
  SEN_ND2_3 U307 ( .A1(n255), .A2(n374), .X(n690) );
  SEN_INV_4 U308 ( .A(n639), .X(n638) );
  SEN_EN2_3 U309 ( .A1(n641), .A2(n642), .X(n639) );
  SEN_ND2_T_4 U310 ( .A1(n324), .A2(n422), .X(n847) );
  SEN_ND2_T_4 U311 ( .A1(n254), .A2(n421), .X(n846) );
  SEN_OR2_5 U312 ( .A1(n303), .A2(n238), .X(n535) );
  SEN_INV_4 U313 ( .A(n200), .X(n203) );
  SEN_AN2_DG_4 U314 ( .A1(n279), .A2(n698), .X(n311) );
  SEN_AN2_3 U315 ( .A1(n405), .A2(n315), .X(n317) );
  SEN_INV_0P8 U316 ( .A(n405), .X(n710) );
  SEN_ND2_S_2 U317 ( .A1(A_qual[31]), .A2(INST_qual[2]), .X(n345) );
  SEN_ND2_2 U318 ( .A1(n324), .A2(n402), .X(n803) );
  SEN_MUXI2_DG_1 U319 ( .D0(n202), .D1(n320), .S(A_qual[15]), .X(n367) );
  SEN_INV_5 U320 ( .A(n323), .X(n320) );
  SEN_INV_2 U321 ( .A(n472), .X(n326) );
  SEN_MUXI2_S_3 U322 ( .D0(n330), .D1(n473), .S(B_qual[9]), .X(n378) );
  SEN_ND2_S_4 U323 ( .A1(n613), .A2(n289), .X(n438) );
  SEN_INV_S_3 U324 ( .A(n288), .X(n289) );
  SEN_INV_2P5 U325 ( .A(n341), .X(n474) );
  SEN_INV_S_6 U326 ( .A(n341), .X(n330) );
  SEN_INV_6 U327 ( .A(n458), .X(n200) );
  SEN_EN2_S_2 U328 ( .A1(n660), .A2(n661), .X(n658) );
  SEN_ND2_3 U329 ( .A1(n255), .A2(n366), .X(n660) );
  SEN_ND2_4 U330 ( .A1(n807), .A2(n810), .X(n745) );
  SEN_ND2B_V1DG_4 U331 ( .A(INST_qual[2]), .B(n346), .X(n467) );
  SEN_ND2_T_1P5 U332 ( .A1(n255), .A2(n244), .X(n851) );
  SEN_ND2_3 U333 ( .A1(n255), .A2(n378), .X(n738) );
  SEN_ND2_6 U334 ( .A1(n255), .A2(n370), .X(n731) );
  SEN_INV_3 U335 ( .A(n332), .X(n255) );
  SEN_MUXI2_S_2 U336 ( .D0(n474), .D1(n473), .S(B_qual[12]), .X(n376) );
  SEN_MUXI2_S_0P5 U337 ( .D0(n474), .D1(n473), .S(B_qual[14]), .X(n368) );
  SEN_INV_6 U338 ( .A(n473), .X(n329) );
  SEN_AO21B_6 U339 ( .A1(n480), .A2(n484), .B(n428), .X(n473) );
  SEN_ND2_T_2 U340 ( .A1(INST_qual[3]), .A2(INST_qual[0]), .X(n346) );
  SEN_INV_S_6 U341 ( .A(n416), .X(n764) );
  SEN_AOI211_G_2 U342 ( .A1(n793), .A2(n432), .B1(n417), .B2(n416), .X(n418)
         );
  SEN_ND2_S_4 U343 ( .A1(n223), .A2(n224), .X(n416) );
  SEN_ND2B_3 U344 ( .A(INST_qual[2]), .B(INST_qual[3]), .X(n342) );
  SEN_INV_3 U345 ( .A(INST_qual[0]), .X(n480) );
  SEN_OAI21_3 U346 ( .A1(n684), .A2(n681), .B(n705), .X(n380) );
  SEN_INV_S_8 U347 ( .A(n200), .X(n202) );
  SEN_INV_S_2 U348 ( .A(n731), .X(n261) );
  SEN_ND2_2 U349 ( .A1(n731), .A2(n262), .X(n263) );
  SEN_EO2_3 U350 ( .A1(n430), .A2(n853), .X(n852) );
  SEN_INV_S_6 U351 ( .A(n833), .X(n832) );
  SEN_EN2_S_3 U352 ( .A1(n835), .A2(n836), .X(n833) );
  SEN_ND2_T_4 U353 ( .A1(n714), .A2(n305), .X(n646) );
  SEN_INV_2 U354 ( .A(n658), .X(n215) );
  SEN_ND3_T_4 U355 ( .A1(n468), .A2(n347), .A3(n467), .X(n457) );
  SEN_ND2_S_1P5 U356 ( .A1(n517), .A2(n516), .X(n259) );
  SEN_ND2_S_4 U357 ( .A1(n496), .A2(n513), .X(n525) );
  SEN_INV_4 U358 ( .A(n432), .X(n815) );
  SEN_ND2_S_4 U359 ( .A1(n286), .A2(n287), .X(n432) );
  SEN_ND2_T_1P5 U360 ( .A1(n486), .A2(n299), .X(n300) );
  SEN_ND2_T_4 U361 ( .A1(n255), .A2(n409), .X(n821) );
  SEN_INV_4 U362 ( .A(n228), .X(n409) );
  SEN_NR2_4 U363 ( .A1(n307), .A2(n809), .X(n434) );
  SEN_NR2B_V1DG_6 U364 ( .A(n828), .B(n827), .X(n307) );
  SEN_AOI21_G_2 U365 ( .A1(n624), .A2(n614), .B(n609), .X(n393) );
  SEN_EN2_1 U366 ( .A1(n618), .A2(n617), .X(n609) );
  SEN_ND2_3 U367 ( .A1(n633), .A2(n197), .X(n610) );
  SEN_ND2_3 U368 ( .A1(n698), .A2(n276), .X(n715) );
  SEN_ND2_T_2 U369 ( .A1(n274), .A2(n275), .X(n276) );
  SEN_MUXI2_DG_3 U370 ( .D0(n201), .D1(n320), .S(A_qual[11]), .X(n373) );
  SEN_ND2_T_4 U371 ( .A1(n815), .A2(n832), .X(n752) );
  SEN_INV_S_8 U372 ( .A(n854), .X(n430) );
  SEN_AN2_S_2 U373 ( .A1(n406), .A2(n309), .X(n313) );
  SEN_ND2_2 U374 ( .A1(n324), .A2(n414), .X(n836) );
  SEN_OAI211_3 U375 ( .A1(n385), .A2(n384), .B1(n676), .B2(n383), .X(n633) );
  SEN_OA21B_8 U376 ( .A1(n447), .A2(n592), .B(n209), .X(n208) );
  SEN_ND2_S_1 U377 ( .A1(n726), .A2(n405), .X(n681) );
  SEN_OAI21_G_1 U378 ( .A1(n311), .A2(n666), .B(n406), .X(n384) );
  SEN_MUXI2_S_3 U379 ( .D0(n330), .D1(n327), .S(B_qual[4]), .X(n411) );
  SEN_ND2_3 U380 ( .A1(n255), .A2(n411), .X(n813) );
  SEN_ND2_4 U381 ( .A1(n828), .A2(n829), .X(n754) );
  SEN_ND2_4 U382 ( .A1(n842), .A2(n431), .X(n829) );
  SEN_INV_S_0P5 U383 ( .A(n681), .X(n683) );
  SEN_NR3_T_0P5 U384 ( .A1(n681), .A2(n740), .A3(n684), .X(n667) );
  SEN_INV_S_3 U385 ( .A(n813), .X(n284) );
  SEN_AN2_S_4 U386 ( .A1(n311), .A2(n317), .X(n309) );
  SEN_MUXI2_DG_3 U387 ( .D0(n203), .D1(n320), .S(A_qual[12]), .X(n377) );
  SEN_ND2_4 U388 ( .A1(n762), .A2(n761), .X(n723) );
  SEN_ND2_2 U389 ( .A1(n256), .A2(n376), .X(n703) );
  SEN_ND2_2 U390 ( .A1(n256), .A2(n413), .X(n835) );
  SEN_ND2_S_4 U391 ( .A1(n703), .A2(n702), .X(n279) );
  SEN_INV_S_3 U392 ( .A(n702), .X(n278) );
  SEN_ND2_S_3 U393 ( .A1(n324), .A2(n377), .X(n702) );
  SEN_ND2_3 U394 ( .A1(n324), .A2(n379), .X(n737) );
  SEN_MUXI2_DG_3 U395 ( .D0(n201), .D1(n320), .S(A_qual[9]), .X(n379) );
  SEN_ND2_T_1 U396 ( .A1(n504), .A2(n506), .X(n293) );
  SEN_ND2_S_4 U397 ( .A1(n493), .A2(n258), .X(n260) );
  SEN_INV_S_6 U398 ( .A(n516), .X(n258) );
  SEN_OAI21_3 U399 ( .A1(n503), .A2(n502), .B(n501), .X(n504) );
  SEN_MUXI2_DG_5 U400 ( .D0(n330), .D1(n327), .S(B_qual[8]), .X(n399) );
  SEN_ND2_2 U401 ( .A1(n477), .A2(n478), .X(n301) );
  SEN_OAI211_3 U402 ( .A1(n542), .A2(n339), .B1(n541), .B2(n540), .X(Z[27]) );
  SEN_OAI21_S_8 U403 ( .A1(n208), .A2(n584), .B(n450), .X(n576) );
  SEN_ND2_T_4 U404 ( .A1(n852), .A2(n840), .X(n827) );
  SEN_INV_2 U405 ( .A(n408), .X(n613) );
  SEN_INV_S_3 U406 ( .A(n722), .X(n407) );
  SEN_ND2_T_1 U407 ( .A1(n627), .A2(n626), .X(n614) );
  SEN_ND2_3 U408 ( .A1(n480), .A2(n343), .X(n428) );
  SEN_ND2_G_1 U409 ( .A1(n690), .A2(n689), .X(n406) );
  SEN_ND2_2 U410 ( .A1(n614), .A2(n611), .X(n394) );
  SEN_ND2_T_1P5 U411 ( .A1(n813), .A2(n812), .X(n793) );
  SEN_EN2_S_2 U412 ( .A1(n802), .A2(n803), .X(n800) );
  SEN_EN2_3 U413 ( .A1(n778), .A2(n779), .X(n776) );
  SEN_ND2_G_1 U414 ( .A1(n778), .A2(n779), .X(n748) );
  SEN_ND2_2 U415 ( .A1(n221), .A2(n222), .X(n224) );
  SEN_ND2_G_2 U416 ( .A1(n738), .A2(n737), .X(n726) );
  SEN_ND2_G_1 U417 ( .A1(n277), .A2(n278), .X(n280) );
  SEN_ND2_2 U418 ( .A1(n251), .A2(n252), .X(n651) );
  SEN_ND2_G_1 U419 ( .A1(n249), .A2(n250), .X(n252) );
  SEN_EN2_0P5 U420 ( .A1(n627), .A2(n626), .X(n624) );
  SEN_NR2_T_2 U421 ( .A1(n610), .A2(n394), .X(n440) );
  SEN_ND2_S_3 U422 ( .A1(n696), .A2(n437), .X(n288) );
  SEN_AN2_S_1 U423 ( .A1(n578), .A2(n577), .X(n211) );
  SEN_OR2_1 U424 ( .A1(n302), .A2(n304), .X(n238) );
  SEN_ND2_G_2 U425 ( .A1(n291), .A2(n292), .X(n294) );
  SEN_INV_2 U426 ( .A(n504), .X(n292) );
  SEN_INV_2 U427 ( .A(Z[31]), .X(n881) );
  SEN_INV_S_1 U428 ( .A(n793), .X(n415) );
  SEN_INV_1 U429 ( .A(n761), .X(n222) );
  SEN_INV_S_3 U430 ( .A(n709), .X(n436) );
  SEN_ND2_G_1 U431 ( .A1(n536), .A2(n547), .X(n515) );
  SEN_INV_S_4 U432 ( .A(n754), .X(n809) );
  SEN_ND2_T_1 U433 ( .A1(n821), .A2(n820), .X(n272) );
  SEN_INV_S_1 U434 ( .A(n820), .X(n271) );
  SEN_ND2_G_1 U435 ( .A1(n330), .A2(n225), .X(n226) );
  SEN_ND2_G_1 U436 ( .A1(n793), .A2(n795), .X(n747) );
  SEN_ND2_G_1 U437 ( .A1(n775), .A2(n420), .X(n749) );
  SEN_ND2_G_1 U438 ( .A1(n474), .A2(n245), .X(n246) );
  SEN_INV_S_1 U439 ( .A(n718), .X(n275) );
  SEN_ND2_2 U440 ( .A1(n717), .A2(n718), .X(n698) );
  SEN_AN2_3 U441 ( .A1(n726), .A2(n723), .X(n315) );
  SEN_INV_S_1 U442 ( .A(n698), .X(n684) );
  SEN_INV_S_1 U443 ( .A(n406), .X(n669) );
  SEN_INV_S_1 U444 ( .A(n390), .X(n634) );
  SEN_AN2_3 U445 ( .A1(n253), .A2(n313), .X(n318) );
  SEN_ND2_G_4 U446 ( .A1(n216), .A2(n403), .X(n722) );
  SEN_OAI21_G_2 U447 ( .A1(n312), .A2(n776), .B(n748), .X(n403) );
  SEN_ND2_G_1 U448 ( .A1(n641), .A2(n642), .X(n611) );
  SEN_OA21_1 U449 ( .A1(n634), .A2(n215), .B(n638), .X(n308) );
  SEN_INV_S_8 U450 ( .A(n323), .X(n321) );
  SEN_AN2_S_1 U451 ( .A1(n569), .A2(n568), .X(n206) );
  SEN_ND3_1 U452 ( .A1(n866), .A2(n865), .A3(n864), .X(n876) );
  SEN_MUXI2_D_1 U453 ( .D0(n201), .D1(n321), .S(A_qual[2]), .X(n414) );
  SEN_ND2_2 U454 ( .A1(n226), .A2(n227), .X(n228) );
  SEN_ND2_2 U455 ( .A1(n327), .A2(B_qual[3]), .X(n227) );
  SEN_INV_2 U456 ( .A(n800), .X(n799) );
  SEN_MUXI2_S_1 U457 ( .D0(n201), .D1(n321), .S(A_qual[5]), .X(n402) );
  SEN_INV_2 U458 ( .A(n776), .X(n775) );
  SEN_INV_S_1 U459 ( .A(n727), .X(n740) );
  SEN_INV_3 U460 ( .A(n715), .X(n714) );
  SEN_INV_2 U461 ( .A(n648), .X(n705) );
  SEN_INV_2 U462 ( .A(n651), .X(n676) );
  SEN_ND2_G_1 U463 ( .A1(n324), .A2(n369), .X(n673) );
  SEN_ND2_G_1 U464 ( .A1(n255), .A2(n368), .X(n674) );
  SEN_ND2_G_1 U465 ( .A1(n290), .A2(n367), .X(n661) );
  SEN_ND2_G_1 U466 ( .A1(n256), .A2(n388), .X(n641) );
  SEN_MUXI2_S_1 U467 ( .D0(n330), .D1(n327), .S(B_qual[16]), .X(n388) );
  SEN_ND2_2 U468 ( .A1(n220), .A2(n393), .X(n439) );
  SEN_ND2_G_1 U469 ( .A1(n256), .A2(n443), .X(n603) );
  SEN_EN2_0P5 U470 ( .A1(n305), .A2(n728), .X(n735) );
  SEN_EN2_1 U471 ( .A1(n536), .A2(n535), .X(n542) );
  SEN_OAI211_2 U472 ( .A1(n534), .A2(n339), .B1(n533), .B2(n532), .X(Z[29]) );
  SEN_EN2_1 U473 ( .A1(n527), .A2(n526), .X(n534) );
  SEN_OAI211_3 U474 ( .A1(n512), .A2(n338), .B1(n511), .B2(n510), .X(Z[30]) );
  SEN_ND2_T_2 U475 ( .A1(n229), .A2(n198), .X(Z[31]) );
  SEN_ND2_G_1 U476 ( .A1(n762), .A2(n761), .X(n223) );
  SEN_INV_S_1 U477 ( .A(n762), .X(n221) );
  SEN_INV_S_0P5 U478 ( .A(n453), .X(n196) );
  SEN_ND2_T_2 U479 ( .A1(n300), .A2(n301), .X(n490) );
  SEN_AN2_S_1 U480 ( .A1(n253), .A2(n390), .X(n197) );
  SEN_INV_2 U481 ( .A(n478), .X(n299) );
  SEN_AN3_1 U482 ( .A1(n489), .A2(n488), .A3(n487), .X(n198) );
  SEN_INV_S_2 U483 ( .A(n326), .X(n290) );
  SEN_INV_S_1 U484 ( .A(n493), .X(n517) );
  SEN_ND2_G_1 U485 ( .A1(n696), .A2(n281), .X(n724) );
  SEN_AN2_S_1 U486 ( .A1(n524), .A2(n314), .X(n199) );
  SEN_INV_S_1 U487 ( .A(n513), .X(n543) );
  SEN_INV_3 U488 ( .A(n423), .X(n343) );
  SEN_AN2_2 U489 ( .A1(n770), .A2(n773), .X(n312) );
  SEN_ND2_G_1 U490 ( .A1(n802), .A2(n803), .X(n770) );
  SEN_ND2B_3 U491 ( .A(INST_qual[2]), .B(INST_qual[1]), .X(n423) );
  SEN_ND2_3 U492 ( .A1(n293), .A2(n294), .X(n512) );
  SEN_INV_S_8 U493 ( .A(n200), .X(n201) );
  SEN_OAI211_8 U494 ( .A1(n523), .A2(n339), .B1(n522), .B2(n521), .X(Z[28]) );
  SEN_ND2_6 U495 ( .A1(n259), .A2(n260), .X(n523) );
  SEN_ND2_G_3 U496 ( .A1(n324), .A2(n398), .X(n779) );
  SEN_INV_2 U497 ( .A(n329), .X(n328) );
  SEN_INV_12 U498 ( .A(n329), .X(n327) );
  SEN_BUF_1 U499 ( .A(n196), .X(n204) );
  SEN_INV_4 U500 ( .A(n576), .X(n453) );
  SEN_INV_S_3 U501 ( .A(Z[30]), .X(n880) );
  SEN_OA21B_4 U502 ( .A1(n210), .A2(n567), .B(n206), .X(n205) );
  SEN_BUF_1 U503 ( .A(n593), .X(n207) );
  SEN_AN2_DG_16 U504 ( .A1(n595), .A2(n594), .X(n209) );
  SEN_OA21B_4 U505 ( .A1(n453), .A2(n575), .B(n211), .X(n210) );
  SEN_INV_S_0P5 U506 ( .A(n210), .X(n212) );
  SEN_INV_S_0P5 U507 ( .A(n205), .X(n213) );
  SEN_INV_S_0P5 U508 ( .A(n208), .X(n214) );
  SEN_ND2_G_3 U509 ( .A1(n272), .A2(n273), .X(n807) );
  SEN_ND2_T_2 U510 ( .A1(n270), .A2(n271), .X(n273) );
  SEN_INV_1P25 U511 ( .A(n821), .X(n270) );
  SEN_OAI21_S_0P5 U512 ( .A1(n667), .A2(n648), .B(n279), .X(n649) );
  SEN_INV_0P8 U513 ( .A(n703), .X(n277) );
  SEN_INV_4 U514 ( .A(n342), .X(n484) );
  SEN_NR2_S_8 U515 ( .A1(n430), .A2(n429), .X(n282) );
  SEN_INV_5 U516 ( .A(n298), .X(n429) );
  SEN_ND2_3 U517 ( .A1(n296), .A2(n297), .X(n298) );
  SEN_INV_4 U518 ( .A(n269), .X(n422) );
  SEN_ND2_3 U519 ( .A1(n267), .A2(n268), .X(n269) );
  SEN_ND2_T_1P5 U520 ( .A1(n201), .A2(n266), .X(n267) );
  SEN_INV_2 U521 ( .A(n812), .X(n285) );
  SEN_ND2_G_1 U522 ( .A1(n835), .A2(n836), .X(n808) );
  SEN_INV_6 U523 ( .A(n457), .X(n323) );
  SEN_INV_4 U524 ( .A(n242), .X(n412) );
  SEN_ND2_4 U525 ( .A1(n324), .A2(n412), .X(n812) );
  SEN_ND2_G_2 U526 ( .A1(n846), .A2(n847), .X(n828) );
  SEN_ND2_T_4 U527 ( .A1(n290), .A2(n410), .X(n820) );
  SEN_INV_3 U528 ( .A(n233), .X(n410) );
  SEN_INV_S_0P5 U529 ( .A(n807), .X(n823) );
  SEN_ND2_0P8 U530 ( .A1(n325), .A2(n387), .X(n626) );
  SEN_OR3B_4 U531 ( .B1(A_qual[31]), .B2(INST_qual[3]), .A(n480), .X(n347) );
  SEN_ND2_0P8 U532 ( .A1(n525), .A2(n199), .X(n526) );
  SEN_ND2_3 U533 ( .A1(n256), .A2(n395), .X(n786) );
  SEN_EN2_S_3 U534 ( .A1(n786), .A2(n785), .X(n783) );
  SEN_MUXI2_DG_3 U535 ( .D0(n330), .D1(n327), .S(B_qual[1]), .X(n421) );
  SEN_ND2_T_3 U536 ( .A1(n325), .A2(n400), .X(n761) );
  SEN_ND2_S_3 U537 ( .A1(n821), .A2(n820), .X(n810) );
  SEN_MUXI2_DG_2 U538 ( .D0(n203), .D1(n320), .S(A_qual[10]), .X(n371) );
  SEN_ND3B_1 U539 ( .A(n346), .B1(INST_qual[1]), .B2(INST_qual[2]), .X(n472)
         );
  SEN_INV_5 U540 ( .A(n326), .X(n324) );
  SEN_NR2_T_6 U541 ( .A1(n750), .A2(n751), .X(n435) );
  SEN_OAI21_S_0P5 U542 ( .A1(n736), .A2(n727), .B(n726), .X(n728) );
  SEN_INV_S_0P5 U543 ( .A(n726), .X(n697) );
  SEN_OAI31_3 U544 ( .A1(n345), .A2(INST_qual[0]), .A3(INST_qual[3]), .B(n466), 
        .X(n458) );
  SEN_ND2_4 U545 ( .A1(n263), .A2(n264), .X(n305) );
  SEN_INV_S_3 U546 ( .A(n420), .X(n751) );
  SEN_ND2_6 U547 ( .A1(n255), .A2(n425), .X(n854) );
  SEN_MUXI2_DG_8 U548 ( .D0(n424), .D1(n327), .S(B_qual[0]), .X(n425) );
  SEN_OR4B_4 U549 ( .B1(n382), .B2(n669), .B3(n381), .A(n380), .X(n383) );
  SEN_OR2_2 U550 ( .A1(n423), .A2(n480), .X(n235) );
  SEN_OA21_2 U551 ( .A1(n420), .A2(n404), .B(n764), .X(n216) );
  SEN_ND2_S_4 U552 ( .A1(n773), .A2(n783), .X(n420) );
  SEN_INV_S_1 U553 ( .A(n748), .X(n404) );
  SEN_AN3B_8 U554 ( .B1(n775), .B2(n764), .A(n752), .X(n433) );
  SEN_MUXI2_DG_2 U555 ( .D0(n201), .D1(n321), .S(A_qual[6]), .X(n396) );
  SEN_ND3_T_4 U556 ( .A1(n435), .A2(n434), .A3(n433), .X(n709) );
  SEN_MUXI2_DG_3 U557 ( .D0(n202), .D1(n321), .S(A_qual[8]), .X(n400) );
  SEN_AOI31_0P75 U558 ( .A1(n807), .A2(n793), .A3(n810), .B(n800), .X(n419) );
  SEN_ND3_S_4 U559 ( .A1(n419), .A2(n759), .A3(n418), .X(n696) );
  SEN_ND2_S_0P5 U560 ( .A1(n793), .A2(n794), .X(n746) );
  SEN_INV_2 U561 ( .A(n326), .X(n325) );
  SEN_INV_S_0P5 U562 ( .A(n666), .X(n692) );
  SEN_ND2_S_4 U563 ( .A1(n525), .A2(n500), .X(n503) );
  SEN_ND2_T_6 U564 ( .A1(n237), .A2(n514), .X(n516) );
  SEN_INV_S_2 U565 ( .A(Z[18]), .X(n865) );
  SEN_AOAI211_1 U566 ( .A1(n613), .A2(n653), .B(n612), .C(n611), .X(n625) );
  SEN_ND3_S_0P5 U567 ( .A1(n435), .A2(n433), .A3(n434), .X(n281) );
  SEN_MUXI2_S_2 U568 ( .D0(n202), .D1(n321), .S(A_qual[7]), .X(n398) );
  SEN_ND2_T_1 U569 ( .A1(n321), .A2(A_qual[0]), .X(n297) );
  SEN_ND2_T_2 U570 ( .A1(n256), .A2(n397), .X(n778) );
  SEN_BUF_2 U571 ( .A(n476), .X(n256) );
  SEN_AN2_6 U572 ( .A1(n442), .A2(n441), .X(n217) );
  SEN_INV_S_2 U573 ( .A(Z[29]), .X(n882) );
  SEN_EO2_1 U574 ( .A1(n547), .A2(n543), .X(n550) );
  SEN_OR4B_4 U575 ( .B1(Z[27]), .B2(Z[26]), .B3(Z[28]), .A(n878), .X(n879) );
  SEN_OAOI211_1 U576 ( .A1(n636), .A2(n724), .B(n635), .C(n634), .X(n637) );
  SEN_ND2_2 U577 ( .A1(n218), .A2(n219), .X(n220) );
  SEN_INV_2 U578 ( .A(n308), .X(n218) );
  SEN_INV_S_0P5 U579 ( .A(n394), .X(n219) );
  SEN_ND2_T_1 U580 ( .A1(n201), .A2(n295), .X(n296) );
  SEN_INV_S_0P5 U581 ( .A(n745), .X(n794) );
  SEN_OR3B_4 U582 ( .B1(n440), .B2(n439), .A(n438), .X(n442) );
  SEN_MUXI2_DG_2 U583 ( .D0(n203), .D1(n320), .S(A_qual[13]), .X(n375) );
  SEN_ND2_G_1 U584 ( .A1(n813), .A2(n812), .X(n286) );
  SEN_ND2_T_2 U585 ( .A1(n325), .A2(n375), .X(n689) );
  SEN_ND2_2 U586 ( .A1(n261), .A2(n732), .X(n264) );
  SEN_OR3B_4 U587 ( .B1(n407), .B2(n634), .A(n318), .X(n408) );
  SEN_ND2_T_2 U588 ( .A1(n254), .A2(n372), .X(n717) );
  SEN_MUXI2_DG_3 U589 ( .D0(n474), .D1(n327), .S(B_qual[11]), .X(n372) );
  SEN_ND2_S_1P5 U590 ( .A1(n674), .A2(n673), .X(n654) );
  SEN_BUF_S_3 U591 ( .A(n654), .X(n253) );
  SEN_ND2_2 U592 ( .A1(n284), .A2(n285), .X(n287) );
  SEN_AO2BB2_8 U593 ( .A1(n217), .A2(n601), .B1(n603), .B2(n602), .X(n593) );
  SEN_AN4B_2 U594 ( .B1(n880), .B2(n882), .B3(n881), .A(n879), .X(FLAGS[2]) );
  SEN_NR4_6 U595 ( .A1(n877), .A2(n876), .A3(n875), .A4(n874), .X(n878) );
  SEN_ND3_S_4 U596 ( .A1(n863), .A2(n862), .A3(n861), .X(n877) );
  SEN_MUXI2_DG_3 U597 ( .D0(n330), .D1(n327), .S(B_qual[5]), .X(n401) );
  SEN_AN3B_4 U598 ( .B1(n611), .B2(n614), .A(n436), .X(n437) );
  SEN_OR2_5 U599 ( .A1(n282), .A2(n283), .X(n431) );
  SEN_MUXI2_DG_3 U600 ( .D0(n330), .D1(n327), .S(B_qual[6]), .X(n395) );
  SEN_MUXI2_DG_2 U601 ( .D0(n330), .D1(n327), .S(B_qual[2]), .X(n413) );
  SEN_OAI211_2 U602 ( .A1(n550), .A2(n339), .B1(n549), .B2(n548), .X(Z[26]) );
  SEN_MUXI2_DG_2 U603 ( .D0(n330), .D1(n327), .S(B_qual[7]), .X(n397) );
  SEN_MUXI2_DG_3 U604 ( .D0(n474), .D1(n328), .S(B_qual[15]), .X(n366) );
  SEN_ND2_3 U605 ( .A1(n325), .A2(n371), .X(n732) );
  SEN_INV_0P5 U606 ( .A(B_qual[3]), .X(n225) );
  SEN_ND2_T_2 U607 ( .A1(n490), .A2(n505), .X(n229) );
  SEN_ND2_T_1 U608 ( .A1(n201), .A2(n230), .X(n231) );
  SEN_ND2_2 U609 ( .A1(n231), .A2(n232), .X(n233) );
  SEN_INV_S_1 U610 ( .A(A_qual[3]), .X(n230) );
  SEN_OR2_DG_1 U611 ( .A1(n479), .A2(INST_qual[3]), .X(n234) );
  SEN_ND2_2 U612 ( .A1(n234), .A2(n235), .X(n424) );
  SEN_ND2_T_4 U613 ( .A1(n513), .A2(n236), .X(n237) );
  SEN_INV_4 U614 ( .A(n515), .X(n236) );
  SEN_NR2_6 U615 ( .A1(n316), .A2(n319), .X(n514) );
  SEN_ND2_T_2 U616 ( .A1(n321), .A2(A_qual[4]), .X(n241) );
  SEN_INV_1 U617 ( .A(A_qual[4]), .X(n239) );
  SEN_ND2_S_0P5 U618 ( .A1(n428), .A2(n427), .X(n243) );
  SEN_INV_1 U619 ( .A(n243), .X(n244) );
  SEN_INV_2 U620 ( .A(n851), .X(n283) );
  SEN_ND2_G_0P65 U621 ( .A1(n660), .A2(n661), .X(n390) );
  SEN_ND2_T_3 U622 ( .A1(n327), .A2(B_qual[10]), .X(n247) );
  SEN_ND2_4 U623 ( .A1(n246), .A2(n247), .X(n248) );
  SEN_INV_1 U624 ( .A(B_qual[10]), .X(n245) );
  SEN_INV_S_6 U625 ( .A(n248), .X(n370) );
  SEN_ND2_S_1 U626 ( .A1(n674), .A2(n673), .X(n251) );
  SEN_INV_0P65 U627 ( .A(n674), .X(n249) );
  SEN_INV_S_0P5 U628 ( .A(n673), .X(n250) );
  SEN_MUXI2_DG_2 U629 ( .D0(n474), .D1(n327), .S(B_qual[13]), .X(n374) );
  SEN_ND2_T_2 U630 ( .A1(n256), .A2(n401), .X(n802) );
  SEN_OR3B_2 U631 ( .B1(INST_qual[1]), .B2(INST_qual[0]), .A(INST_qual[3]), 
        .X(n468) );
  SEN_ND2_2 U632 ( .A1(INST_qual[0]), .A2(INST_qual[1]), .X(n479) );
  SEN_ND2_2 U633 ( .A1(n324), .A2(n373), .X(n718) );
  SEN_EN2_DG_4 U634 ( .A1(n738), .A2(n737), .X(n727) );
  SEN_OR4B_4 U635 ( .B1(n465), .B2(n464), .B3(n463), .A(n462), .X(n478) );
  SEN_OR4B_4 U636 ( .B1(n493), .B2(n461), .B3(n491), .A(n535), .X(n462) );
  SEN_INV_1 U637 ( .A(n749), .X(n759) );
  SEN_OAI21_S_0P5 U638 ( .A1(n784), .A2(n783), .B(n773), .X(n774) );
  SEN_INV_S_0P5 U639 ( .A(n783), .X(n788) );
  SEN_ND2_G_1 U640 ( .A1(n254), .A2(n386), .X(n627) );
  SEN_ND2_G_1 U641 ( .A1(n324), .A2(n389), .X(n642) );
  SEN_OR3B_0P5 U642 ( .B1(INST_qual[1]), .B2(INST_qual[0]), .A(n484), .X(n561)
         );
  SEN_ND2_S_0P5 U643 ( .A1(n723), .A2(n722), .X(n725) );
  SEN_ND2_S_0P5 U644 ( .A1(n722), .A2(n696), .X(n711) );
  SEN_NR2_S_0P5 U645 ( .A1(n844), .A2(n833), .X(n834) );
  SEN_INV_1 U646 ( .A(n717), .X(n274) );
  SEN_NR3_0P5 U647 ( .A1(n755), .A2(n792), .A3(n307), .X(n756) );
  SEN_ND2B_S_0P5 U648 ( .A(n307), .B(n768), .X(n771) );
  SEN_NR3_0P5 U649 ( .A1(n792), .A2(n307), .A3(n794), .X(n797) );
  SEN_OAI21_S_8 U650 ( .A1(n205), .A2(n551), .B(n460), .X(n559) );
  SEN_ND3B_2 U651 ( .A(INST_qual[1]), .B1(INST_qual[0]), .B2(INST_qual[2]), 
        .X(n466) );
  SEN_ND2_G_1 U652 ( .A1(n290), .A2(n444), .X(n602) );
  SEN_ND2_S_0P5 U653 ( .A1(n290), .A2(n459), .X(n552) );
  SEN_INV_1 U654 ( .A(n332), .X(n254) );
  SEN_OR3B_1 U655 ( .B1(INST_qual[1]), .B2(INST_qual[2]), .A(INST_qual[0]), 
        .X(n476) );
  SEN_INV_S_2 U656 ( .A(n476), .X(n332) );
  SEN_INV_S_1 U657 ( .A(n844), .X(n257) );
  SEN_OR3B_0P5 U658 ( .B1(n485), .B2(INST_qual[0]), .A(n484), .X(n844) );
  SEN_INV_1 U659 ( .A(n732), .X(n262) );
  SEN_ND2_S_0P5 U660 ( .A1(n842), .A2(n431), .X(n265) );
  SEN_INV_S_1 U661 ( .A(A_qual[1]), .X(n266) );
  SEN_INV_1 U662 ( .A(n625), .X(n615) );
  SEN_NR3_0P5 U663 ( .A1(n538), .A2(n561), .A3(n537), .X(n539) );
  SEN_EN2_0P5 U664 ( .A1(n508), .A2(n509), .X(n506) );
  SEN_INV_1 U665 ( .A(n491), .X(n536) );
  SEN_ND2_T_0P5 U666 ( .A1(n517), .A2(n316), .X(n524) );
  SEN_INV_S_0P5 U667 ( .A(n575), .X(n580) );
  SEN_NR2B_V1DG_1 U668 ( .A(n536), .B(n499), .X(n316) );
  SEN_AN2_1 U669 ( .A1(n498), .A2(n497), .X(n314) );
  SEN_NR3_T_0P5 U670 ( .A1(n519), .A2(n561), .A3(n518), .X(n520) );
  SEN_MUXI2_D_1 U671 ( .D0(n203), .D1(n322), .S(A_qual[22]), .X(n452) );
  SEN_INV_S_0P5 U672 ( .A(n506), .X(n291) );
  SEN_EN2_0P5 U673 ( .A1(n545), .A2(n544), .X(n492) );
  SEN_AN2_S_0P5 U674 ( .A1(n358), .A2(n359), .X(n319) );
  SEN_ND2_S_0P5 U675 ( .A1(n586), .A2(n585), .X(n450) );
  SEN_ND2_S_0P5 U676 ( .A1(n536), .A2(n257), .X(n541) );
  SEN_OR2_DG_1 U677 ( .A1(A_qual[20]), .A2(B_qual[20]), .X(n596) );
  SEN_INV_S_1 U678 ( .A(A_qual[0]), .X(n295) );
  SEN_INV_S_0P5 U679 ( .A(n752), .X(n753) );
  SEN_ND2_S_1 U680 ( .A1(n314), .A2(n524), .X(n502) );
  SEN_NR2_S_0P5 U681 ( .A1(n497), .A2(n461), .X(n465) );
  SEN_INV_S_1 U682 ( .A(n477), .X(n486) );
  SEN_NR3_T_0P5 U683 ( .A1(n562), .A2(n561), .A3(n560), .X(n563) );
  SEN_ND2_S_0P5 U684 ( .A1(n356), .A2(n355), .X(n498) );
  SEN_ND2_0P8 U685 ( .A1(n508), .A2(n509), .X(n357) );
  SEN_ND2_S_0P5 U686 ( .A1(n310), .A2(n856), .X(n565) );
  SEN_NR2_S_0P5 U687 ( .A1(n492), .A2(n495), .X(n302) );
  SEN_INV_S_1 U688 ( .A(n499), .X(n304) );
  SEN_ND2_S_0P5 U689 ( .A1(n364), .A2(n365), .X(n495) );
  SEN_ND2_S_0P5 U690 ( .A1(n545), .A2(n544), .X(n499) );
  SEN_INV_S_0P5 U691 ( .A(n750), .X(n768) );
  SEN_OAOI211_1 U692 ( .A1(n712), .A2(n711), .B(n306), .C(n710), .X(n713) );
  SEN_ND4_S_1 U693 ( .A1(n870), .A2(n869), .A3(n868), .A4(n867), .X(n875) );
  SEN_AOI31_0P5 U694 ( .A1(n650), .A2(n649), .A3(n692), .B(n669), .X(n652) );
  SEN_INV_S_0P5 U695 ( .A(n253), .X(n655) );
  SEN_OAOI211_0P5 U696 ( .A1(n668), .A2(n667), .B(n279), .C(n666), .X(n670) );
  SEN_OAOI211_0P5 U697 ( .A1(n671), .A2(n724), .B(n670), .C(n669), .X(n672) );
  SEN_ND2_S_0P5 U698 ( .A1(n309), .A2(n722), .X(n671) );
  SEN_OAI21_S_0P5 U699 ( .A1(n306), .A2(n710), .B(n714), .X(n699) );
  SEN_OAI21_S_0P5 U700 ( .A1(n700), .A2(n699), .B(n698), .X(n701) );
  SEN_NR2_S_0P5 U701 ( .A1(n725), .A2(n724), .X(n736) );
  SEN_NR3_1 U702 ( .A1(Z[21]), .A2(Z[20]), .A3(Z[19]), .X(n862) );
  SEN_INV_S_0P5 U703 ( .A(n601), .X(n605) );
  SEN_AOI21B_0P5 U704 ( .A1(n823), .A2(n819), .B(n810), .X(n811) );
  SEN_INV_S_0P5 U705 ( .A(n584), .X(n588) );
  SEN_INV_S_0P5 U706 ( .A(n609), .X(n620) );
  SEN_OAI21_S_0P5 U707 ( .A1(n615), .A2(n624), .B(n614), .X(n616) );
  SEN_OAI21_S_0P5 U708 ( .A1(n685), .A2(n684), .B(n705), .X(n686) );
  SEN_AN4B_0P5 U709 ( .B1(n315), .B2(n680), .B3(n722), .A(n724), .X(n687) );
  SEN_AOI21_S_0P5 U710 ( .A1(n683), .A2(n727), .B(n682), .X(n685) );
  SEN_INV_S_0P5 U711 ( .A(n624), .X(n629) );
  SEN_OAI21_S_0P5 U712 ( .A1(n795), .A2(n794), .B(n793), .X(n796) );
  SEN_NR2_S_1 U713 ( .A1(Z[8]), .A2(Z[6]), .X(n873) );
  SEN_NR2_S_1 U714 ( .A1(Z[23]), .A2(Z[22]), .X(n863) );
  SEN_OAI211_0P5 U715 ( .A1(n771), .A2(n792), .B1(n770), .B2(n769), .X(n772)
         );
  SEN_OA21_1 U716 ( .A1(n740), .A2(n697), .B(n305), .X(n306) );
  SEN_OR3B_0P5 U717 ( .B1(n776), .B2(n751), .A(n768), .X(n755) );
  SEN_INV_S_0P5 U718 ( .A(n279), .X(n381) );
  SEN_AOI22_0P5 U719 ( .A1(n815), .A2(n856), .B1(n336), .B2(n814), .X(n816) );
  SEN_AOI22_0P5 U720 ( .A1(n705), .A2(n856), .B1(n336), .B2(n704), .X(n706) );
  SEN_AOI22_0P5 U721 ( .A1(n764), .A2(n856), .B1(n336), .B2(n763), .X(n765) );
  SEN_AOI22_0P5 U722 ( .A1(n676), .A2(n856), .B1(n336), .B2(n675), .X(n677) );
  SEN_AOI22_0P5 U723 ( .A1(n740), .A2(n856), .B1(n336), .B2(n739), .X(n741) );
  SEN_INV_S_1 U724 ( .A(n481), .X(n336) );
  SEN_EN2_0P5 U725 ( .A1(n731), .A2(n732), .X(n729) );
  SEN_NR2_S_0P5 U726 ( .A1(n844), .A2(n800), .X(n801) );
  SEN_NR2_S_0P5 U727 ( .A1(n844), .A2(n776), .X(n777) );
  SEN_NR2_S_0P5 U728 ( .A1(n844), .A2(n658), .X(n659) );
  SEN_NR2_S_0P5 U729 ( .A1(n844), .A2(n639), .X(n640) );
  SEN_NR2_S_1 U730 ( .A1(Z[5]), .A2(Z[3]), .X(n868) );
  SEN_INV_S_0P5 U731 ( .A(n341), .X(n331) );
  SEN_INV_S_0P5 U732 ( .A(n323), .X(n322) );
  SEN_ND2_S_0P5 U733 ( .A1(n479), .A2(n484), .X(n505) );
  SEN_ND2_S_0P5 U734 ( .A1(n618), .A2(n617), .X(n441) );
  SEN_INV_S_0P5 U735 ( .A(INST_qual[1]), .X(n485) );
  SEN_MUXI2_S_0P5 U736 ( .D0(n201), .D1(n321), .S(A_qual[16]), .X(n389) );
  SEN_ND2_S_0P5 U737 ( .A1(n324), .A2(n392), .X(n617) );
  SEN_MUXI2_S_0P5 U738 ( .D0(n203), .D1(n321), .S(A_qual[18]), .X(n392) );
  SEN_ND2_S_0P5 U739 ( .A1(n324), .A2(n446), .X(n594) );
  SEN_MUXI2_S_0P5 U740 ( .D0(n203), .D1(n321), .S(A_qual[20]), .X(n446) );
  SEN_ND2_S_0P5 U741 ( .A1(n325), .A2(n449), .X(n585) );
  SEN_MUXI2_S_0P5 U742 ( .D0(n203), .D1(n321), .S(A_qual[21]), .X(n449) );
  SEN_MUXI2_S_0P5 U743 ( .D0(n474), .D1(n327), .S(B_qual[17]), .X(n386) );
  SEN_ND2_S_0P5 U744 ( .A1(n256), .A2(n475), .X(n483) );
  SEN_MUXI2_S_0P5 U745 ( .D0(n202), .D1(n321), .S(A_qual[19]), .X(n444) );
  SEN_ND2_T_0P5 U746 ( .A1(n254), .A2(n391), .X(n618) );
  SEN_MUXI2_S_0P5 U747 ( .D0(n330), .D1(n328), .S(B_qual[18]), .X(n391) );
  SEN_ND2_S_0P5 U748 ( .A1(n256), .A2(n445), .X(n595) );
  SEN_MUXI2_S_0P5 U749 ( .D0(n330), .D1(n328), .S(B_qual[20]), .X(n445) );
  SEN_ND2_S_0P5 U750 ( .A1(n255), .A2(n448), .X(n586) );
  SEN_MUXI2_S_0P5 U751 ( .D0(n330), .D1(n328), .S(B_qual[21]), .X(n448) );
  SEN_ND2_S_0P5 U752 ( .A1(n255), .A2(n451), .X(n578) );
  SEN_MUXI2_S_0P5 U753 ( .D0(n330), .D1(n328), .S(B_qual[22]), .X(n451) );
  SEN_ND2_S_0P5 U754 ( .A1(n254), .A2(n454), .X(n569) );
  SEN_ND2_S_0P5 U755 ( .A1(n255), .A2(n456), .X(n553) );
  SEN_MUXI2_S_0P5 U756 ( .D0(n330), .D1(n328), .S(B_qual[19]), .X(n443) );
  SEN_OAOI211_0P5 U757 ( .A1(B_qual[15]), .A2(A_qual[15]), .B(n335), .C(n659), 
        .X(n663) );
  SEN_EO2_S_0P5 U758 ( .A1(n215), .A2(n657), .X(n664) );
  SEN_OAOI211_0P5 U759 ( .A1(B_qual[5]), .A2(A_qual[5]), .B(n335), .C(n801), 
        .X(n805) );
  SEN_ND2_S_0P5 U760 ( .A1(n255), .A2(n349), .X(n356) );
  SEN_MUXI2_S_0P5 U761 ( .D0(n331), .D1(n328), .S(B_qual[28]), .X(n349) );
  SEN_OAOI211_0P5 U762 ( .A1(B_qual[11]), .A2(A_qual[11]), .B(n335), .C(n716), 
        .X(n720) );
  SEN_NR2_S_0P5 U763 ( .A1(n426), .A2(INST_qual[3]), .X(n427) );
  SEN_ND2_S_0P5 U764 ( .A1(n255), .A2(n344), .X(n358) );
  SEN_MUXI2_S_0P5 U765 ( .D0(n331), .D1(n328), .S(B_qual[27]), .X(n344) );
  SEN_MUXI2_S_0P5 U766 ( .D0(n202), .D1(n320), .S(A_qual[17]), .X(n387) );
  SEN_OAOI211_0P5 U767 ( .A1(B_qual[1]), .A2(A_qual[1]), .B(n335), .C(n845), 
        .X(n849) );
  SEN_OAOI211_0P5 U768 ( .A1(B_qual[7]), .A2(A_qual[7]), .B(n335), .C(n777), 
        .X(n781) );
  SEN_OAOI211_0P5 U769 ( .A1(B_qual[10]), .A2(A_qual[10]), .B(n335), .C(n730), 
        .X(n734) );
  SEN_ND2_S_0P5 U770 ( .A1(n325), .A2(n361), .X(n544) );
  SEN_MUXI2_S_0P5 U771 ( .D0(n202), .D1(n320), .S(A_qual[26]), .X(n361) );
  SEN_ND2_S_0P5 U772 ( .A1(n324), .A2(n350), .X(n355) );
  SEN_MUXI2_S_0P5 U773 ( .D0(n202), .D1(n320), .S(A_qual[28]), .X(n350) );
  SEN_ND2_S_0P5 U774 ( .A1(n290), .A2(n354), .X(n509) );
  SEN_MUXI2_S_0P5 U775 ( .D0(n203), .D1(n320), .S(A_qual[30]), .X(n354) );
  SEN_INV_S_0P5 U776 ( .A(n466), .X(n470) );
  SEN_MUXI2_S_0P5 U777 ( .D0(n470), .D1(n469), .S(A_qual[31]), .X(n471) );
  SEN_MUXI2_S_0P5 U778 ( .D0(n202), .D1(n320), .S(A_qual[14]), .X(n369) );
  SEN_ND2_S_0P5 U779 ( .A1(n290), .A2(n352), .X(n531) );
  SEN_MUXI2_S_0P5 U780 ( .D0(n203), .D1(n320), .S(A_qual[29]), .X(n352) );
  SEN_ND2_S_0P5 U781 ( .A1(n325), .A2(n363), .X(n365) );
  SEN_MUXI2_S_0P5 U782 ( .D0(n203), .D1(n320), .S(A_qual[25]), .X(n363) );
  SEN_ND2_S_0P5 U783 ( .A1(n325), .A2(n348), .X(n359) );
  SEN_MUXI2_S_0P5 U784 ( .D0(n202), .D1(n320), .S(A_qual[27]), .X(n348) );
  SEN_ND2_S_0P5 U785 ( .A1(n256), .A2(n351), .X(n530) );
  SEN_MUXI2_S_0P5 U786 ( .D0(n331), .D1(n328), .S(B_qual[29]), .X(n351) );
  SEN_ND2_S_0P5 U787 ( .A1(n256), .A2(n353), .X(n508) );
  SEN_MUXI2_S_0P5 U788 ( .D0(n331), .D1(n328), .S(B_qual[30]), .X(n353) );
  SEN_ND2_S_0P5 U789 ( .A1(n254), .A2(n360), .X(n545) );
  SEN_MUXI2_S_0P5 U790 ( .D0(n331), .D1(n328), .S(B_qual[26]), .X(n360) );
  SEN_ND2_S_0P5 U791 ( .A1(n254), .A2(n362), .X(n364) );
  SEN_MUXI2_S_0P5 U792 ( .D0(n331), .D1(n328), .S(B_qual[25]), .X(n362) );
  SEN_OAI21_S_0P5 U793 ( .A1(A_qual[31]), .A2(B_qual[31]), .B(n337), .X(n489)
         );
  SEN_OR3B_0P5 U794 ( .B1(n480), .B2(INST_qual[1]), .A(n484), .X(n481) );
  SEN_OR2_DG_1 U795 ( .A1(B_qual[0]), .A2(A_qual[0]), .X(n855) );
  SEN_OR2_DG_1 U796 ( .A1(A_qual[4]), .A2(B_qual[4]), .X(n814) );
  SEN_OR2_DG_1 U797 ( .A1(A_qual[3]), .A2(B_qual[3]), .X(n822) );
  SEN_OR2_DG_1 U798 ( .A1(A_qual[6]), .A2(B_qual[6]), .X(n787) );
  SEN_OR2_DG_1 U799 ( .A1(A_qual[8]), .A2(B_qual[8]), .X(n763) );
  SEN_OR2_DG_1 U800 ( .A1(A_qual[9]), .A2(B_qual[9]), .X(n739) );
  SEN_OR2_DG_1 U801 ( .A1(A_qual[12]), .A2(B_qual[12]), .X(n704) );
  SEN_OR2_DG_1 U802 ( .A1(A_qual[13]), .A2(B_qual[13]), .X(n691) );
  SEN_OR2_DG_1 U803 ( .A1(A_qual[14]), .A2(B_qual[14]), .X(n675) );
  SEN_OR2_DG_1 U804 ( .A1(A_qual[17]), .A2(B_qual[17]), .X(n628) );
  SEN_OR2_DG_1 U805 ( .A1(A_qual[18]), .A2(B_qual[18]), .X(n619) );
  SEN_OR2_DG_1 U806 ( .A1(A_qual[19]), .A2(B_qual[19]), .X(n604) );
  SEN_INV_S_1 U807 ( .A(n724), .X(n653) );
  SEN_INV_S_1 U808 ( .A(n682), .X(n665) );
  SEN_ND3_S_0P5 U809 ( .A1(n647), .A2(n646), .A3(n311), .X(n650) );
  SEN_NR2_1 U810 ( .A1(n515), .A2(n493), .X(n496) );
  SEN_INV_S_1 U811 ( .A(n505), .X(n339) );
  SEN_INV_S_1 U812 ( .A(n505), .X(n338) );
  SEN_INV_S_1 U813 ( .A(n505), .X(n340) );
  SEN_OAI21_G_1 U814 ( .A1(n687), .A2(n686), .B(n279), .X(n688) );
  SEN_EN2_0P5 U815 ( .A1(n518), .A2(n519), .X(n493) );
  SEN_ND2_S_0P5 U816 ( .A1(n318), .A2(n722), .X(n636) );
  SEN_EN2_0P5 U817 ( .A1(n537), .A2(n538), .X(n491) );
  SEN_AOI211_0P5 U818 ( .A1(n759), .A2(n758), .B1(n757), .B2(n756), .X(n760)
         );
  SEN_OAI21_S_0P5 U819 ( .A1(n749), .A2(n312), .B(n748), .X(n757) );
  SEN_INV_S_1 U820 ( .A(n769), .X(n758) );
  SEN_EN2_0P5 U821 ( .A1(n299), .A2(FLAGS[1]), .X(FLAGS[0]) );
  SEN_EO2_S_0P5 U822 ( .A1(n560), .A2(n562), .X(n310) );
  SEN_INV_S_1 U823 ( .A(n492), .X(n547) );
  SEN_NR2_1 U824 ( .A1(n656), .A2(n655), .X(n657) );
  SEN_ND2_G_1 U825 ( .A1(n527), .A2(n291), .X(n461) );
  SEN_INV_S_1 U826 ( .A(n551), .X(n555) );
  SEN_INV_S_1 U827 ( .A(n592), .X(n597) );
  SEN_INV_S_1 U828 ( .A(n772), .X(n784) );
  SEN_INV_S_1 U829 ( .A(n528), .X(n527) );
  SEN_NR2_1 U830 ( .A1(n797), .A2(n796), .X(n798) );
  SEN_ND2_G_1 U831 ( .A1(n486), .A2(n257), .X(n487) );
  SEN_INV_S_1 U832 ( .A(n567), .X(n571) );
  SEN_OAI21_G_1 U833 ( .A1(n830), .A2(n265), .B(n828), .X(n831) );
  SEN_INV_S_1 U834 ( .A(n827), .X(n830) );
  SEN_OAI21_G_1 U835 ( .A1(n500), .A2(n506), .B(n357), .X(n463) );
  SEN_NR2_1 U836 ( .A1(n498), .A2(n461), .X(n464) );
  SEN_ND3_S_0P5 U837 ( .A1(n799), .A2(n747), .A3(n746), .X(n769) );
  SEN_ND2_G_1 U838 ( .A1(n528), .A2(n500), .X(n501) );
  SEN_ND2_G_1 U839 ( .A1(n319), .A2(n517), .X(n497) );
  SEN_INV_S_1 U840 ( .A(Z[4]), .X(n869) );
  SEN_INV_S_1 U841 ( .A(n561), .X(n333) );
  SEN_INV_S_1 U842 ( .A(n561), .X(n334) );
  SEN_INV_S_1 U843 ( .A(n844), .X(n856) );
  SEN_OAI211_1 U844 ( .A1(n826), .A2(n338), .B1(n825), .B2(n824), .X(Z[3]) );
  SEN_ND3_S_0P5 U845 ( .A1(n821), .A2(n333), .A3(n820), .X(n825) );
  SEN_AOI22_1 U846 ( .A1(n823), .A2(n856), .B1(n336), .B2(n822), .X(n824) );
  SEN_EN2_0P5 U847 ( .A1(n823), .A2(n819), .X(n826) );
  SEN_NR2_S_0P5 U848 ( .A1(n844), .A2(n729), .X(n730) );
  SEN_NR2_1 U849 ( .A1(n844), .A2(n528), .X(n529) );
  SEN_NR2_1 U850 ( .A1(n844), .A2(n506), .X(n507) );
  SEN_EN2_0P5 U851 ( .A1(n553), .A2(n552), .X(n551) );
  SEN_EN2_0P5 U852 ( .A1(n595), .A2(n594), .X(n592) );
  SEN_EN2_0P5 U853 ( .A1(n530), .A2(n531), .X(n528) );
  SEN_EN2_0P5 U854 ( .A1(n603), .A2(n602), .X(n601) );
  SEN_EN2_0P5 U855 ( .A1(n578), .A2(n577), .X(n575) );
  SEN_EN2_0P5 U856 ( .A1(n569), .A2(n568), .X(n567) );
  SEN_EN2_0P5 U857 ( .A1(n586), .A2(n585), .X(n584) );
  SEN_OAI211_1 U858 ( .A1(n791), .A2(n338), .B1(n790), .B2(n789), .X(Z[6]) );
  SEN_AOI22_1 U859 ( .A1(n788), .A2(n856), .B1(n336), .B2(n787), .X(n789) );
  SEN_EO2_S_0P5 U860 ( .A1(n788), .A2(n784), .X(n791) );
  SEN_OAI211_1 U861 ( .A1(n591), .A2(n339), .B1(n590), .B2(n589), .X(Z[21]) );
  SEN_ND3_S_0P5 U862 ( .A1(n586), .A2(n334), .A3(n585), .X(n590) );
  SEN_AOI22_1 U863 ( .A1(n588), .A2(n856), .B1(n336), .B2(n587), .X(n589) );
  SEN_EN2_0P5 U864 ( .A1(n588), .A2(n214), .X(n591) );
  SEN_EN2_0P5 U865 ( .A1(n482), .A2(n483), .X(n477) );
  SEN_OAI211_1 U866 ( .A1(n860), .A2(n339), .B1(n859), .B2(n858), .X(Z[0]) );
  SEN_ND3_S_0P5 U867 ( .A1(n854), .A2(n333), .A3(n853), .X(n859) );
  SEN_AOI22_1 U868 ( .A1(n857), .A2(n856), .B1(n336), .B2(n855), .X(n858) );
  SEN_EN2_0P5 U869 ( .A1(n283), .A2(n857), .X(n860) );
  SEN_OAI211_1 U870 ( .A1(n767), .A2(n338), .B1(n766), .B2(n765), .X(Z[8]) );
  SEN_ND3_S_0P5 U871 ( .A1(n762), .A2(n333), .A3(n761), .X(n766) );
  SEN_EO2_S_0P5 U872 ( .A1(n764), .A2(n760), .X(n767) );
  SEN_OAI211_1 U873 ( .A1(n608), .A2(n339), .B1(n607), .B2(n606), .X(Z[19]) );
  SEN_ND3_S_0P5 U874 ( .A1(n603), .A2(n333), .A3(n602), .X(n607) );
  SEN_AOI22_1 U875 ( .A1(n605), .A2(n856), .B1(n336), .B2(n604), .X(n606) );
  SEN_EO2_S_0P5 U876 ( .A1(n605), .A2(n217), .X(n608) );
  SEN_OAI211_1 U877 ( .A1(n743), .A2(n338), .B1(n742), .B2(n741), .X(Z[9]) );
  SEN_ND3_S_0P5 U878 ( .A1(n738), .A2(n333), .A3(n737), .X(n742) );
  SEN_EO2_S_0P5 U879 ( .A1(n740), .A2(n736), .X(n743) );
  SEN_OAI211_1 U880 ( .A1(n583), .A2(n339), .B1(n582), .B2(n581), .X(Z[22]) );
  SEN_ND3_S_0P5 U881 ( .A1(n578), .A2(n333), .A3(n577), .X(n582) );
  SEN_AOI22_1 U882 ( .A1(n580), .A2(n257), .B1(n336), .B2(n579), .X(n581) );
  SEN_EN2_0P5 U883 ( .A1(n580), .A2(n204), .X(n583) );
  SEN_OAI211_1 U884 ( .A1(n818), .A2(n338), .B1(n817), .B2(n816), .X(Z[4]) );
  SEN_ND3_S_0P5 U885 ( .A1(n813), .A2(n333), .A3(n812), .X(n817) );
  SEN_OAI211_1 U886 ( .A1(n600), .A2(n339), .B1(n599), .B2(n598), .X(Z[20]) );
  SEN_ND3_S_0P5 U887 ( .A1(n595), .A2(n334), .A3(n594), .X(n599) );
  SEN_AOI22_1 U888 ( .A1(n597), .A2(n856), .B1(n336), .B2(n596), .X(n598) );
  SEN_EN2_0P5 U889 ( .A1(n597), .A2(n207), .X(n600) );
  SEN_OAI211_1 U890 ( .A1(n695), .A2(n338), .B1(n694), .B2(n693), .X(Z[13]) );
  SEN_ND3_S_0P5 U891 ( .A1(n690), .A2(n333), .A3(n689), .X(n694) );
  SEN_AOI22_1 U892 ( .A1(n692), .A2(n856), .B1(n336), .B2(n691), .X(n693) );
  SEN_EN2_0P5 U893 ( .A1(n692), .A2(n688), .X(n695) );
  SEN_OAI211_1 U894 ( .A1(n679), .A2(n338), .B1(n678), .B2(n677), .X(Z[14]) );
  SEN_ND3_S_0P5 U895 ( .A1(n674), .A2(n333), .A3(n673), .X(n678) );
  SEN_EO2_S_0P5 U896 ( .A1(n676), .A2(n672), .X(n679) );
  SEN_ND3_S_0P5 U897 ( .A1(n545), .A2(n334), .A3(n544), .X(n549) );
  SEN_AOI22_1 U898 ( .A1(n547), .A2(n257), .B1(n337), .B2(n546), .X(n548) );
  SEN_AO2BB2_1 U899 ( .A1(n299), .A2(n477), .B1(n483), .B2(n482), .X(FLAGS[1])
         );
  SEN_OAI211_1 U900 ( .A1(n558), .A2(n339), .B1(n557), .B2(n556), .X(Z[24]) );
  SEN_ND3_S_0P5 U901 ( .A1(n553), .A2(n333), .A3(n552), .X(n557) );
  SEN_AOI22_1 U902 ( .A1(n555), .A2(n257), .B1(n337), .B2(n554), .X(n556) );
  SEN_EN2_0P5 U903 ( .A1(n555), .A2(n213), .X(n558) );
  SEN_OAI211_1 U904 ( .A1(n632), .A2(n339), .B1(n631), .B2(n630), .X(Z[17]) );
  SEN_ND3_S_0P5 U905 ( .A1(n627), .A2(n333), .A3(n626), .X(n631) );
  SEN_AOI22_1 U906 ( .A1(n629), .A2(n856), .B1(n336), .B2(n628), .X(n630) );
  SEN_EN2_0P5 U907 ( .A1(n629), .A2(n625), .X(n632) );
  SEN_OAI211_1 U908 ( .A1(n708), .A2(n338), .B1(n707), .B2(n706), .X(Z[12]) );
  SEN_ND3_S_0P5 U909 ( .A1(n703), .A2(n333), .A3(n702), .X(n707) );
  SEN_EN2_0P5 U910 ( .A1(n705), .A2(n701), .X(n708) );
  SEN_OAI211_1 U911 ( .A1(n574), .A2(n339), .B1(n573), .B2(n572), .X(Z[23]) );
  SEN_ND3_S_0P5 U912 ( .A1(n569), .A2(n334), .A3(n568), .X(n573) );
  SEN_AOI22_1 U913 ( .A1(n571), .A2(n257), .B1(n337), .B2(n570), .X(n572) );
  SEN_EN2_0P5 U914 ( .A1(n571), .A2(n212), .X(n574) );
  SEN_OAI211_1 U915 ( .A1(n623), .A2(n339), .B1(n622), .B2(n621), .X(Z[18]) );
  SEN_ND3_S_0P5 U916 ( .A1(n618), .A2(n333), .A3(n617), .X(n622) );
  SEN_AOI22_1 U917 ( .A1(n620), .A2(n856), .B1(n336), .B2(n619), .X(n621) );
  SEN_EN2_0P5 U918 ( .A1(n620), .A2(n616), .X(n623) );
  SEN_ND2_G_1 U919 ( .A1(n530), .A2(n531), .X(n500) );
  SEN_ND2_G_1 U920 ( .A1(n553), .A2(n552), .X(n460) );
  SEN_INV_S_1 U921 ( .A(n356), .X(n518) );
  SEN_INV_S_1 U922 ( .A(n358), .X(n537) );
  SEN_INV_S_1 U923 ( .A(n364), .X(n560) );
  SEN_INV_S_1 U924 ( .A(n355), .X(n519) );
  SEN_INV_S_1 U925 ( .A(n359), .X(n538) );
  SEN_INV_S_1 U926 ( .A(n365), .X(n562) );
  SEN_NR3_G_1 U927 ( .A1(Z[2]), .A2(Z[1]), .A3(Z[0]), .X(n870) );
  SEN_NR2_S_1 U928 ( .A1(Z[17]), .A2(Z[16]), .X(n864) );
  SEN_NR3_1 U929 ( .A1(Z[14]), .A2(Z[13]), .A3(Z[15]), .X(n866) );
  SEN_ND3_S_0P5 U930 ( .A1(n334), .A2(n483), .A3(n482), .X(n488) );
  SEN_INV_S_1 U931 ( .A(n481), .X(n335) );
  SEN_NR2_S_1 U932 ( .A1(Z[12]), .A2(Z[11]), .X(n871) );
  SEN_NR2_S_1 U933 ( .A1(Z[10]), .A2(Z[9]), .X(n867) );
  SEN_INV_S_1 U934 ( .A(Z[7]), .X(n872) );
  SEN_INV_S_1 U935 ( .A(n481), .X(n337) );
  SEN_OAI211_1 U936 ( .A1(n340), .A2(n782), .B1(n781), .B2(n780), .X(Z[7]) );
  SEN_ND3_S_0P5 U937 ( .A1(n334), .A2(n779), .A3(n778), .X(n780) );
  SEN_ND2_G_1 U938 ( .A1(n324), .A2(n471), .X(n482) );
  SEN_MUXI2_S_1 U939 ( .D0(n331), .D1(n328), .S(B_qual[31]), .X(n475) );
  SEN_ND2_G_1 U940 ( .A1(n290), .A2(n452), .X(n577) );
  SEN_ND2_G_1 U941 ( .A1(n324), .A2(n455), .X(n568) );
  SEN_MUXI2_S_1 U942 ( .D0(n202), .D1(n322), .S(A_qual[23]), .X(n455) );
  SEN_MUXI2_S_1 U943 ( .D0(n202), .D1(n322), .S(A_qual[24]), .X(n459) );
  SEN_OAI211_1 U944 ( .A1(n340), .A2(n850), .B1(n849), .B2(n848), .X(Z[1]) );
  SEN_ND3_S_0P5 U945 ( .A1(n334), .A2(n847), .A3(n846), .X(n848) );
  SEN_EN2_0P5 U946 ( .A1(n842), .A2(n841), .X(n850) );
  SEN_OAI211_1 U947 ( .A1(n664), .A2(n338), .B1(n663), .B2(n662), .X(Z[15]) );
  SEN_ND3_S_0P5 U948 ( .A1(n334), .A2(n661), .A3(n660), .X(n662) );
  SEN_OAI211_1 U949 ( .A1(n340), .A2(n735), .B1(n734), .B2(n733), .X(Z[10]) );
  SEN_ND3_S_0P5 U950 ( .A1(n334), .A2(n732), .A3(n731), .X(n733) );
  SEN_OAOI211_G_1 U951 ( .A1(B_qual[25]), .A2(A_qual[25]), .B(n335), .C(n563), 
        .X(n564) );
  SEN_OAI211_1 U952 ( .A1(n645), .A2(n338), .B1(n644), .B2(n643), .X(Z[16]) );
  SEN_ND3_S_0P5 U953 ( .A1(n334), .A2(n642), .A3(n641), .X(n643) );
  SEN_OAOI211_G_1 U954 ( .A1(B_qual[16]), .A2(A_qual[16]), .B(n335), .C(n640), 
        .X(n644) );
  SEN_EO2_S_0P5 U955 ( .A1(n638), .A2(n637), .X(n645) );
  SEN_OAI211_1 U956 ( .A1(n721), .A2(n338), .B1(n720), .B2(n719), .X(Z[11]) );
  SEN_ND3_S_0P5 U957 ( .A1(n334), .A2(n718), .A3(n717), .X(n719) );
  SEN_EO2_S_0P5 U958 ( .A1(n714), .A2(n713), .X(n721) );
  SEN_OAI211_1 U959 ( .A1(n839), .A2(n338), .B1(n838), .B2(n837), .X(Z[2]) );
  SEN_ND3_S_0P5 U960 ( .A1(n334), .A2(n836), .A3(n835), .X(n837) );
  SEN_OAOI211_G_1 U961 ( .A1(B_qual[2]), .A2(A_qual[2]), .B(n335), .C(n834), 
        .X(n838) );
  SEN_EN2_0P5 U962 ( .A1(n832), .A2(n831), .X(n839) );
  SEN_OAOI211_G_1 U963 ( .A1(B_qual[27]), .A2(A_qual[27]), .B(n335), .C(n539), 
        .X(n540) );
  SEN_OAI211_1 U964 ( .A1(n806), .A2(n338), .B1(n805), .B2(n804), .X(Z[5]) );
  SEN_ND3_S_0P5 U965 ( .A1(n334), .A2(n803), .A3(n802), .X(n804) );
  SEN_EO2_S_0P5 U966 ( .A1(n799), .A2(n798), .X(n806) );
  SEN_ND3_S_0P5 U967 ( .A1(n334), .A2(n531), .A3(n530), .X(n532) );
  SEN_OAOI211_G_1 U968 ( .A1(B_qual[29]), .A2(A_qual[29]), .B(n335), .C(n529), 
        .X(n533) );
  SEN_ND3_S_0P5 U969 ( .A1(n334), .A2(n509), .A3(n508), .X(n510) );
  SEN_OAOI211_G_1 U970 ( .A1(B_qual[30]), .A2(A_qual[30]), .B(n335), .C(n507), 
        .X(n511) );
  SEN_OAOI211_G_1 U971 ( .A1(B_qual[28]), .A2(A_qual[28]), .B(n335), .C(n520), 
        .X(n521) );
  SEN_ND2_G_1 U972 ( .A1(n517), .A2(n257), .X(n522) );
  SEN_MUXI2_S_1 U973 ( .D0(n331), .D1(n328), .S(B_qual[23]), .X(n454) );
  SEN_MUXI2_S_1 U974 ( .D0(n331), .D1(n328), .S(B_qual[24]), .X(n456) );
  SEN_OR2_1 U975 ( .A1(A_qual[21]), .A2(B_qual[21]), .X(n587) );
  SEN_OR2_1 U976 ( .A1(A_qual[22]), .A2(B_qual[22]), .X(n579) );
  SEN_OR2_1 U977 ( .A1(A_qual[23]), .A2(B_qual[23]), .X(n570) );
  SEN_OR2_1 U978 ( .A1(A_qual[24]), .A2(B_qual[24]), .X(n554) );
  SEN_OR2_1 U979 ( .A1(A_qual[26]), .A2(B_qual[26]), .X(n546) );
  SEN_TIE0_1 U980 ( .X(\*Logic0* ) );
  SEN_AOI311_1 U981 ( .A1(n313), .A2(n722), .A3(n653), .B1(n652), .B2(n651), 
        .X(n656) );
  SEN_OAI31_0P5 U982 ( .A1(n307), .A2(n833), .A3(n809), .B(n808), .X(n819) );
  SEN_NR2_S_0P5 U983 ( .A1(n844), .A2(n715), .X(n716) );
  SEN_ND2_S_0P5 U984 ( .A1(n468), .A2(n467), .X(n469) );
  SEN_EN2_0P5 U985 ( .A1(n775), .A2(n774), .X(n782) );
  SEN_EO2_S_0P5 U986 ( .A1(n815), .A2(n811), .X(n818) );
  SEN_INV_S_0P5 U987 ( .A(n852), .X(n857) );
  SEN_OAI21_S_0P5 U988 ( .A1(n852), .A2(n851), .B(n840), .X(n841) );
  SEN_OAI21_S_0P5 U989 ( .A1(n305), .A2(n710), .B(n714), .X(n682) );
  SEN_NR2_1 U990 ( .A1(n684), .A2(n710), .X(n680) );
  SEN_NR3B_1 U991 ( .A(INST_qual[2]), .B1(A_qual[31]), .B2(INST_qual[0]), .X(
        n426) );
  SEN_ND2_S_0P5 U992 ( .A1(n754), .A2(n753), .X(n792) );
  SEN_NR2_S_0P5 U993 ( .A1(n844), .A2(n843), .X(n845) );
  SEN_ND2_S_0P5 U994 ( .A1(n308), .A2(n610), .X(n612) );
  SEN_AOI21_S_0P5 U995 ( .A1(n633), .A2(n253), .B(n658), .X(n635) );
  SEN_OAI21_S_0P5 U996 ( .A1(n665), .A2(n684), .B(n705), .X(n668) );
  SEN_ND2_S_0P5 U997 ( .A1(n315), .A2(n281), .X(n712) );
  SEN_AN3B_0P5 U998 ( .B1(n281), .B2(n317), .A(n711), .X(n700) );
  SEN_ND3_S_0P5 U999 ( .A1(n786), .A2(n333), .A3(n785), .X(n790) );
  SEN_AO21_2 U1000 ( .A1(INST_qual[3]), .A2(INST_qual[2]), .B(n479), .X(n341)
         );
endmodule

