
module ShiftLR ( Z, X, S, LEFT, LOG );
  output [31:0] Z;
  input [31:0] X;
  input [4:0] S;
  input LEFT, LOG;
  wire   n2, n3, n4, n5, n6, n7, n8, n10, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n89, n90, n92, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355;

  SEN_OAI222_1 U289 ( .A1(n38), .A2(n261), .B1(n150), .B2(n281), .C1(n36), 
        .C2(n123), .X(n131) );
  SEN_EO2_DG_4 U290 ( .A1(S[2]), .A2(n256), .X(n123) );
  SEN_NR2B_V1DG_2 U291 ( .A(n342), .B(n294), .X(n256) );
  SEN_BUF_S_1 U292 ( .A(n104), .X(n281) );
  SEN_INV_2 U293 ( .A(n137), .X(n78) );
  SEN_BUF_S_1 U294 ( .A(n99), .X(n275) );
  SEN_ND2_0P5 U295 ( .A1(n349), .A2(n167), .X(n333) );
  SEN_NR3_G_1 U296 ( .A1(n268), .A2(n269), .A3(n152), .X(n190) );
  SEN_BUF_S_1 U297 ( .A(n104), .X(n280) );
  SEN_INV_S_1 U298 ( .A(n207), .X(n23) );
  SEN_OAI211_1 U299 ( .A1(n66), .A2(n158), .B1(n39), .B2(n172), .X(n151) );
  SEN_AOI22_1 U300 ( .A1(n160), .A2(n344), .B1(n173), .B2(n37), .X(n172) );
  SEN_AO222_1 U301 ( .A1(n115), .A2(n81), .B1(n50), .B2(n83), .C1(n200), .C2(
        n84), .X(n321) );
  SEN_AOI221_1 U302 ( .A1(n115), .A2(n79), .B1(n170), .B2(n81), .C(n226), .X(
        n213) );
  SEN_AOI221_1 U303 ( .A1(n24), .A2(n79), .B1(n164), .B2(n81), .C(n223), .X(
        n209) );
  SEN_AOI221_1 U304 ( .A1(n17), .A2(n79), .B1(n178), .B2(n81), .C(n215), .X(
        n201) );
  SEN_OR3_1 U305 ( .A1(n285), .A2(n286), .A3(n259), .X(n167) );
  SEN_INV_S_1 U306 ( .A(n148), .X(n34) );
  SEN_INV_S_1 U307 ( .A(n279), .X(n81) );
  SEN_BUF_S_1 U308 ( .A(n104), .X(n279) );
  SEN_INV_2 U309 ( .A(n123), .X(n84) );
  SEN_INV_S_1 U310 ( .A(n108), .X(n83) );
  SEN_AOI222_1 U311 ( .A1(n355), .A2(n179), .B1(n350), .B2(n183), .C1(n347), 
        .C2(n22), .X(n184) );
  SEN_ND3_1 U312 ( .A1(n266), .A2(n267), .A3(n149), .X(Z[29]) );
  SEN_AN3_1 U313 ( .A1(n318), .A2(n319), .A3(n320), .X(n149) );
  SEN_OAI221_1 U314 ( .A1(n116), .A2(n317), .B1(n188), .B2(n280), .C(n237), 
        .X(n94) );
  SEN_AN2_S_1 U315 ( .A1(n79), .A2(n258), .X(n257) );
  SEN_INV_S_0P5 U316 ( .A(n257), .X(n352) );
  SEN_INV_S_0P5 U317 ( .A(n257), .X(n351) );
  SEN_AN3_0P5 U318 ( .A1(n130), .A2(n212), .A3(n86), .X(n258) );
  SEN_OAI221_1 U319 ( .A1(n113), .A2(n317), .B1(n190), .B2(n280), .C(n211), 
        .X(n195) );
  SEN_INV_2 U320 ( .A(n238), .X(n355) );
  SEN_INV_1 U321 ( .A(n152), .X(n39) );
  SEN_INV_S_1 U322 ( .A(n338), .X(n349) );
  SEN_AO22_1 U323 ( .A1(n79), .A2(n28), .B1(n81), .B2(n133), .X(n259) );
  SEN_INV_1 U324 ( .A(n216), .X(n32) );
  SEN_INV_S_1 U325 ( .A(n195), .X(n284) );
  SEN_ND2_G_1 U326 ( .A1(n212), .A2(n342), .X(n137) );
  SEN_AOI222_1 U327 ( .A1(n133), .A2(n83), .B1(n134), .B2(n81), .C1(n135), 
        .C2(n84), .X(n132) );
  SEN_OA2BB2_0P5 U328 ( .A1(n130), .A2(n131), .B1(n130), .B2(n132), .X(n129)
         );
  SEN_AOI221_1 U329 ( .A1(n345), .A2(X[21]), .B1(n337), .B2(X[5]), .C(n32), 
        .X(n103) );
  SEN_INV_2 U330 ( .A(n331), .X(n337) );
  SEN_OA2BB2_DG_1 U331 ( .A1(n83), .A2(n24), .B1(n106), .B2(n103), .X(n235) );
  SEN_AN2_DG_1 U332 ( .A1(n197), .A2(n130), .X(n340) );
  SEN_ND2_G_1 U333 ( .A1(n173), .A2(n123), .X(n261) );
  SEN_INV_S_1 U334 ( .A(n80), .X(n260) );
  SEN_OAI22_S_0P5 U335 ( .A1(n261), .A2(n193), .B1(n106), .B2(n175), .X(n215)
         );
  SEN_AO2BB2_0P5 U336 ( .A1(n106), .A2(n166), .B1(n83), .B2(n164), .X(n185) );
  SEN_ND2_G_1 U337 ( .A1(n84), .A2(n82), .X(n106) );
  SEN_ND2_G_0P65 U338 ( .A1(n173), .A2(n123), .X(n108) );
  SEN_OAI211_0P5 U339 ( .A1(n64), .A2(n158), .B1(n39), .B2(n159), .X(n135) );
  SEN_ND2_T_0P5 U340 ( .A1(n78), .A2(n82), .X(n158) );
  SEN_AOI221_1 U341 ( .A1(n346), .A2(X[27]), .B1(n337), .B2(X[11]), .C(n32), 
        .X(n175) );
  SEN_ND2_G_1 U342 ( .A1(n345), .A2(X[22]), .X(n262) );
  SEN_ND2_G_1 U343 ( .A1(n336), .A2(X[6]), .X(n263) );
  SEN_AN3_1 U344 ( .A1(n262), .A2(n263), .A3(n297), .X(n203) );
  SEN_INV_2 U345 ( .A(n331), .X(n336) );
  SEN_AN2_S_1 U346 ( .A1(n346), .A2(X[19]), .X(n264) );
  SEN_AN2_S_0P5 U347 ( .A1(n337), .A2(X[3]), .X(n265) );
  SEN_NR3_0P8 U348 ( .A1(n264), .A2(n265), .A3(n32), .X(n120) );
  SEN_INV_1 U349 ( .A(n341), .X(n346) );
  SEN_OA22_DG_1 U350 ( .A1(n106), .A2(n120), .B1(n261), .B2(n229), .X(n236) );
  SEN_OR2_1 U351 ( .A1(n148), .A2(n354), .X(n266) );
  SEN_OR2_1 U352 ( .A1(n44), .A2(n351), .X(n267) );
  SEN_NR3_T_1 U353 ( .A1(n300), .A2(n301), .A3(n302), .X(n148) );
  SEN_INV_S_1 U354 ( .A(n340), .X(n354) );
  SEN_AN2_S_0P5 U355 ( .A1(X[0]), .A2(n78), .X(n268) );
  SEN_AN2_S_0P5 U356 ( .A1(n337), .A2(X[16]), .X(n269) );
  SEN_NR3_0P8 U357 ( .A1(LOG), .A2(n342), .A3(n40), .X(n152) );
  SEN_AN2_S_0P5 U358 ( .A1(n316), .A2(n117), .X(n270) );
  SEN_AN2_S_0P5 U359 ( .A1(n349), .A2(n321), .X(n271) );
  SEN_AN2_S_1 U360 ( .A1(n347), .A2(n110), .X(n272) );
  SEN_NR3_T_2 U361 ( .A1(n270), .A2(n271), .A3(n272), .X(n124) );
  SEN_OAI222_0P75 U362 ( .A1(n107), .A2(n280), .B1(n101), .B2(n261), .C1(n147), 
        .C2(n123), .X(n117) );
  SEN_OAI222_1 U363 ( .A1(n125), .A2(n280), .B1(n126), .B2(n261), .C1(n127), 
        .C2(n123), .X(n110) );
  SEN_OAI221_0P5 U364 ( .A1(n41), .A2(n354), .B1(n71), .B2(n351), .C(n124), 
        .X(Z[3]) );
  SEN_AN2_S_0P5 U365 ( .A1(n346), .A2(X[13]), .X(n273) );
  SEN_AN2_S_0P5 U366 ( .A1(n246), .A2(X[29]), .X(n274) );
  SEN_NR2_1 U367 ( .A1(n273), .A2(n274), .X(n109) );
  SEN_NR2_T_0P5 U368 ( .A1(n212), .A2(n342), .X(n246) );
  SEN_OA222_1 U369 ( .A1(n69), .A2(n247), .B1(n53), .B2(n248), .C1(n109), .C2(
        n173), .X(n147) );
  SEN_EO2_5 U370 ( .A1(n254), .A2(S[4]), .X(n212) );
  SEN_OAI21_4 U371 ( .A1(S[3]), .A2(n253), .B(n342), .X(n254) );
  SEN_NR2_S_0P5 U372 ( .A1(n193), .A2(n317), .X(n276) );
  SEN_NR2_S_0P5 U373 ( .A1(n155), .A2(n280), .X(n277) );
  SEN_INV_S_1 U374 ( .A(n194), .X(n278) );
  SEN_OR3_1 U375 ( .A1(n276), .A2(n277), .A3(n278), .X(n183) );
  SEN_OA2BB2_0P5 U376 ( .A1(n80), .A2(n178), .B1(n261), .B2(n175), .X(n194) );
  SEN_OA22_1 U377 ( .A1(n261), .A2(n120), .B1(n106), .B2(n193), .X(n230) );
  SEN_ND2_S_0P5 U378 ( .A1(n123), .A2(n82), .X(n104) );
  SEN_OR2_DG_1 U379 ( .A1(n121), .A2(n106), .X(n282) );
  SEN_OR2_DG_1 U380 ( .A1(n122), .A2(n84), .X(n283) );
  SEN_ND3_1 U381 ( .A1(n282), .A2(n283), .A3(n249), .X(n146) );
  SEN_NR2_S_0P5 U382 ( .A1(n181), .A2(n261), .X(n285) );
  SEN_NR2_S_0P5 U383 ( .A1(n161), .A2(n260), .X(n286) );
  SEN_AOI221_1 U384 ( .A1(X[2]), .A2(n78), .B1(X[18]), .B2(n74), .C(n152), .X(
        n161) );
  SEN_OAI221_0P5 U385 ( .A1(n125), .A2(n317), .B1(n181), .B2(n281), .C(n218), 
        .X(n208) );
  SEN_OAI221_0P5 U386 ( .A1(n126), .A2(n317), .B1(n203), .B2(n280), .C(n239), 
        .X(n92) );
  SEN_OAI221_0P5 U387 ( .A1(n101), .A2(n317), .B1(n103), .B2(n280), .C(n105), 
        .X(n95) );
  SEN_OAI221_0P5 U388 ( .A1(n229), .A2(n317), .B1(n175), .B2(n280), .C(n230), 
        .X(n221) );
  SEN_OAI221_0P5 U389 ( .A1(n112), .A2(n317), .B1(n113), .B2(n280), .C(n114), 
        .X(n97) );
  SEN_OAI222_0P5 U390 ( .A1(n120), .A2(n281), .B1(n121), .B2(n261), .C1(n122), 
        .C2(n123), .X(n99) );
  SEN_OAI221_1 U391 ( .A1(n109), .A2(n317), .B1(n207), .B2(n280), .C(n235), 
        .X(n227) );
  SEN_NR2_S_0P5 U392 ( .A1(n73), .A2(n40), .X(n287) );
  SEN_NR2_S_0P5 U393 ( .A1(n136), .A2(n59), .X(n288) );
  SEN_OR3_2 U394 ( .A1(n287), .A2(n288), .A3(n32), .X(n178) );
  SEN_INV_S_2 U395 ( .A(n345), .X(n73) );
  SEN_INV_1 U396 ( .A(X[31]), .X(n40) );
  SEN_ND2_G_1 U397 ( .A1(n75), .A2(n342), .X(n136) );
  SEN_ND2_G_1 U398 ( .A1(n152), .A2(n75), .X(n216) );
  SEN_AOI22_0P75 U399 ( .A1(n160), .A2(X[23]), .B1(n173), .B2(n178), .X(n177)
         );
  SEN_ND2_G_1 U400 ( .A1(n346), .A2(X[18]), .X(n289) );
  SEN_ND2_S_0P5 U401 ( .A1(n336), .A2(X[2]), .X(n290) );
  SEN_INV_S_0P5 U402 ( .A(n32), .X(n291) );
  SEN_AN3_1 U403 ( .A1(n289), .A2(n290), .A3(n291), .X(n125) );
  SEN_OA22_DG_1 U404 ( .A1(n106), .A2(n203), .B1(n261), .B2(n125), .X(n233) );
  SEN_ND2_S_0P5 U405 ( .A1(n346), .A2(X[25]), .X(n292) );
  SEN_ND2_S_0P5 U406 ( .A1(n337), .A2(X[9]), .X(n293) );
  SEN_AN3_1 U407 ( .A1(n292), .A2(n293), .A3(n291), .X(n207) );
  SEN_OAI22_0P5 U408 ( .A1(n261), .A2(n103), .B1(n106), .B2(n207), .X(n223) );
  SEN_BUF_2 U409 ( .A(n355), .X(n316) );
  SEN_ND2_0P5 U410 ( .A1(n84), .A2(n173), .X(n102) );
  SEN_ND2_0P5 U411 ( .A1(n84), .A2(n173), .X(n317) );
  SEN_NR2_S_0P5 U412 ( .A1(S[1]), .A2(S[0]), .X(n294) );
  SEN_ND2_S_0P5 U413 ( .A1(n345), .A2(X[20]), .X(n295) );
  SEN_ND2_S_0P5 U414 ( .A1(n336), .A2(X[4]), .X(n296) );
  SEN_INV_S_0P5 U415 ( .A(n32), .X(n297) );
  SEN_AN3_1 U416 ( .A1(n295), .A2(n296), .A3(n297), .X(n113) );
  SEN_OAI22_S_0P5 U417 ( .A1(n261), .A2(n113), .B1(n106), .B2(n188), .X(n226)
         );
  SEN_OA2BB2_DG_1 U418 ( .A1(n83), .A2(n115), .B1(n106), .B2(n113), .X(n237)
         );
  SEN_NR2_G_0P5 U419 ( .A1(n175), .A2(n317), .X(n326) );
  SEN_OA2BB2_0P5 U420 ( .A1(n160), .A2(X[25]), .B1(n82), .B2(n166), .X(n165)
         );
  SEN_ND2_2 U421 ( .A1(n324), .A2(n325), .X(n173) );
  SEN_ND2_0P65 U422 ( .A1(n349), .A2(n33), .X(n309) );
  SEN_ND2_G_1 U423 ( .A1(n348), .A2(n33), .X(n334) );
  SEN_OAI221_1 U424 ( .A1(n168), .A2(n354), .B1(n48), .B2(n351), .C(n169), .X(
        Z[25]) );
  SEN_ND2_S_0P5 U425 ( .A1(X[1]), .A2(n78), .X(n303) );
  SEN_ND2_S_0P5 U426 ( .A1(n74), .A2(X[17]), .X(n304) );
  SEN_AN3_1 U427 ( .A1(n303), .A2(n304), .A3(n39), .X(n166) );
  SEN_NR2_T_2 U428 ( .A1(S[1]), .A2(S[0]), .X(n255) );
  SEN_INV_1 U429 ( .A(n102), .X(n79) );
  SEN_INV_2 U430 ( .A(n136), .X(n74) );
  SEN_AN3_S_1 U431 ( .A1(n305), .A2(n306), .A3(n307), .X(n153) );
  SEN_INV_4 U432 ( .A(n212), .X(n75) );
  SEN_INV_S_0P5 U433 ( .A(n252), .X(n322) );
  SEN_AN3_1 U434 ( .A1(n308), .A2(n309), .A3(n310), .X(n157) );
  SEN_AN3_1 U435 ( .A1(n332), .A2(n333), .A3(n334), .X(n169) );
  SEN_ND2_S_0P5 U436 ( .A1(n346), .A2(n344), .X(n298) );
  SEN_ND2_S_0P5 U437 ( .A1(n336), .A2(X[8]), .X(n299) );
  SEN_AN3_1 U438 ( .A1(n298), .A2(n299), .A3(n291), .X(n188) );
  SEN_OA2BB2_0P5 U439 ( .A1(n80), .A2(n170), .B1(n108), .B2(n188), .X(n211) );
  SEN_AN2_S_0P5 U440 ( .A1(n164), .A2(n79), .X(n300) );
  SEN_AN2_S_1 U441 ( .A1(n144), .A2(n80), .X(n301) );
  SEN_AN2_DG_1 U442 ( .A1(n142), .A2(n123), .X(n302) );
  SEN_OAI221_0P5 U443 ( .A1(n69), .A2(n137), .B1(n331), .B2(n53), .C(n39), .X(
        n144) );
  SEN_INV_1 U444 ( .A(n106), .X(n80) );
  SEN_INV_2 U445 ( .A(n341), .X(n345) );
  SEN_INV_1 U446 ( .A(n153), .X(n33) );
  SEN_OAI221_1 U447 ( .A1(n153), .A2(n354), .B1(n45), .B2(n351), .C(n154), .X(
        Z[28]) );
  SEN_ND2_S_0P5 U448 ( .A1(n151), .A2(n123), .X(n307) );
  SEN_AOI221_0P5 U449 ( .A1(X[3]), .A2(n78), .B1(n337), .B2(X[19]), .C(n152), 
        .X(n155) );
  SEN_ND2_S_0P5 U450 ( .A1(n170), .A2(n79), .X(n305) );
  SEN_ND2_S_0P5 U451 ( .A1(n171), .A2(n80), .X(n306) );
  SEN_OAI221_0P5 U452 ( .A1(n73), .A2(n45), .B1(n331), .B2(n62), .C(n216), .X(
        n170) );
  SEN_NR2B_V1DG_1 U453 ( .A(n246), .B(n102), .X(n244) );
  SEN_INV_S_1 U454 ( .A(n339), .X(n347) );
  SEN_INV_S_0P5 U455 ( .A(S[3]), .X(n323) );
  SEN_ND2B_V1_3 U456 ( .A(S[2]), .B(n255), .X(n253) );
  SEN_ND2_S_0P5 U457 ( .A1(n316), .A2(n34), .X(n308) );
  SEN_ND2_S_0P5 U458 ( .A1(n347), .A2(n335), .X(n310) );
  SEN_ND2_S_0P5 U459 ( .A1(n355), .A2(n208), .X(n311) );
  SEN_ND2_S_0P5 U460 ( .A1(n350), .A2(n20), .X(n312) );
  SEN_ND2_S_0P5 U461 ( .A1(n347), .A2(n15), .X(n313) );
  SEN_AN3_S_1 U462 ( .A1(n311), .A2(n312), .A3(n313), .X(n214) );
  SEN_ND2_S_0P5 U463 ( .A1(n345), .A2(X[23]), .X(n314) );
  SEN_ND2_S_0P5 U464 ( .A1(n336), .A2(X[7]), .X(n315) );
  SEN_AN3_1 U465 ( .A1(n314), .A2(n315), .A3(n297), .X(n193) );
  SEN_OAI221_1 U466 ( .A1(n121), .A2(n317), .B1(n193), .B2(n280), .C(n236), 
        .X(n90) );
  SEN_OA2BB2_DG_1 U467 ( .A1(n140), .A2(n130), .B1(n141), .B2(n130), .X(n128)
         );
  SEN_NR2_S_0P5 U468 ( .A1(n35), .A2(n84), .X(n328) );
  SEN_ND2_S_0P5 U469 ( .A1(n252), .A2(n323), .X(n324) );
  SEN_AOI222_1 U470 ( .A1(n355), .A2(n167), .B1(n350), .B2(n22), .C1(n347), 
        .C2(n162), .X(n174) );
  SEN_ND3_S_1 U471 ( .A1(n329), .A2(n330), .A3(n204), .X(n186) );
  SEN_ND2_S_0P5 U472 ( .A1(n246), .A2(n173), .X(n248) );
  SEN_ND2_S_0P5 U473 ( .A1(n345), .A2(n173), .X(n247) );
  SEN_OAI222_0P5 U474 ( .A1(n70), .A2(n247), .B1(n54), .B2(n248), .C1(n116), 
        .C2(n173), .X(n200) );
  SEN_ND2_S_0P5 U475 ( .A1(n355), .A2(n140), .X(n318) );
  SEN_ND2_G_1 U476 ( .A1(n348), .A2(n131), .X(n320) );
  SEN_OA222_0P5 U477 ( .A1(n67), .A2(n247), .B1(n51), .B2(n248), .C1(n229), 
        .C2(n173), .X(n122) );
  SEN_INV_S_0P5 U478 ( .A(n173), .X(n82) );
  SEN_AOI221_0P5 U479 ( .A1(X[30]), .A2(n346), .B1(X[14]), .B2(n337), .C(n32), 
        .X(n181) );
  SEN_ND2_S_0P5 U480 ( .A1(n316), .A2(n162), .X(n332) );
  SEN_ND2_S_0P5 U481 ( .A1(n349), .A2(n335), .X(n319) );
  SEN_ND2_2 U482 ( .A1(n322), .A2(S[3]), .X(n325) );
  SEN_OA222_0P5 U483 ( .A1(n68), .A2(n247), .B1(n52), .B2(n248), .C1(n232), 
        .C2(n173), .X(n127) );
  SEN_INV_S_1 U484 ( .A(n340), .X(n353) );
  SEN_OA22_DG_1 U485 ( .A1(n106), .A2(n107), .B1(n108), .B2(n109), .X(n105) );
  SEN_OA22_DG_1 U486 ( .A1(n106), .A2(n125), .B1(n108), .B2(n232), .X(n239) );
  SEN_AOI22_0P5 U487 ( .A1(n83), .A2(n170), .B1(n80), .B2(n37), .X(n189) );
  SEN_AOI222_0P5 U488 ( .A1(n115), .A2(n81), .B1(n50), .B2(n83), .C1(n200), 
        .C2(n84), .X(n118) );
  SEN_NR2_G_1 U489 ( .A1(n257), .A2(n343), .X(n197) );
  SEN_AOI222_1 U490 ( .A1(n316), .A2(n275), .B1(n349), .B2(n110), .C1(n348), 
        .C2(n97), .X(n111) );
  SEN_AOI22_0P5 U491 ( .A1(n83), .A2(n28), .B1(n80), .B2(n31), .X(n204) );
  SEN_OR3_1 U492 ( .A1(n326), .A2(n327), .A3(n328), .X(n162) );
  SEN_OAI22_S_0P5 U493 ( .A1(n147), .A2(n84), .B1(n101), .B2(n106), .X(n245)
         );
  SEN_AOI221_0P5 U494 ( .A1(n346), .A2(X[26]), .B1(n336), .B2(X[10]), .C(n32), 
        .X(n219) );
  SEN_AOI22_0P5 U495 ( .A1(n343), .A2(n196), .B1(n257), .B2(X[0]), .X(n241) );
  SEN_OAI221_0P5 U496 ( .A1(n240), .A2(n353), .B1(n43), .B2(n238), .C(n241), 
        .X(Z[0]) );
  SEN_INV_1 U497 ( .A(n176), .X(n35) );
  SEN_EO2_S_0P5 U498 ( .A1(n251), .A2(S[1]), .X(n130) );
  SEN_AO221_0P5 U499 ( .A1(n196), .A2(n197), .B1(n198), .B2(n350), .C(n199), 
        .X(Z[1]) );
  SEN_AO22_DG_1 U500 ( .A1(n348), .A2(n321), .B1(n257), .B2(X[1]), .X(n199) );
  SEN_NR2_S_0P5 U501 ( .A1(n155), .A2(n106), .X(n327) );
  SEN_INV_1 U502 ( .A(n162), .X(n29) );
  SEN_AOI222_1 U503 ( .A1(n355), .A2(n183), .B1(n350), .B2(n186), .C1(n347), 
        .C2(n179), .X(n187) );
  SEN_AOI22_0P5 U504 ( .A1(n83), .A2(n23), .B1(n80), .B2(n164), .X(n206) );
  SEN_INV_S_0P5 U505 ( .A(n130), .X(n85) );
  SEN_INV_S_0P5 U506 ( .A(n186), .X(n5) );
  SEN_AOI222_0P5 U507 ( .A1(n31), .A2(n79), .B1(n133), .B2(n80), .C1(n135), 
        .C2(n123), .X(n138) );
  SEN_INV_S_0P5 U508 ( .A(n120), .X(n17) );
  SEN_AOI222_0P5 U509 ( .A1(n84), .A2(n142), .B1(n81), .B2(n143), .C1(n83), 
        .C2(n144), .X(n141) );
  SEN_OAI221_0P5 U510 ( .A1(n61), .A2(n137), .B1(n331), .B2(n44), .C(n39), .X(
        n143) );
  SEN_INV_1 U511 ( .A(n107), .X(n24) );
  SEN_INV_1 U512 ( .A(n112), .X(n50) );
  SEN_OR2_DG_1 U513 ( .A1(n86), .A2(n130), .X(n339) );
  SEN_AO222_1 U514 ( .A1(n31), .A2(n79), .B1(n133), .B2(n80), .C1(n135), .C2(
        n123), .X(n335) );
  SEN_AOI22_0P5 U515 ( .A1(n346), .A2(X[15]), .B1(n246), .B2(X[31]), .X(n229)
         );
  SEN_OR2_DG_1 U516 ( .A1(n203), .A2(n317), .X(n329) );
  SEN_OR2_DG_1 U517 ( .A1(n161), .A2(n281), .X(n330) );
  SEN_INV_S_6 U518 ( .A(n74), .X(n331) );
  SEN_NR2_S_0P5 U519 ( .A1(n102), .A2(n73), .X(n243) );
  SEN_INV_1 U520 ( .A(n168), .X(n22) );
  SEN_INV_2 U521 ( .A(n209), .X(n20) );
  SEN_INV_2 U522 ( .A(n201), .X(n15) );
  SEN_INV_2 U523 ( .A(n213), .X(n8) );
  SEN_NR2_S_0P5 U524 ( .A1(n331), .A2(n173), .X(n160) );
  SEN_OAI221_0P5 U525 ( .A1(n73), .A2(n44), .B1(n331), .B2(n61), .C(n216), .X(
        n164) );
  SEN_OAI221_0P5 U526 ( .A1(n70), .A2(n137), .B1(n331), .B2(n54), .C(n39), .X(
        n171) );
  SEN_AOI221_1 U527 ( .A1(n23), .A2(n79), .B1(n144), .B2(n81), .C(n185), .X(
        n168) );
  SEN_INV_S_0P5 U528 ( .A(n191), .X(n21) );
  SEN_INV_S_0P5 U529 ( .A(n92), .X(n2) );
  SEN_INV_S_0P5 U530 ( .A(n183), .X(n16) );
  SEN_INV_S_0P5 U531 ( .A(n94), .X(n7) );
  SEN_INV_S_0P5 U532 ( .A(n221), .X(n14) );
  SEN_INV_S_0P5 U533 ( .A(n110), .X(n6) );
  SEN_INV_S_0P5 U534 ( .A(n179), .X(n10) );
  SEN_INV_S_0P5 U535 ( .A(n117), .X(n25) );
  SEN_INV_S_0P5 U536 ( .A(n227), .X(n19) );
  SEN_INV_S_0P5 U537 ( .A(n224), .X(n3) );
  SEN_INV_S_0P5 U538 ( .A(n95), .X(n26) );
  SEN_INV_S_0P5 U539 ( .A(n97), .X(n12) );
  SEN_INV_1 U540 ( .A(n146), .X(n41) );
  SEN_INV_1 U541 ( .A(n190), .X(n37) );
  SEN_OR2_DG_1 U542 ( .A1(n75), .A2(n342), .X(n341) );
  SEN_AOI221_0P5 U543 ( .A1(X[28]), .A2(n337), .B1(n78), .B2(X[12]), .C(n152), 
        .X(n150) );
  SEN_INV_S_0P5 U544 ( .A(n151), .X(n36) );
  SEN_OAI222_0P5 U545 ( .A1(n155), .A2(n261), .B1(n156), .B2(n281), .C1(n35), 
        .C2(n123), .X(n140) );
  SEN_AOI221_0P5 U546 ( .A1(X[27]), .A2(n336), .B1(n78), .B2(X[11]), .C(n152), 
        .X(n156) );
  SEN_ND2_S_0P5 U547 ( .A1(n343), .A2(n342), .X(n251) );
  SEN_INV_S_0P5 U548 ( .A(n167), .X(n27) );
  SEN_AOI22_0P5 U549 ( .A1(n345), .A2(X[12]), .B1(n246), .B2(X[28]), .X(n116)
         );
  SEN_OAI221_0P5 U550 ( .A1(n126), .A2(n260), .B1(n127), .B2(n84), .C(n250), 
        .X(n198) );
  SEN_AOI22_0P5 U551 ( .A1(n345), .A2(X[14]), .B1(n246), .B2(X[30]), .X(n232)
         );
  SEN_AOI22_0P5 U552 ( .A1(n345), .A2(X[11]), .B1(n246), .B2(X[27]), .X(n121)
         );
  SEN_AOI22_0P5 U553 ( .A1(n346), .A2(X[10]), .B1(n246), .B2(X[26]), .X(n126)
         );
  SEN_AOI22_0P5 U554 ( .A1(n345), .A2(X[9]), .B1(n246), .B2(X[25]), .X(n101)
         );
  SEN_AOI22_0P5 U555 ( .A1(n346), .A2(X[8]), .B1(n246), .B2(n344), .X(n112) );
  SEN_AO221_0P5 U556 ( .A1(n345), .A2(X[16]), .B1(n337), .B2(X[0]), .C(n32), 
        .X(n115) );
  SEN_INV_S_0P5 U557 ( .A(n208), .X(n4) );
  SEN_AOI222_0P5 U558 ( .A1(n123), .A2(n200), .B1(n244), .B2(X[16]), .C1(n80), 
        .C2(n50), .X(n240) );
  SEN_BUF_6 U559 ( .A(LEFT), .X(n342) );
  SEN_OAI211_1 U560 ( .A1(n65), .A2(n158), .B1(n39), .B2(n165), .X(n142) );
  SEN_BUF_1 U561 ( .A(S[0]), .X(n343) );
  SEN_INV_1 U562 ( .A(n181), .X(n31) );
  SEN_INV_S_1 U563 ( .A(n338), .X(n350) );
  SEN_INV_S_1 U564 ( .A(n171), .X(n38) );
  SEN_OR2_1 U565 ( .A1(n85), .A2(n86), .X(n338) );
  SEN_ND2_G_1 U566 ( .A1(n197), .A2(n85), .X(n238) );
  SEN_INV_S_1 U567 ( .A(n339), .X(n348) );
  SEN_OAI221_1 U568 ( .A1(n188), .A2(n317), .B1(n38), .B2(n281), .C(n189), .X(
        n179) );
  SEN_OA2BB2_1 U569 ( .A1(n80), .A2(n28), .B1(n261), .B2(n203), .X(n218) );
  SEN_OAI221_1 U570 ( .A1(n103), .A2(n317), .B1(n166), .B2(n281), .C(n206), 
        .X(n191) );
  SEN_OAI221_1 U571 ( .A1(n232), .A2(n317), .B1(n219), .B2(n280), .C(n233), 
        .X(n224) );
  SEN_OA2BB2_1 U572 ( .A1(n80), .A2(n115), .B1(n108), .B2(n116), .X(n114) );
  SEN_OAI221_1 U573 ( .A1(n68), .A2(n137), .B1(n331), .B2(n52), .C(n39), .X(
        n133) );
  SEN_OAI222_1 U574 ( .A1(n343), .A2(n128), .B1(n129), .B2(n86), .C1(n40), 
        .C2(n351), .X(Z[31]) );
  SEN_OAI221_0P5 U575 ( .A1(n331), .A2(n42), .B1(n137), .B2(n60), .C(n39), .X(
        n134) );
  SEN_OAI221_1 U576 ( .A1(n118), .A2(n354), .B1(n70), .B2(n351), .C(n119), .X(
        Z[4]) );
  SEN_AOI222_1 U577 ( .A1(n316), .A2(n110), .B1(n349), .B2(n117), .C1(n348), 
        .C2(n275), .X(n119) );
  SEN_OAI221_1 U578 ( .A1(n138), .A2(n354), .B1(n42), .B2(n351), .C(n139), .X(
        Z[30]) );
  SEN_OA2BB2_1 U579 ( .A1(n316), .A2(n131), .B1(n86), .B2(n128), .X(n139) );
  SEN_AOI222_1 U580 ( .A1(n316), .A2(n335), .B1(n349), .B2(n34), .C1(n348), 
        .C2(n140), .X(n154) );
  SEN_OAI221_1 U581 ( .A1(n6), .A2(n354), .B1(n68), .B2(n351), .C(n100), .X(
        Z[6]) );
  SEN_AOI222_1 U582 ( .A1(n316), .A2(n97), .B1(n349), .B2(n275), .C1(n348), 
        .C2(n95), .X(n100) );
  SEN_OAI221_1 U583 ( .A1(n18), .A2(n354), .B1(n67), .B2(n351), .C(n98), .X(
        Z[7]) );
  SEN_INV_S_1 U584 ( .A(n275), .X(n18) );
  SEN_AOI222_1 U585 ( .A1(n316), .A2(n95), .B1(n349), .B2(n97), .C1(n348), 
        .C2(n92), .X(n98) );
  SEN_OAI221_1 U586 ( .A1(n25), .A2(n354), .B1(n69), .B2(n351), .C(n111), .X(
        Z[5]) );
  SEN_INV_1 U587 ( .A(n219), .X(n28) );
  SEN_OAI221_1 U588 ( .A1(n10), .A2(n354), .B1(n49), .B2(n352), .C(n174), .X(
        Z[24]) );
  SEN_INV_S_1 U589 ( .A(n344), .X(n49) );
  SEN_OAI221_1 U590 ( .A1(n26), .A2(n353), .B1(n65), .B2(n352), .C(n89), .X(
        Z[9]) );
  SEN_AOI222_1 U591 ( .A1(n355), .A2(n90), .B1(n350), .B2(n92), .C1(n347), 
        .C2(n94), .X(n89) );
  SEN_OAI221_1 U592 ( .A1(n2), .A2(n353), .B1(n64), .B2(n351), .C(n234), .X(
        Z[10]) );
  SEN_AOI222_1 U593 ( .A1(n316), .A2(n94), .B1(n349), .B2(n90), .C1(n348), 
        .C2(n227), .X(n234) );
  SEN_OAI221_1 U594 ( .A1(n284), .A2(n353), .B1(n54), .B2(n352), .C(n192), .X(
        Z[20]) );
  SEN_AOI222_1 U595 ( .A1(n355), .A2(n186), .B1(n350), .B2(n191), .C1(n347), 
        .C2(n183), .X(n192) );
  SEN_OAI221_1 U596 ( .A1(n21), .A2(n353), .B1(n53), .B2(n352), .C(n187), .X(
        Z[21]) );
  SEN_OAI221_1 U597 ( .A1(n16), .A2(n354), .B1(n51), .B2(n352), .C(n180), .X(
        Z[23]) );
  SEN_AOI222_1 U598 ( .A1(n355), .A2(n22), .B1(n350), .B2(n179), .C1(n347), 
        .C2(n167), .X(n180) );
  SEN_OAI221_1 U599 ( .A1(n7), .A2(n353), .B1(n62), .B2(n352), .C(n228), .X(
        Z[12]) );
  SEN_AOI222_1 U600 ( .A1(n316), .A2(n224), .B1(n349), .B2(n227), .C1(n348), 
        .C2(n221), .X(n228) );
  SEN_OAI221_1 U601 ( .A1(n19), .A2(n353), .B1(n61), .B2(n352), .C(n225), .X(
        Z[13]) );
  SEN_AOI222_1 U602 ( .A1(n355), .A2(n221), .B1(n350), .B2(n224), .C1(n347), 
        .C2(n8), .X(n225) );
  SEN_OAI221_1 U603 ( .A1(n3), .A2(n353), .B1(n60), .B2(n352), .C(n222), .X(
        Z[14]) );
  SEN_AOI222_1 U604 ( .A1(n355), .A2(n8), .B1(n350), .B2(n221), .C1(n347), 
        .C2(n20), .X(n222) );
  SEN_OAI221_1 U605 ( .A1(n14), .A2(n353), .B1(n59), .B2(n352), .C(n217), .X(
        Z[15]) );
  SEN_AOI222_1 U606 ( .A1(n355), .A2(n20), .B1(n350), .B2(n8), .C1(n347), .C2(
        n208), .X(n217) );
  SEN_OAI221_1 U607 ( .A1(n5), .A2(n353), .B1(n52), .B2(n352), .C(n184), .X(
        Z[22]) );
  SEN_OAI221_1 U608 ( .A1(n12), .A2(n354), .B1(n66), .B2(n351), .C(n96), .X(
        Z[8]) );
  SEN_AOI222_1 U609 ( .A1(n316), .A2(n92), .B1(n349), .B2(n95), .C1(n348), 
        .C2(n90), .X(n96) );
  SEN_INV_S_1 U610 ( .A(n343), .X(n86) );
  SEN_INV_S_1 U611 ( .A(n198), .X(n43) );
  SEN_AOI221_1 U612 ( .A1(n345), .A2(X[17]), .B1(n336), .B2(X[1]), .C(n32), 
        .X(n107) );
  SEN_AOI22_1 U613 ( .A1(n243), .A2(X[3]), .B1(n244), .B2(X[19]), .X(n249) );
  SEN_OA2BB2_1 U614 ( .A1(n160), .A2(X[26]), .B1(n82), .B2(n161), .X(n159) );
  SEN_AOI22_1 U615 ( .A1(n243), .A2(X[2]), .B1(n244), .B2(X[18]), .X(n250) );
  SEN_ND2_S_0P5 U616 ( .A1(n342), .A2(n253), .X(n252) );
  SEN_OAI221_1 U617 ( .A1(n213), .A2(n353), .B1(n58), .B2(n352), .C(n214), .X(
        Z[16]) );
  SEN_INV_S_1 U618 ( .A(X[16]), .X(n58) );
  SEN_OAI221_1 U619 ( .A1(n209), .A2(n353), .B1(n57), .B2(n352), .C(n210), .X(
        Z[17]) );
  SEN_INV_S_1 U620 ( .A(X[17]), .X(n57) );
  SEN_AOI222_1 U621 ( .A1(n355), .A2(n15), .B1(n350), .B2(n208), .C1(n347), 
        .C2(n195), .X(n210) );
  SEN_OAI22_1 U622 ( .A1(n41), .A2(n130), .B1(n242), .B2(n85), .X(n196) );
  SEN_AOI221_1 U623 ( .A1(n243), .A2(X[1]), .B1(n244), .B2(X[17]), .C(n245), 
        .X(n242) );
  SEN_INV_S_1 U624 ( .A(X[25]), .X(n48) );
  SEN_OAI221_1 U625 ( .A1(n201), .A2(n353), .B1(n55), .B2(n352), .C(n202), .X(
        Z[19]) );
  SEN_INV_S_1 U626 ( .A(X[19]), .X(n55) );
  SEN_AOI222_1 U627 ( .A1(n355), .A2(n191), .B1(n350), .B2(n195), .C1(n347), 
        .C2(n186), .X(n202) );
  SEN_OAI221_1 U628 ( .A1(n29), .A2(n354), .B1(n46), .B2(n351), .C(n157), .X(
        Z[27]) );
  SEN_INV_S_1 U629 ( .A(X[27]), .X(n46) );
  SEN_INV_S_1 U630 ( .A(X[3]), .X(n71) );
  SEN_OAI221_1 U631 ( .A1(n4), .A2(n353), .B1(n56), .B2(n352), .C(n205), .X(
        Z[18]) );
  SEN_INV_S_1 U632 ( .A(X[18]), .X(n56) );
  SEN_AOI222_1 U633 ( .A1(n355), .A2(n195), .B1(n350), .B2(n15), .C1(n347), 
        .C2(n191), .X(n205) );
  SEN_OAI221_1 U634 ( .A1(n13), .A2(n353), .B1(n63), .B2(n352), .C(n231), .X(
        Z[11]) );
  SEN_INV_S_1 U635 ( .A(X[11]), .X(n63) );
  SEN_INV_S_1 U636 ( .A(n90), .X(n13) );
  SEN_AOI222_1 U637 ( .A1(n316), .A2(n227), .B1(n349), .B2(n94), .C1(n348), 
        .C2(n224), .X(n231) );
  SEN_OAI221_1 U638 ( .A1(n27), .A2(n354), .B1(n47), .B2(n351), .C(n163), .X(
        Z[26]) );
  SEN_INV_S_1 U639 ( .A(X[26]), .X(n47) );
  SEN_AOI222_1 U640 ( .A1(n316), .A2(n33), .B1(n349), .B2(n162), .C1(n348), 
        .C2(n34), .X(n163) );
  SEN_OAI221_1 U641 ( .A1(n43), .A2(n354), .B1(n72), .B2(n351), .C(n145), .X(
        Z[2]) );
  SEN_INV_S_1 U642 ( .A(X[2]), .X(n72) );
  SEN_AOI222_1 U643 ( .A1(n316), .A2(n321), .B1(n349), .B2(n146), .C1(n348), 
        .C2(n117), .X(n145) );
  SEN_INV_S_1 U644 ( .A(X[28]), .X(n45) );
  SEN_INV_S_1 U645 ( .A(X[30]), .X(n42) );
  SEN_INV_S_1 U646 ( .A(X[29]), .X(n44) );
  SEN_INV_S_1 U647 ( .A(X[12]), .X(n62) );
  SEN_INV_S_1 U648 ( .A(X[14]), .X(n60) );
  SEN_INV_S_1 U649 ( .A(X[9]), .X(n65) );
  SEN_INV_S_1 U650 ( .A(X[8]), .X(n66) );
  SEN_INV_S_1 U651 ( .A(X[10]), .X(n64) );
  SEN_INV_S_1 U652 ( .A(X[13]), .X(n61) );
  SEN_INV_S_1 U653 ( .A(X[23]), .X(n51) );
  SEN_INV_S_1 U654 ( .A(X[20]), .X(n54) );
  SEN_INV_S_1 U655 ( .A(X[4]), .X(n70) );
  SEN_INV_S_1 U656 ( .A(X[21]), .X(n53) );
  SEN_INV_S_1 U657 ( .A(X[22]), .X(n52) );
  SEN_INV_S_1 U658 ( .A(X[15]), .X(n59) );
  SEN_INV_S_1 U659 ( .A(X[7]), .X(n67) );
  SEN_INV_S_1 U660 ( .A(X[5]), .X(n69) );
  SEN_INV_S_1 U661 ( .A(X[6]), .X(n68) );
  SEN_OAI211_1 U662 ( .A1(n67), .A2(n158), .B1(n39), .B2(n177), .X(n176) );
  SEN_BUF_S_1 U663 ( .A(X[24]), .X(n344) );
endmodule

