
module ShiftLR ( Z, X, S, LEFT, LOG, clock );
  output [31:0] Z;
  input [31:0] X;
  input [4:0] S;
  input LEFT, LOG, clock;
  wire   clocked_left, clocked_log, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249;
  wire   [31:0] clocked_input;
  wire   [4:0] clocked_shift;

  SEN_FDPQ_D_1 \clocked_input_reg[7]  ( .D(X[7]), .CK(clock), .Q(
        clocked_input[7]) );
  SEN_FDPQ_D_1 \clocked_input_reg[6]  ( .D(X[6]), .CK(clock), .Q(
        clocked_input[6]) );
  SEN_FDPQ_D_1 \clocked_input_reg[5]  ( .D(X[5]), .CK(clock), .Q(
        clocked_input[5]) );
  SEN_FDPQ_D_1 \clocked_input_reg[4]  ( .D(X[4]), .CK(clock), .Q(
        clocked_input[4]) );
  SEN_FDPQ_D_1 clocked_log_reg ( .D(LOG), .CK(clock), .Q(clocked_log) );
  SEN_FDPQ_D_1 \clocked_input_reg[3]  ( .D(X[3]), .CK(clock), .Q(
        clocked_input[3]) );
  SEN_FDPQ_D_1 \clocked_input_reg[2]  ( .D(X[2]), .CK(clock), .Q(
        clocked_input[2]) );
  SEN_FDPQ_D_1 \clocked_input_reg[1]  ( .D(X[1]), .CK(clock), .Q(
        clocked_input[1]) );
  SEN_FDPQ_D_1 \clocked_input_reg[0]  ( .D(X[0]), .CK(clock), .Q(
        clocked_input[0]) );
  SEN_FDPQ_D_1 \clocked_input_reg[23]  ( .D(X[23]), .CK(clock), .Q(
        clocked_input[23]) );
  SEN_FDPQ_D_1 \clocked_input_reg[22]  ( .D(X[22]), .CK(clock), .Q(
        clocked_input[22]) );
  SEN_FDPQ_D_1 \clocked_input_reg[21]  ( .D(X[21]), .CK(clock), .Q(
        clocked_input[21]) );
  SEN_FDPQ_D_1 \clocked_input_reg[20]  ( .D(X[20]), .CK(clock), .Q(
        clocked_input[20]) );
  SEN_FDPQ_D_1 \clocked_input_reg[30]  ( .D(X[30]), .CK(clock), .Q(
        clocked_input[30]) );
  SEN_FDPQ_D_1 \clocked_input_reg[29]  ( .D(X[29]), .CK(clock), .Q(
        clocked_input[29]) );
  SEN_FDPQ_D_1 \clocked_input_reg[28]  ( .D(X[28]), .CK(clock), .Q(
        clocked_input[28]) );
  SEN_FDPQ_D_1 \clocked_input_reg[15]  ( .D(X[15]), .CK(clock), .Q(
        clocked_input[15]) );
  SEN_FDPQ_D_1 \clocked_input_reg[14]  ( .D(X[14]), .CK(clock), .Q(
        clocked_input[14]) );
  SEN_FDPQ_D_1 \clocked_input_reg[13]  ( .D(X[13]), .CK(clock), .Q(
        clocked_input[13]) );
  SEN_FDPQ_D_1 \clocked_input_reg[12]  ( .D(X[12]), .CK(clock), .Q(
        clocked_input[12]) );
  SEN_FDPQB_D_1 \clocked_input_reg[19]  ( .D(X[19]), .CK(clock), .QN(n33) );
  SEN_FDPQB_D_1 \clocked_input_reg[18]  ( .D(X[18]), .CK(clock), .QN(n34) );
  SEN_FDPQB_D_1 \clocked_input_reg[17]  ( .D(X[17]), .CK(clock), .QN(n35) );
  SEN_FDPQB_D_1 \clocked_input_reg[16]  ( .D(X[16]), .CK(clock), .QN(n36) );
  SEN_FDPQ_D_1 \clocked_input_reg[11]  ( .D(X[11]), .CK(clock), .Q(
        clocked_input[11]) );
  SEN_FDPQ_D_1 \clocked_input_reg[10]  ( .D(X[10]), .CK(clock), .Q(
        clocked_input[10]) );
  SEN_FDPQ_D_1 \clocked_input_reg[9]  ( .D(X[9]), .CK(clock), .Q(
        clocked_input[9]) );
  SEN_FDPQ_D_1 \clocked_input_reg[8]  ( .D(X[8]), .CK(clock), .Q(
        clocked_input[8]) );
  SEN_FDPQ_D_1 \clocked_input_reg[27]  ( .D(X[27]), .CK(clock), .Q(
        clocked_input[27]) );
  SEN_FDPQ_D_1 \clocked_input_reg[31]  ( .D(X[31]), .CK(clock), .Q(
        clocked_input[31]) );
  SEN_FDPQ_D_1 \clocked_input_reg[26]  ( .D(X[26]), .CK(clock), .Q(
        clocked_input[26]) );
  SEN_FDPQ_D_1 \clocked_input_reg[25]  ( .D(X[25]), .CK(clock), .Q(
        clocked_input[25]) );
  SEN_FDPQ_D_1 \clocked_input_reg[24]  ( .D(X[24]), .CK(clock), .Q(
        clocked_input[24]) );
  SEN_FDPQ_D_1 \clocked_shift_reg[4]  ( .D(S[4]), .CK(clock), .Q(
        clocked_shift[4]) );
  SEN_FDPQB_3 \clocked_shift_reg[2]  ( .D(S[2]), .CK(clock), .QN(n48) );
  SEN_NR2_1 U224 ( .A1(n107), .A2(n217), .X(n173) );
  SEN_ND2_G_1 U225 ( .A1(n45), .A2(n47), .X(n145) );
  SEN_OAI22_1 U226 ( .A1(n100), .A2(n9), .B1(n101), .B2(n3), .X(n123) );
  SEN_INV_2 U227 ( .A(n196), .X(n241) );
  SEN_AOI22_0P75 U228 ( .A1(clocked_input[5]), .A2(n233), .B1(
        clocked_input[21]), .B2(n241), .X(n185) );
  SEN_INV_2 U229 ( .A(n232), .X(n233) );
  SEN_ND2_0P8 U230 ( .A1(n248), .A2(n225), .X(n107) );
  SEN_AN2_S_1 U232 ( .A1(n49), .A2(n159), .X(n230) );
  SEN_OAI222_1 U233 ( .A1(n17), .A2(n244), .B1(n112), .B2(n145), .C1(n164), 
        .C2(n47), .X(n159) );
  SEN_OR2_1 U234 ( .A1(n15), .A2(n81), .X(n243) );
  SEN_OAI221_1 U235 ( .A1(n112), .A2(n107), .B1(n17), .B2(n237), .C(n153), .X(
        n135) );
  SEN_OAI221_0P5 U236 ( .A1(n7), .A2(n82), .B1(n150), .B2(n81), .C(n151), .X(
        Z[15]) );
  SEN_AN2_DG_1 U237 ( .A1(n52), .A2(n162), .X(n231) );
  SEN_OA2BB2_1 U238 ( .A1(n51), .A2(n162), .B1(n63), .B2(n51), .X(n56) );
  SEN_NR2_S_2 U239 ( .A1(n230), .A2(n231), .X(n161) );
  SEN_AN2_S_0P5 U240 ( .A1(S[3]), .A2(n54), .X(n205) );
  SEN_AN2_1 U241 ( .A1(n193), .A2(clocked_left), .X(n206) );
  SEN_INV_2 U242 ( .A(n217), .X(n245) );
  SEN_EO2_1 U243 ( .A1(n48), .A2(n194), .X(n195) );
  SEN_AO21B_1 U244 ( .A1(n245), .A2(clocked_input[23]), .B(n154), .X(n148) );
  SEN_ND3_1 U245 ( .A1(n221), .A2(n222), .A3(n187), .X(n86) );
  SEN_NR3_G_1 U246 ( .A1(n210), .A2(n211), .A3(n212), .X(n68) );
  SEN_AN2_S_0P5 U247 ( .A1(n225), .A2(n138), .X(n212) );
  SEN_INV_1 U248 ( .A(n145), .X(n44) );
  SEN_ND2_G_1 U249 ( .A1(n44), .A2(n84), .X(n125) );
  SEN_BUF_2 U250 ( .A(n98), .X(n237) );
  SEN_INV_1 U251 ( .A(n67), .X(n47) );
  SEN_NR2_S_0P5 U252 ( .A1(n98), .A2(n217), .X(n174) );
  SEN_NR2_S_2 U253 ( .A1(clocked_shift[1]), .A2(clocked_shift[0]), .X(n194) );
  SEN_INV_S_1 U254 ( .A(n191), .X(n213) );
  SEN_INV_S_1 U255 ( .A(n121), .X(n20) );
  SEN_NR3_G_1 U256 ( .A1(n199), .A2(n200), .A3(n201), .X(n183) );
  SEN_AN2_S_1 U257 ( .A1(clocked_input[1]), .A2(n174), .X(n201) );
  SEN_INV_S_1 U258 ( .A(n136), .X(n9) );
  SEN_ND2_G_1 U259 ( .A1(n234), .A2(n132), .X(n115) );
  SEN_INV_S_1 U260 ( .A(n124), .X(n3) );
  SEN_ND2_G_1 U261 ( .A1(n51), .A2(n55), .X(n82) );
  SEN_OAI22_1 U262 ( .A1(n56), .A2(n55), .B1(n247), .B2(n57), .X(Z[9]) );
  SEN_AO221_1 U263 ( .A1(n106), .A2(n53), .B1(n103), .B2(n50), .C(n110), .X(
        Z[23]) );
  SEN_ND2_G_1 U264 ( .A1(n228), .A2(n229), .X(n110) );
  SEN_OR2_1 U265 ( .A1(n81), .A2(n3), .X(n229) );
  SEN_OR2_1 U266 ( .A1(n82), .A2(n10), .X(n228) );
  SEN_OR2_1 U267 ( .A1(n225), .A2(n245), .X(n196) );
  SEN_OR2_1 U268 ( .A1(clocked_log), .A2(clocked_left), .X(n197) );
  SEN_AN2_1 U269 ( .A1(n243), .A2(n242), .X(n198) );
  SEN_NR3_1 U270 ( .A1(n207), .A2(n208), .A3(n209), .X(n72) );
  SEN_OAI211_1 U271 ( .A1(n120), .A2(n244), .B1(n125), .B2(n140), .X(n122) );
  SEN_AOI222_1 U272 ( .A1(n241), .A2(clocked_input[26]), .B1(n233), .B2(
        clocked_input[10]), .C1(n225), .C2(n165), .X(n79) );
  SEN_OAI221_0P5 U273 ( .A1(n36), .A2(n170), .B1(n248), .B2(n31), .C(n179), 
        .X(n169) );
  SEN_OA22_DG_1 U274 ( .A1(n248), .A2(n164), .B1(n79), .B2(n47), .X(n63) );
  SEN_OA22_DG_1 U275 ( .A1(n248), .A2(n68), .B1(n69), .B2(n47), .X(n61) );
  SEN_OA22_DG_1 U276 ( .A1(n29), .A2(n47), .B1(n248), .B2(n69), .X(n75) );
  SEN_AOI22_1 U277 ( .A1(S[2]), .A2(n54), .B1(n195), .B2(clocked_left), .X(n67) );
  SEN_OA2BB2_1 U278 ( .A1(n129), .A2(n249), .B1(n249), .B2(n78), .X(n85) );
  SEN_OA22_DG_1 U279 ( .A1(n249), .A2(n157), .B1(n60), .B2(n51), .X(n163) );
  SEN_ND2_G_1 U280 ( .A1(n249), .A2(n55), .X(n81) );
  SEN_AOI22_0P75 U281 ( .A1(n86), .A2(n51), .B1(n249), .B2(n182), .X(n128) );
  SEN_OA22_DG_1 U282 ( .A1(n249), .A2(n66), .B1(n75), .B2(n51), .X(n70) );
  SEN_ND2_S_1 U283 ( .A1(n194), .A2(n48), .X(n192) );
  SEN_OAI222_0P5 U284 ( .A1(n14), .A2(n244), .B1(n120), .B2(n145), .C1(n72), 
        .C2(n47), .X(n162) );
  SEN_OAI221_1 U285 ( .A1(n20), .A2(n244), .B1(n120), .B2(n237), .C(n109), .X(
        n106) );
  SEN_AN2_S_1 U286 ( .A1(n172), .A2(clocked_input[25]), .X(n199) );
  SEN_AN2_DG_1 U287 ( .A1(n173), .A2(clocked_input[9]), .X(n200) );
  SEN_NR2_S_0P65 U288 ( .A1(n107), .A2(n245), .X(n172) );
  SEN_NR2_S_5 U290 ( .A1(n205), .A2(n206), .X(n167) );
  SEN_AN2_DG_1 U291 ( .A1(n241), .A2(clocked_input[30]), .X(n202) );
  SEN_AN2_S_0P5 U292 ( .A1(n233), .A2(clocked_input[14]), .X(n203) );
  SEN_AN2_S_0P5 U293 ( .A1(n225), .A2(n133), .X(n204) );
  SEN_NR3_G_1 U294 ( .A1(n202), .A2(n203), .A3(n204), .X(n164) );
  SEN_BUF_3 U295 ( .A(n67), .X(n248) );
  SEN_INV_S_1 U296 ( .A(clocked_left), .X(n54) );
  SEN_INV_S_0P5 U297 ( .A(n167), .X(n45) );
  SEN_AN2_S_0P5 U298 ( .A1(n241), .A2(clocked_input[28]), .X(n207) );
  SEN_AN2_S_0P5 U299 ( .A1(n233), .A2(clocked_input[12]), .X(n208) );
  SEN_AN2_S_0P5 U300 ( .A1(n225), .A2(n141), .X(n209) );
  SEN_OAI22_S_0P5 U301 ( .A1(n163), .A2(n55), .B1(n247), .B2(n56), .X(Z[10])
         );
  SEN_ND2_3 U302 ( .A1(n84), .A2(n217), .X(n154) );
  SEN_AN2_3 U303 ( .A1(n48), .A2(n224), .X(n223) );
  SEN_INV_1 U304 ( .A(clocked_shift[3]), .X(n224) );
  SEN_ND2_T_2 U305 ( .A1(n194), .A2(n223), .X(n191) );
  SEN_AN2_S_1 U306 ( .A1(n241), .A2(clocked_input[29]), .X(n210) );
  SEN_AN2_S_0P5 U307 ( .A1(n233), .A2(clocked_input[13]), .X(n211) );
  SEN_OAI22_1 U308 ( .A1(n57), .A2(n55), .B1(n247), .B2(n58), .X(Z[8]) );
  SEN_OA22_DG_1 U309 ( .A1(n249), .A2(n60), .B1(n61), .B2(n51), .X(n57) );
  SEN_ND2_1P5 U310 ( .A1(n191), .A2(n214), .X(n215) );
  SEN_ND2_4 U311 ( .A1(n213), .A2(clocked_shift[4]), .X(n216) );
  SEN_ND2_S_4 U312 ( .A1(n215), .A2(n216), .X(n190) );
  SEN_INV_0P8 U313 ( .A(clocked_shift[4]), .X(n214) );
  SEN_AO22_8 U314 ( .A1(S[4]), .A2(n54), .B1(n190), .B2(clocked_left), .X(n217) );
  SEN_AN2_S_0P5 U315 ( .A1(n241), .A2(clocked_input[27]), .X(n218) );
  SEN_AN2_S_0P5 U316 ( .A1(n233), .A2(clocked_input[11]), .X(n219) );
  SEN_AN2_S_0P5 U317 ( .A1(n225), .A2(n147), .X(n220) );
  SEN_NR3_G_1 U318 ( .A1(n218), .A2(n219), .A3(n220), .X(n76) );
  SEN_OAI22_T_0P5 U319 ( .A1(n85), .A2(n55), .B1(n247), .B2(n128), .X(Z[1]) );
  SEN_OR2_1 U320 ( .A1(n33), .A2(n170), .X(n221) );
  SEN_OR2_DG_1 U321 ( .A1(n248), .A2(n6), .X(n222) );
  SEN_OA2BB2_1 U322 ( .A1(n86), .A2(n249), .B1(n249), .B2(n75), .X(n77) );
  SEN_OR2_DG_1 U323 ( .A1(n157), .A2(n100), .X(n226) );
  SEN_OR2_DG_1 U324 ( .A1(n150), .A2(n101), .X(n227) );
  SEN_ND3_S_1 U325 ( .A1(n226), .A2(n227), .A3(n161), .X(Z[12]) );
  SEN_ND2_S_0P5 U326 ( .A1(n247), .A2(n59), .X(n100) );
  SEN_AOI222_1 U327 ( .A1(n147), .A2(n46), .B1(n127), .B2(n44), .C1(n5), .C2(
        n248), .X(n150) );
  SEN_BUF_1 U328 ( .A(n111), .X(n244) );
  SEN_AOI22_0P75 U329 ( .A1(n49), .A2(n103), .B1(n52), .B2(n106), .X(n105) );
  SEN_INV_1 U330 ( .A(n159), .X(n15) );
  SEN_NR2_1 U331 ( .A1(n235), .A2(n236), .X(n131) );
  SEN_AOI22_0P5 U332 ( .A1(n53), .A2(n115), .B1(n50), .B2(n106), .X(n119) );
  SEN_ND2_G_1 U333 ( .A1(n155), .A2(n198), .X(Z[14]) );
  SEN_INV_S_2 U334 ( .A(n88), .X(n232) );
  SEN_AOI22_S_1 U336 ( .A1(n49), .A2(n95), .B1(n52), .B2(n103), .X(n102) );
  SEN_AN2_1 U337 ( .A1(n53), .A2(n122), .X(n235) );
  SEN_OAI22_T_0P5 U338 ( .A1(n74), .A2(n55), .B1(n247), .B2(n77), .X(Z[3]) );
  SEN_OR3_1 U339 ( .A1(n238), .A2(n239), .A3(n240), .X(n103) );
  SEN_AOI22_0P5 U340 ( .A1(n43), .A2(n113), .B1(n42), .B2(n133), .X(n132) );
  SEN_OA21_1 U341 ( .A1(n112), .A2(n244), .B(n125), .X(n234) );
  SEN_AOI22_0P5 U342 ( .A1(n53), .A2(n159), .B1(n50), .B2(n152), .X(n158) );
  SEN_INV_1 U343 ( .A(n237), .X(n42) );
  SEN_OAI221_1 U344 ( .A1(n9), .A2(n82), .B1(n2), .B2(n81), .C(n131), .X(Z[19]) );
  SEN_NR2_S_0P5 U345 ( .A1(n24), .A2(n244), .X(n238) );
  SEN_OA22_DG_1 U346 ( .A1(n248), .A2(n72), .B1(n73), .B2(n47), .X(n64) );
  SEN_OA22_DG_1 U347 ( .A1(n27), .A2(n47), .B1(n248), .B2(n79), .X(n71) );
  SEN_OA22_DG_1 U348 ( .A1(n31), .A2(n47), .B1(n248), .B2(n73), .X(n78) );
  SEN_AN2_1 U349 ( .A1(n50), .A2(n115), .X(n236) );
  SEN_INV_1 U350 ( .A(n100), .X(n53) );
  SEN_INV_1 U351 ( .A(n101), .X(n50) );
  SEN_OAI22_T_0P5 U352 ( .A1(n77), .A2(n55), .B1(n247), .B2(n85), .X(Z[2]) );
  SEN_INV_S_1 U353 ( .A(n113), .X(n24) );
  SEN_OAI21_T_0P5 U354 ( .A1(n128), .A2(n55), .B(n168), .X(Z[0]) );
  SEN_AOI22_S_1 U355 ( .A1(n52), .A2(n169), .B1(n49), .B2(n129), .X(n168) );
  SEN_NR2_S_0P5 U356 ( .A1(n112), .A2(n237), .X(n239) );
  SEN_INV_S_1 U357 ( .A(n109), .X(n240) );
  SEN_ND2_S_0P5 U358 ( .A1(n248), .A2(n167), .X(n98) );
  SEN_AOI22_1 U359 ( .A1(n53), .A2(n103), .B1(n50), .B2(n95), .X(n104) );
  SEN_OA222_0P5 U360 ( .A1(n8), .A2(n244), .B1(n117), .B2(n145), .C1(n68), 
        .C2(n47), .X(n157) );
  SEN_ND2_S_0P5 U361 ( .A1(n167), .A2(n47), .X(n111) );
  SEN_INV_1 U362 ( .A(n93), .X(n21) );
  SEN_INV_1 U363 ( .A(n111), .X(n46) );
  SEN_AOI22_0P5 U364 ( .A1(n44), .A2(n113), .B1(n46), .B2(n133), .X(n153) );
  SEN_OAI21_S_0P5 U365 ( .A1(n217), .A2(n33), .B(n154), .X(n147) );
  SEN_OAI21_S_0P5 U366 ( .A1(n217), .A2(n34), .B(n154), .X(n165) );
  SEN_OR2_1 U367 ( .A1(n13), .A2(n82), .X(n242) );
  SEN_INV_S_0P5 U368 ( .A(n152), .X(n13) );
  SEN_AOI22_T_0P5 U369 ( .A1(n53), .A2(n152), .B1(n50), .B2(n135), .X(n151) );
  SEN_AOI22_0P75 U370 ( .A1(n53), .A2(n135), .B1(n50), .B2(n122), .X(n139) );
  SEN_INV_S_0P5 U371 ( .A(n135), .X(n16) );
  SEN_INV_S_0P5 U372 ( .A(n142), .X(n2) );
  SEN_ND2_S_0P5 U373 ( .A1(n84), .A2(n225), .X(n109) );
  SEN_AOI22_0P5 U374 ( .A1(n53), .A2(n91), .B1(n50), .B2(n84), .X(n90) );
  SEN_AOI21_S_0P5 U375 ( .A1(n83), .A2(n249), .B(n84), .X(n80) );
  SEN_AOI22_0P5 U376 ( .A1(n44), .A2(n118), .B1(n46), .B2(n138), .X(n156) );
  SEN_OAI21_G_0P5 U377 ( .A1(n247), .A2(n80), .B(n25), .X(Z[31]) );
  SEN_INV_S_0P5 U378 ( .A(n127), .X(n18) );
  SEN_INV_S_0P5 U379 ( .A(n148), .X(n11) );
  SEN_AOI222_0P5 U380 ( .A1(n241), .A2(clocked_input[24]), .B1(n233), .B2(
        clocked_input[8]), .C1(n130), .C2(n225), .X(n73) );
  SEN_OAI221_1 U381 ( .A1(n3), .A2(n82), .B1(n9), .B2(n81), .C(n119), .X(Z[21]) );
  SEN_OAI221_1 U382 ( .A1(n96), .A2(n82), .B1(n10), .B2(n81), .C(n104), .X(
        Z[25]) );
  SEN_AOI22_0P5 U383 ( .A1(n53), .A2(n95), .B1(n50), .B2(n91), .X(n97) );
  SEN_AOI22_0P5 U384 ( .A1(n43), .A2(n127), .B1(n42), .B2(n147), .X(n146) );
  SEN_INV_S_0P5 U385 ( .A(n84), .X(n25) );
  SEN_AOI22_0P5 U386 ( .A1(n43), .A2(n118), .B1(n42), .B2(n138), .X(n137) );
  SEN_OAI221_0P5 U387 ( .A1(n117), .A2(n107), .B1(n8), .B2(n237), .C(n156), 
        .X(n144) );
  SEN_OAI22_S_0P5 U388 ( .A1(n62), .A2(n55), .B1(n247), .B2(n65), .X(Z[6]) );
  SEN_AOI22_0P5 U389 ( .A1(clocked_input[4]), .A2(n233), .B1(clocked_input[20]), .B2(n241), .X(n181) );
  SEN_AOI22_0P5 U390 ( .A1(clocked_input[6]), .A2(n233), .B1(clocked_input[22]), .B2(n241), .X(n178) );
  SEN_AOI222_0P5 U391 ( .A1(n241), .A2(clocked_input[25]), .B1(n233), .B2(
        clocked_input[9]), .C1(n225), .C2(n89), .X(n69) );
  SEN_OR2_DG_1 U392 ( .A1(n217), .A2(n35), .X(n246) );
  SEN_ND2_S_0P5 U393 ( .A1(n246), .A2(n154), .X(n89) );
  SEN_INV_S_0P5 U394 ( .A(n89), .X(n8) );
  SEN_OAI21_S_0P5 U395 ( .A1(n24), .A2(n237), .B(n99), .X(n91) );
  SEN_OAI221_0P5 U396 ( .A1(n22), .A2(n244), .B1(n117), .B2(n237), .C(n109), 
        .X(n116) );
  SEN_ND2_S_0P5 U397 ( .A1(n84), .A2(n237), .X(n99) );
  SEN_NR2_T_1 U398 ( .A1(n26), .A2(n197), .X(n84) );
  SEN_INV_1 U399 ( .A(n91), .X(n23) );
  SEN_OAI21_S_0P5 U400 ( .A1(n94), .A2(n47), .B(n25), .X(n83) );
  SEN_OAI221_1 U401 ( .A1(n96), .A2(n100), .B1(n21), .B2(n101), .C(n102), .X(
        Z[26]) );
  SEN_OAI221_1 U402 ( .A1(n3), .A2(n100), .B1(n10), .B2(n101), .C(n114), .X(
        Z[22]) );
  SEN_ND2_S_0P5 U403 ( .A1(n42), .A2(n217), .X(n170) );
  SEN_AOI22_0P5 U404 ( .A1(n53), .A2(n93), .B1(n50), .B2(n83), .X(n92) );
  SEN_INV_S_0P5 U405 ( .A(n95), .X(n19) );
  SEN_OAI221_0P5 U406 ( .A1(n21), .A2(n82), .B1(n96), .B2(n81), .C(n97), .X(
        Z[27]) );
  SEN_ND2_S_0P5 U407 ( .A1(n225), .A2(n217), .X(n177) );
  SEN_AOI22_0P5 U408 ( .A1(n53), .A2(n144), .B1(n50), .B2(n142), .X(n143) );
  SEN_INV_1 U409 ( .A(n118), .X(n22) );
  SEN_OA22_1 U410 ( .A1(n101), .A2(n7), .B1(n100), .B2(n150), .X(n155) );
  SEN_OAI21_S_0P5 U411 ( .A1(n217), .A2(n32), .B(n154), .X(n121) );
  SEN_OAI21_S_0P5 U412 ( .A1(n217), .A2(n28), .B(n154), .X(n113) );
  SEN_OAI21_S_0P5 U413 ( .A1(n217), .A2(n30), .B(n154), .X(n118) );
  SEN_INV_S_0P5 U414 ( .A(n162), .X(n12) );
  SEN_OAI221_0P5 U415 ( .A1(n108), .A2(n145), .B1(n11), .B2(n244), .C(n146), 
        .X(n142) );
  SEN_OA2BB2_0P5 U416 ( .A1(n47), .A2(n5), .B1(n76), .B2(n47), .X(n60) );
  SEN_INV_S_0P5 U417 ( .A(n83), .X(n4) );
  SEN_ND2_S_0P5 U418 ( .A1(n245), .A2(n225), .X(n176) );
  SEN_OAI22_S_1 U419 ( .A1(n70), .A2(n55), .B1(n247), .B2(n74), .X(Z[4]) );
  SEN_OAI22_S_1 U420 ( .A1(n65), .A2(n55), .B1(n247), .B2(n70), .X(Z[5]) );
  SEN_OAI22_S_1 U421 ( .A1(n58), .A2(n55), .B1(n247), .B2(n62), .X(Z[7]) );
  SEN_OA22_1 U422 ( .A1(n249), .A2(n64), .B1(n71), .B2(n51), .X(n65) );
  SEN_OA22_1 U423 ( .A1(n249), .A2(n61), .B1(n66), .B2(n51), .X(n62) );
  SEN_OAI211_0P5 U424 ( .A1(n18), .A2(n244), .B1(n125), .B2(n126), .X(n124) );
  SEN_AOI21B_0P5 U425 ( .A1(n245), .A2(clocked_input[24]), .B(n154), .X(n120)
         );
  SEN_AOI21B_0P5 U426 ( .A1(n245), .A2(clocked_input[26]), .B(n154), .X(n112)
         );
  SEN_AOI21B_0P5 U427 ( .A1(n245), .A2(clocked_input[25]), .B(n154), .X(n117)
         );
  SEN_AOI21_S_0P5 U428 ( .A1(n245), .A2(clocked_input[31]), .B(n84), .X(n108)
         );
  SEN_BUF_S_1 U429 ( .A(S[0]), .X(n247) );
  SEN_OAI21_S_0P5 U430 ( .A1(n217), .A2(n36), .B(n154), .X(n130) );
  SEN_BUF_S_1 U431 ( .A(n59), .X(n249) );
  SEN_AOI22_0P5 U432 ( .A1(S[1]), .A2(n54), .B1(clocked_left), .B2(n186), .X(
        n59) );
  SEN_OAI221_1 U433 ( .A1(n120), .A2(n107), .B1(n14), .B2(n237), .C(n160), .X(
        n152) );
  SEN_OA22_DG_1 U434 ( .A1(n237), .A2(n11), .B1(n107), .B2(n108), .X(n126) );
  SEN_INV_S_0P5 U435 ( .A(n107), .X(n43) );
  SEN_INV_S_1 U436 ( .A(n82), .X(n49) );
  SEN_OAI21_S_0P5 U437 ( .A1(n20), .A2(n237), .B(n99), .X(n95) );
  SEN_INV_S_1 U438 ( .A(n81), .X(n52) );
  SEN_OAI222_1 U439 ( .A1(n23), .A2(n81), .B1(n25), .B2(n82), .C1(n80), .C2(
        n55), .X(Z[30]) );
  SEN_OAI221_1 U440 ( .A1(n150), .A2(n82), .B1(n157), .B2(n81), .C(n158), .X(
        Z[13]) );
  SEN_OAI21_S_0P5 U441 ( .A1(n22), .A2(n237), .B(n99), .X(n93) );
  SEN_AOI22_S_1 U442 ( .A1(n49), .A2(n106), .B1(n52), .B2(n115), .X(n114) );
  SEN_OAI221_0P5 U443 ( .A1(n10), .A2(n100), .B1(n96), .B2(n101), .C(n105), 
        .X(Z[24]) );
  SEN_OAI221_1 U444 ( .A1(n2), .A2(n82), .B1(n7), .B2(n81), .C(n139), .X(Z[17]) );
  SEN_OAI221_1 U445 ( .A1(n2), .A2(n100), .B1(n9), .B2(n101), .C(n134), .X(
        Z[18]) );
  SEN_AOI22_S_1 U446 ( .A1(n49), .A2(n122), .B1(n52), .B2(n135), .X(n134) );
  SEN_OAI221_1 U447 ( .A1(n16), .A2(n82), .B1(n13), .B2(n81), .C(n143), .X(
        Z[16]) );
  SEN_OAI221_1 U448 ( .A1(n23), .A2(n82), .B1(n19), .B2(n81), .C(n92), .X(
        Z[28]) );
  SEN_INV_S_1 U449 ( .A(n144), .X(n7) );
  SEN_AO221_1 U450 ( .A1(n115), .A2(n49), .B1(n122), .B2(n52), .C(n123), .X(
        Z[20]) );
  SEN_AOI22_S_1 U451 ( .A1(n43), .A2(n121), .B1(n42), .B2(n141), .X(n140) );
  SEN_AOI22_S_1 U452 ( .A1(n44), .A2(n121), .B1(n46), .B2(n141), .X(n160) );
  SEN_OAI222_1 U453 ( .A1(n15), .A2(n101), .B1(n12), .B2(n100), .C1(n247), 
        .C2(n163), .X(Z[11]) );
  SEN_ND2_G_1 U454 ( .A1(n247), .A2(n51), .X(n101) );
  SEN_OA222_0P5 U455 ( .A1(n18), .A2(n237), .B1(n25), .B2(n107), .C1(n248), 
        .C2(n94), .X(n96) );
  SEN_OAI221_1 U456 ( .A1(n4), .A2(n82), .B1(n21), .B2(n81), .C(n90), .X(Z[29]) );
  SEN_INV_S_1 U457 ( .A(n116), .X(n10) );
  SEN_OAI211_1 U458 ( .A1(n117), .A2(n244), .B1(n125), .B2(n137), .X(n136) );
  SEN_INV_S_1 U459 ( .A(S[0]), .X(n55) );
  SEN_OA22_DG_1 U460 ( .A1(n249), .A2(n63), .B1(n64), .B2(n51), .X(n58) );
  SEN_OA22_DG_1 U461 ( .A1(n249), .A2(n71), .B1(n78), .B2(n51), .X(n74) );
  SEN_OA22_DG_1 U462 ( .A1(n6), .A2(n47), .B1(n248), .B2(n76), .X(n66) );
  SEN_INV_S_1 U463 ( .A(n165), .X(n17) );
  SEN_INV_S_1 U464 ( .A(n130), .X(n14) );
  SEN_OA21_1 U465 ( .A1(n108), .A2(n225), .B(n109), .X(n94) );
  SEN_INV_1 U466 ( .A(n249), .X(n51) );
  SEN_OAI221_1 U467 ( .A1(n34), .A2(n170), .B1(n248), .B2(n27), .C(n171), .X(
        n129) );
  SEN_AOI222_1 U468 ( .A1(n172), .A2(clocked_input[26]), .B1(n173), .B2(
        clocked_input[10]), .C1(clocked_input[2]), .C2(n174), .X(n171) );
  SEN_AOI222_1 U469 ( .A1(n172), .A2(clocked_input[27]), .B1(n173), .B2(
        clocked_input[11]), .C1(clocked_input[3]), .C2(n174), .X(n187) );
  SEN_OAI221_1 U470 ( .A1(n35), .A2(n170), .B1(n248), .B2(n29), .C(n183), .X(
        n182) );
  SEN_EO2_S_0P5 U471 ( .A1(clocked_shift[1]), .A2(clocked_shift[0]), .X(n186)
         );
  SEN_AO21B_1 U472 ( .A1(n245), .A2(clocked_input[20]), .B(n154), .X(n141) );
  SEN_AO21B_1 U473 ( .A1(n245), .A2(clocked_input[21]), .B(n154), .X(n138) );
  SEN_AO21B_1 U474 ( .A1(n245), .A2(clocked_input[22]), .B(n154), .X(n133) );
  SEN_AO21B_1 U475 ( .A1(n245), .A2(clocked_input[27]), .B(n154), .X(n127) );
  SEN_INV_S_1 U476 ( .A(n166), .X(n5) );
  SEN_AOI222_1 U477 ( .A1(n241), .A2(clocked_input[31]), .B1(n233), .B2(
        clocked_input[15]), .C1(n225), .C2(n148), .X(n166) );
  SEN_INV_S_1 U478 ( .A(n180), .X(n31) );
  SEN_OAI221_1 U479 ( .A1(n40), .A2(n176), .B1(n32), .B2(n177), .C(n181), .X(
        n180) );
  SEN_INV_S_1 U480 ( .A(clocked_input[12]), .X(n40) );
  SEN_INV_S_1 U481 ( .A(n184), .X(n29) );
  SEN_OAI221_1 U482 ( .A1(n39), .A2(n176), .B1(n30), .B2(n177), .C(n185), .X(
        n184) );
  SEN_INV_S_1 U483 ( .A(clocked_input[13]), .X(n39) );
  SEN_INV_S_1 U484 ( .A(n175), .X(n27) );
  SEN_OAI221_1 U485 ( .A1(n38), .A2(n176), .B1(n28), .B2(n177), .C(n178), .X(
        n175) );
  SEN_INV_S_1 U486 ( .A(clocked_input[14]), .X(n38) );
  SEN_INV_S_1 U487 ( .A(n188), .X(n6) );
  SEN_OAI221_1 U488 ( .A1(n37), .A2(n176), .B1(n26), .B2(n177), .C(n189), .X(
        n188) );
  SEN_INV_S_1 U489 ( .A(clocked_input[15]), .X(n37) );
  SEN_AOI22_1 U490 ( .A1(clocked_input[7]), .A2(n233), .B1(clocked_input[23]), 
        .B2(n241), .X(n189) );
  SEN_INV_S_1 U491 ( .A(clocked_input[31]), .X(n26) );
  SEN_AOI222_1 U492 ( .A1(n172), .A2(clocked_input[24]), .B1(n173), .B2(
        clocked_input[8]), .C1(clocked_input[0]), .C2(n174), .X(n179) );
  SEN_INV_S_1 U493 ( .A(clocked_input[29]), .X(n30) );
  SEN_INV_S_1 U494 ( .A(clocked_input[28]), .X(n32) );
  SEN_INV_S_1 U495 ( .A(clocked_input[30]), .X(n28) );
  SEN_FDPQ_2 clocked_left_reg ( .D(LEFT), .CK(clock), .Q(clocked_left) );
  SEN_FDPQ_2 \clocked_shift_reg[3]  ( .D(S[3]), .CK(clock), .Q(
        clocked_shift[3]) );
  SEN_FDPQ_2 \clocked_shift_reg[1]  ( .D(S[1]), .CK(clock), .Q(
        clocked_shift[1]) );
  SEN_FDPQ_2 \clocked_shift_reg[0]  ( .D(S[0]), .CK(clock), .Q(
        clocked_shift[0]) );
  SEN_EO2_1 U231 ( .A1(n192), .A2(clocked_shift[3]), .X(n193) );
  SEN_NR2_1 U289 ( .A1(n217), .A2(n225), .X(n88) );
  SEN_INV_4 U335 ( .A(n167), .X(n225) );
endmodule

