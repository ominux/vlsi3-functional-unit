/*
 Testbench for the functional verification of the 
 functional unit top level using VCS simulator

 Author: Corey Olson
 Date: 4/29/2010
*/
module functional_unit_tb();

endmodule
