#----------------------------------------------------------------------------
# Description	: Cell LEF definitions for cp65npksdst
#		  (Common Platform 65nm LP LowK Std Vt High Density Tapless Library)
# Date		: $Date: 2008/11/28 11:38:38 $
# Copyright	: 1997-2008 by Virage Logic Corporation
# Revision	: Version $Revision: 1.7 $
#----------------------------------------------------------------------------

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

# Placement site definition for this library.
SITE cp65_dst
  SYMMETRY Y ;
  CLASS core ;
  SIZE 0.2 BY 1.8 ;
END cp65_dst

#----------------------------------------------------------------------------
# Cell macro definitions.
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_D_1
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_D_1
  CLASS CORE ;
  FOREIGN SEN_ADDF_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.24 0.71 0.45 0.88 ;
      RECT  0.35 0.88 0.45 1.07 ;
      RECT  0.35 1.07 0.84 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0585 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.885 ;
      RECT  0.55 0.885 1.05 0.975 ;
      RECT  0.95 0.975 1.05 1.185 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0585 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.31 0.91 5.41 1.34 ;
      RECT  2.325 0.78 2.425 1.115 ;
      RECT  2.325 1.115 2.55 1.21 ;
      LAYER M2 ;
      RECT  2.285 0.95 5.45 1.05 ;
      LAYER V1 ;
      RECT  5.31 0.95 5.41 1.05 ;
      RECT  2.325 0.95 2.425 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0837 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.245 2.85 1.05 ;
      RECT  2.73 1.05 2.85 1.25 ;
    END
    ANTENNADIFFAREA 0.143 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.5 5.95 0.69 ;
      RECT  5.75 0.69 5.85 1.42 ;
      RECT  5.75 1.42 5.95 1.6 ;
    END
    ANTENNADIFFAREA 0.139 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  5.52 0.98 5.645 1.22 ;
      RECT  5.555 1.22 5.645 1.75 ;
      RECT  0.045 1.465 0.215 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.565 1.465 0.735 1.75 ;
      RECT  2.47 1.44 2.6 1.75 ;
      RECT  3.22 1.44 3.35 1.75 ;
      RECT  3.77 1.4 3.9 1.75 ;
      RECT  4.28 1.43 4.41 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  0.575 0.05 0.745 0.2 ;
      RECT  1.165 0.05 1.335 0.2 ;
      RECT  4.29 0.05 4.42 0.25 ;
      RECT  3.31 0.05 3.44 0.36 ;
      RECT  2.47 0.05 2.6 0.39 ;
      RECT  5.56 0.05 5.69 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.555 0.23 5.45 0.32 ;
      RECT  4.555 0.32 4.645 0.34 ;
      RECT  5.36 0.32 5.45 0.58 ;
      RECT  4.04 0.34 4.645 0.43 ;
      RECT  4.04 0.43 4.48 0.51 ;
      RECT  4.39 0.51 4.48 0.63 ;
      RECT  4.39 0.63 4.53 0.8 ;
      RECT  4.39 0.8 4.48 1.25 ;
      RECT  4.025 1.25 4.62 1.34 ;
      RECT  4.53 1.34 4.62 1.455 ;
      RECT  4.025 1.34 4.145 1.52 ;
      RECT  4.53 1.455 4.95 1.575 ;
      RECT  0.06 0.29 1.525 0.38 ;
      RECT  1.435 0.38 1.525 0.46 ;
      RECT  0.06 0.38 0.175 0.48 ;
      RECT  0.06 0.48 0.15 1.285 ;
      RECT  0.06 1.285 1.16 1.375 ;
      RECT  1.055 1.375 1.16 1.57 ;
      RECT  0.34 1.375 0.44 1.6 ;
      RECT  1.055 1.57 2.085 1.66 ;
      RECT  1.915 1.48 2.085 1.57 ;
      RECT  1.925 0.285 2.045 0.455 ;
      RECT  1.925 0.455 2.025 1.31 ;
      RECT  0.87 0.5 1.18 0.555 ;
      RECT  0.87 0.555 1.385 0.59 ;
      RECT  1.09 0.59 1.385 0.645 ;
      RECT  1.285 0.645 1.385 1.3 ;
      RECT  1.285 1.3 1.455 1.48 ;
      RECT  2.195 0.2 2.305 0.575 ;
      RECT  2.115 0.575 2.305 0.665 ;
      RECT  2.115 0.665 2.235 1.3 ;
      RECT  2.115 1.3 2.325 1.39 ;
      RECT  2.205 1.39 2.325 1.58 ;
      RECT  2.395 0.51 2.495 0.59 ;
      RECT  2.395 0.59 2.655 0.69 ;
      RECT  2.555 0.69 2.655 0.985 ;
      RECT  3.775 0.2 3.895 0.6 ;
      RECT  3.56 0.6 4.235 0.69 ;
      RECT  4.145 0.69 4.235 0.83 ;
      RECT  3.56 0.69 3.65 0.99 ;
      RECT  3.48 0.99 3.65 1.13 ;
      RECT  2.98 0.19 3.07 0.64 ;
      RECT  2.98 0.64 3.445 0.73 ;
      RECT  3.355 0.73 3.445 0.87 ;
      RECT  2.98 0.73 3.07 1.515 ;
      RECT  5.075 0.41 5.18 0.73 ;
      RECT  5.075 0.73 5.66 0.82 ;
      RECT  5.49 0.82 5.66 0.84 ;
      RECT  5.075 0.82 5.195 1.16 ;
      RECT  4.85 0.44 4.955 0.89 ;
      RECT  4.67 0.52 4.76 0.99 ;
      RECT  4.57 0.99 4.76 1.07 ;
      RECT  4.57 1.07 4.895 1.16 ;
      RECT  4.805 1.16 4.895 1.25 ;
      RECT  4.805 1.25 5.16 1.34 ;
      RECT  5.07 1.34 5.16 1.515 ;
      RECT  5.07 1.515 5.465 1.61 ;
      RECT  5.345 1.43 5.465 1.515 ;
      RECT  1.475 0.685 1.585 1.21 ;
      RECT  3.74 1.135 3.83 1.22 ;
      RECT  3.49 1.22 3.83 1.31 ;
      RECT  3.49 1.31 3.59 1.51 ;
      RECT  1.695 0.27 1.795 1.32 ;
      RECT  1.59 1.32 1.795 1.44 ;
      RECT  3.16 0.885 3.26 1.335 ;
      LAYER M2 ;
      RECT  1.655 0.55 2.535 0.65 ;
      RECT  1.445 0.75 4.99 0.85 ;
      RECT  1.245 1.15 3.3 1.25 ;
      RECT  1.02 1.35 3.63 1.45 ;
      LAYER V1 ;
      RECT  1.695 0.55 1.795 0.65 ;
      RECT  2.395 0.55 2.495 0.65 ;
      RECT  1.485 0.75 1.585 0.85 ;
      RECT  2.115 0.75 2.215 0.85 ;
      RECT  4.85 0.75 4.95 0.85 ;
      RECT  1.285 1.15 1.385 1.25 ;
      RECT  1.925 1.15 2.025 1.25 ;
      RECT  3.16 1.15 3.26 1.25 ;
      RECT  1.06 1.35 1.16 1.45 ;
      RECT  3.49 1.35 3.59 1.45 ;
  END
END SEN_ADDF_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_D_2
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_D_2
  CLASS CORE ;
  FOREIGN SEN_ADDF_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.645 ;
      RECT  0.27 0.645 0.86 0.735 ;
      RECT  0.75 0.51 0.85 0.645 ;
      RECT  0.27 0.735 0.45 0.9 ;
      RECT  0.75 0.735 0.86 0.93 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.135 0.88 ;
      RECT  0.95 0.88 1.05 1.045 ;
      RECT  0.55 0.91 0.65 1.0 ;
      RECT  0.47 1.0 0.65 1.045 ;
      RECT  0.47 1.045 1.05 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1053 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.295 0.91 5.395 1.335 ;
      RECT  2.325 0.49 2.425 1.09 ;
      LAYER M2 ;
      RECT  2.285 0.95 5.435 1.05 ;
      LAYER V1 ;
      RECT  5.295 0.95 5.395 1.05 ;
      RECT  2.325 0.95 2.425 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.093 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.735 0.17 2.85 0.36 ;
      RECT  2.75 0.36 2.85 0.51 ;
      RECT  2.75 0.51 3.05 0.69 ;
      RECT  2.75 0.69 2.85 1.16 ;
      RECT  2.505 1.16 2.85 1.25 ;
      RECT  2.505 1.25 2.65 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 5.87 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.045 1.445 0.215 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.655 1.475 0.825 1.75 ;
      RECT  2.225 1.405 2.355 1.75 ;
      RECT  2.745 1.37 2.875 1.75 ;
      RECT  3.245 1.445 3.415 1.75 ;
      RECT  3.79 1.36 3.92 1.75 ;
      RECT  4.3 1.44 4.43 1.75 ;
      RECT  5.52 0.99 5.61 1.75 ;
      RECT  6.02 1.41 6.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  4.455 0.05 4.545 0.215 ;
      RECT  2.455 0.05 2.585 0.345 ;
      RECT  1.195 0.05 1.325 0.36 ;
      RECT  0.675 0.05 0.805 0.39 ;
      RECT  3.485 0.05 3.615 0.39 ;
      RECT  5.5 0.05 5.63 0.39 ;
      RECT  6.02 0.05 6.145 0.39 ;
      RECT  2.975 0.05 3.105 0.42 ;
      RECT  4.375 0.215 4.545 0.305 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.64 0.14 5.405 0.23 ;
      RECT  4.64 0.23 4.73 0.395 ;
      RECT  5.315 0.23 5.405 0.61 ;
      RECT  4.455 0.395 4.73 0.485 ;
      RECT  4.455 0.485 4.545 0.6 ;
      RECT  4.155 0.52 4.245 0.6 ;
      RECT  4.155 0.6 4.545 0.69 ;
      RECT  4.45 0.69 4.545 0.745 ;
      RECT  4.45 0.745 4.58 0.825 ;
      RECT  4.375 0.825 4.58 0.915 ;
      RECT  4.375 0.915 4.465 1.26 ;
      RECT  4.06 1.26 4.62 1.35 ;
      RECT  4.53 1.35 4.62 1.47 ;
      RECT  4.06 1.35 4.15 1.5 ;
      RECT  4.53 1.47 4.94 1.57 ;
      RECT  1.445 0.14 1.615 0.25 ;
      RECT  1.445 0.25 1.545 0.49 ;
      RECT  2.215 0.175 2.305 0.285 ;
      RECT  2.145 0.285 2.305 0.375 ;
      RECT  2.145 0.375 2.235 0.71 ;
      RECT  2.135 0.71 2.235 0.89 ;
      RECT  2.145 0.89 2.235 1.18 ;
      RECT  1.97 1.18 2.235 1.27 ;
      RECT  1.97 1.27 2.09 1.53 ;
      RECT  5.0 0.335 5.205 0.425 ;
      RECT  5.115 0.425 5.205 0.73 ;
      RECT  5.115 0.73 5.66 0.82 ;
      RECT  5.57 0.82 5.66 0.9 ;
      RECT  5.115 0.82 5.205 0.99 ;
      RECT  5.05 0.99 5.205 1.16 ;
      RECT  1.94 0.19 2.055 0.43 ;
      RECT  1.94 0.43 2.04 1.09 ;
      RECT  0.955 0.2 1.045 0.47 ;
      RECT  0.955 0.47 1.345 0.56 ;
      RECT  1.245 0.56 1.345 0.91 ;
      RECT  1.245 0.91 1.425 1.09 ;
      RECT  1.245 1.09 1.345 1.355 ;
      RECT  1.15 1.355 1.345 1.475 ;
      RECT  0.085 0.31 0.25 0.49 ;
      RECT  0.085 0.49 0.175 1.25 ;
      RECT  0.085 1.25 1.005 1.355 ;
      RECT  0.915 1.355 1.005 1.565 ;
      RECT  0.915 1.565 1.835 1.655 ;
      RECT  1.72 1.42 1.835 1.565 ;
      RECT  3.245 0.19 3.335 0.575 ;
      RECT  3.245 0.575 3.675 0.665 ;
      RECT  3.58 0.49 3.675 0.575 ;
      RECT  3.245 0.665 3.335 0.78 ;
      RECT  3.02 0.78 3.335 0.87 ;
      RECT  3.02 0.87 3.11 1.58 ;
      RECT  4.635 0.575 4.805 0.665 ;
      RECT  4.675 0.665 4.765 1.06 ;
      RECT  4.555 1.06 4.765 1.08 ;
      RECT  4.555 1.08 4.81 1.17 ;
      RECT  4.72 1.17 4.81 1.29 ;
      RECT  4.72 1.29 5.12 1.38 ;
      RECT  5.03 1.38 5.12 1.43 ;
      RECT  5.03 1.43 5.425 1.52 ;
      RECT  5.335 1.52 5.425 1.6 ;
      RECT  4.895 0.515 5.025 0.77 ;
      RECT  4.855 0.77 5.025 0.9 ;
      RECT  3.965 0.17 4.055 0.795 ;
      RECT  3.965 0.795 4.285 0.885 ;
      RECT  4.195 0.885 4.285 1.06 ;
      RECT  3.55 1.06 4.285 1.15 ;
      RECT  3.55 1.15 3.64 1.59 ;
      RECT  3.775 0.29 3.875 0.855 ;
      RECT  3.695 0.855 3.875 0.96 ;
      RECT  2.545 0.44 2.645 0.95 ;
      RECT  1.515 0.58 1.615 1.08 ;
      RECT  1.705 0.19 1.83 1.205 ;
      RECT  1.46 1.205 1.83 1.295 ;
      RECT  1.46 1.295 1.58 1.47 ;
      RECT  3.2 0.96 3.31 1.355 ;
      LAYER M2 ;
      RECT  0.11 0.35 3.93 0.45 ;
      RECT  1.69 0.55 2.685 0.65 ;
      RECT  1.475 0.75 5.035 0.85 ;
      RECT  1.285 0.95 2.16 1.05 ;
      RECT  2.06 1.05 2.16 1.15 ;
      RECT  2.06 1.15 3.34 1.25 ;
      LAYER V1 ;
      RECT  0.15 0.35 0.25 0.45 ;
      RECT  1.445 0.35 1.545 0.45 ;
      RECT  3.775 0.35 3.875 0.45 ;
      RECT  1.73 0.55 1.83 0.65 ;
      RECT  2.545 0.55 2.645 0.65 ;
      RECT  1.515 0.75 1.615 0.85 ;
      RECT  2.135 0.75 2.235 0.85 ;
      RECT  4.895 0.75 4.995 0.85 ;
      RECT  1.325 0.95 1.425 1.05 ;
      RECT  1.94 0.95 2.04 1.05 ;
      RECT  3.2 1.15 3.3 1.25 ;
  END
END SEN_ADDF_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_D_4
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_D_4
  CLASS CORE ;
  FOREIGN SEN_ADDF_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 0.705 ;
      RECT  0.35 0.705 1.65 0.81 ;
      RECT  0.35 0.81 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  0.95 0.91 2.25 1.0 ;
      RECT  0.95 1.0 1.05 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.91 0.85 8.08 0.94 ;
      RECT  7.91 0.94 8.05 1.29 ;
      RECT  3.63 0.685 3.73 1.15 ;
      LAYER M2 ;
      RECT  3.59 0.95 8.05 1.05 ;
      LAYER V1 ;
      RECT  7.91 0.95 8.01 1.05 ;
      RECT  3.63 0.95 3.73 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.183 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.045 0.36 4.135 0.51 ;
      RECT  4.045 0.51 4.655 0.6 ;
      RECT  4.55 0.6 4.655 1.025 ;
      RECT  3.98 1.025 4.655 1.115 ;
      RECT  4.55 1.115 4.655 1.49 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.42 0.28 8.54 0.43 ;
      RECT  8.42 0.43 9.055 0.52 ;
      RECT  8.945 0.52 9.055 1.11 ;
      RECT  8.41 1.11 9.055 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.45 0.205 1.75 ;
      RECT  0.0 1.75 9.4 1.85 ;
      RECT  0.575 1.47 0.745 1.75 ;
      RECT  1.095 1.485 1.265 1.75 ;
      RECT  1.625 1.485 1.795 1.75 ;
      RECT  3.77 1.24 3.89 1.75 ;
      RECT  4.29 1.205 4.41 1.75 ;
      RECT  4.81 1.19 4.93 1.75 ;
      RECT  5.335 1.44 5.465 1.75 ;
      RECT  5.885 1.215 6.005 1.75 ;
      RECT  6.135 1.215 6.255 1.75 ;
      RECT  6.65 1.44 6.78 1.75 ;
      RECT  7.17 1.44 7.28 1.75 ;
      RECT  8.175 0.99 8.265 1.75 ;
      RECT  8.675 1.41 8.805 1.75 ;
      RECT  9.2 1.21 9.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      RECT  0.835 0.05 1.005 0.325 ;
      RECT  2.08 0.05 2.25 0.335 ;
      RECT  8.655 0.05 8.825 0.34 ;
      RECT  8.155 0.05 8.285 0.36 ;
      RECT  7.195 0.05 7.33 0.38 ;
      RECT  1.395 0.05 1.525 0.39 ;
      RECT  3.765 0.05 3.895 0.39 ;
      RECT  4.285 0.05 4.415 0.39 ;
      RECT  6.7 0.05 6.81 0.39 ;
      RECT  5.335 0.05 5.465 0.43 ;
      RECT  6.13 0.05 6.26 0.43 ;
      RECT  4.81 0.05 4.93 0.59 ;
      RECT  9.2 0.05 9.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.08 0.14 0.705 0.23 ;
      RECT  0.08 0.23 0.2 0.39 ;
      RECT  0.615 0.23 0.705 0.47 ;
      RECT  0.615 0.47 1.235 0.56 ;
      RECT  1.13 0.38 1.235 0.47 ;
      RECT  7.725 0.185 8.05 0.28 ;
      RECT  7.95 0.28 8.05 0.49 ;
      RECT  7.95 0.49 8.12 0.58 ;
      RECT  6.37 0.22 6.61 0.34 ;
      RECT  6.51 0.34 6.61 0.76 ;
      RECT  6.51 0.76 6.935 0.865 ;
      RECT  6.51 0.865 6.61 1.26 ;
      RECT  6.41 1.26 7.46 1.35 ;
      RECT  7.37 1.35 7.46 1.44 ;
      RECT  6.41 1.35 6.5 1.5 ;
      RECT  7.37 1.44 7.63 1.53 ;
      RECT  3.25 0.235 3.355 0.405 ;
      RECT  3.25 0.405 3.35 1.29 ;
      RECT  1.755 0.19 1.845 0.425 ;
      RECT  1.755 0.425 2.47 0.515 ;
      RECT  2.38 0.515 2.47 0.81 ;
      RECT  2.38 0.81 2.72 0.9 ;
      RECT  2.63 0.9 2.72 1.29 ;
      RECT  2.63 1.29 3.35 1.305 ;
      RECT  2.12 1.305 3.35 1.395 ;
      RECT  2.73 0.145 2.83 0.43 ;
      RECT  2.59 0.43 2.83 0.54 ;
      RECT  7.455 0.32 7.575 0.47 ;
      RECT  6.96 0.47 7.575 0.56 ;
      RECT  6.96 0.56 7.155 0.64 ;
      RECT  7.065 0.64 7.155 1.05 ;
      RECT  6.86 1.05 7.155 1.08 ;
      RECT  6.86 1.08 7.64 1.17 ;
      RECT  7.55 1.17 7.64 1.26 ;
      RECT  7.55 1.26 7.81 1.35 ;
      RECT  7.72 1.35 7.81 1.48 ;
      RECT  7.72 1.48 8.08 1.57 ;
      RECT  7.975 1.4 8.08 1.48 ;
      RECT  0.315 0.34 0.495 0.48 ;
      RECT  0.17 0.48 0.495 0.57 ;
      RECT  0.17 0.57 0.26 1.22 ;
      RECT  0.17 1.22 1.005 1.305 ;
      RECT  0.17 1.305 2.03 1.34 ;
      RECT  0.895 1.34 2.03 1.395 ;
      RECT  1.94 1.395 2.03 1.485 ;
      RECT  1.94 1.485 3.42 1.58 ;
      RECT  3.515 0.19 3.605 0.495 ;
      RECT  3.44 0.495 3.605 0.585 ;
      RECT  3.44 0.585 3.54 1.305 ;
      RECT  3.44 1.305 3.615 1.395 ;
      RECT  3.525 1.395 3.615 1.6 ;
      RECT  5.885 0.32 6.005 0.55 ;
      RECT  5.885 0.55 6.395 0.64 ;
      RECT  6.305 0.64 6.395 1.015 ;
      RECT  5.64 1.015 6.395 1.105 ;
      RECT  5.64 1.105 5.73 1.485 ;
      RECT  7.73 0.4 7.82 0.67 ;
      RECT  7.73 0.67 8.42 0.76 ;
      RECT  8.33 0.76 8.835 0.87 ;
      RECT  7.73 0.76 7.82 1.17 ;
      RECT  5.075 0.19 5.165 0.7 ;
      RECT  5.075 0.7 5.575 0.79 ;
      RECT  5.485 0.79 5.575 0.925 ;
      RECT  5.075 0.79 5.165 1.54 ;
      RECT  2.635 0.63 2.91 0.72 ;
      RECT  2.81 0.72 2.91 1.02 ;
      RECT  5.665 0.29 5.765 0.755 ;
      RECT  5.665 0.755 5.885 0.925 ;
      RECT  3.82 0.51 3.92 0.795 ;
      RECT  3.82 0.795 4.44 0.905 ;
      RECT  7.255 0.71 7.64 0.89 ;
      RECT  3.0 0.235 3.1 1.11 ;
      RECT  2.9 1.11 3.1 1.2 ;
      RECT  2.45 0.99 2.54 1.115 ;
      RECT  1.36 1.115 2.54 1.215 ;
      RECT  5.255 0.89 5.355 1.35 ;
      LAYER M2 ;
      RECT  0.315 0.35 5.805 0.45 ;
      RECT  6.47 0.35 8.09 0.45 ;
      RECT  2.96 0.55 3.96 0.65 ;
      RECT  2.77 0.75 7.43 0.85 ;
      RECT  3.21 1.15 5.395 1.25 ;
      LAYER V1 ;
      RECT  0.355 0.35 0.455 0.45 ;
      RECT  2.73 0.35 2.83 0.45 ;
      RECT  5.665 0.35 5.765 0.45 ;
      RECT  6.51 0.35 6.61 0.45 ;
      RECT  7.95 0.35 8.05 0.45 ;
      RECT  3.0 0.55 3.1 0.65 ;
      RECT  3.82 0.55 3.92 0.65 ;
      RECT  2.81 0.75 2.91 0.85 ;
      RECT  3.44 0.75 3.54 0.85 ;
      RECT  7.29 0.75 7.39 0.85 ;
      RECT  3.25 1.15 3.35 1.25 ;
      RECT  5.255 1.15 5.355 1.25 ;
  END
END SEN_ADDF_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_D_6
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_D_6
  CLASS CORE ;
  FOREIGN SEN_ADDF_D_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.745 2.94 0.9 ;
      RECT  0.355 0.74 0.74 0.85 ;
      LAYER M2 ;
      RECT  0.36 0.75 2.74 0.85 ;
      LAYER V1 ;
      RECT  2.6 0.75 2.7 0.85 ;
      RECT  0.4 0.75 0.5 0.85 ;
      RECT  0.6 0.75 0.7 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.309 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.51 ;
      RECT  1.15 0.51 1.45 0.69 ;
      RECT  1.15 0.69 1.245 0.76 ;
      RECT  0.855 0.76 1.245 0.865 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.309 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.635 0.98 10.91 1.085 ;
      RECT  10.635 1.085 10.735 1.39 ;
      RECT  4.4 0.81 4.84 0.92 ;
      RECT  4.4 0.92 4.5 1.35 ;
      LAYER M2 ;
      RECT  4.36 1.15 10.775 1.25 ;
      LAYER V1 ;
      RECT  10.635 1.15 10.735 1.25 ;
      RECT  4.4 1.15 4.5 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2724 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.25 0.19 5.42 0.36 ;
      RECT  5.33 0.36 5.42 0.51 ;
      RECT  5.33 0.51 6.45 0.69 ;
      RECT  6.35 0.69 6.45 1.075 ;
      RECT  5.15 1.075 6.45 1.19 ;
      RECT  5.75 1.19 5.86 1.49 ;
      RECT  6.35 1.19 6.45 1.49 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  11.665 0.475 12.85 0.595 ;
      RECT  12.72 0.595 12.85 1.11 ;
      RECT  11.69 1.11 12.85 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.44 0.19 1.75 ;
      RECT  0.0 1.75 13.2 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  2.37 1.48 2.54 1.75 ;
      RECT  2.91 1.44 3.04 1.75 ;
      RECT  4.45 1.44 4.58 1.75 ;
      RECT  4.97 1.375 5.1 1.75 ;
      RECT  5.49 1.435 5.62 1.75 ;
      RECT  6.01 1.375 6.14 1.75 ;
      RECT  6.55 1.24 6.655 1.75 ;
      RECT  7.055 1.41 7.185 1.75 ;
      RECT  7.575 1.41 7.705 1.75 ;
      RECT  8.095 1.41 8.225 1.75 ;
      RECT  8.63 1.44 8.76 1.75 ;
      RECT  9.13 1.48 9.3 1.75 ;
      RECT  9.65 1.48 9.82 1.75 ;
      RECT  11.43 1.21 11.55 1.75 ;
      RECT  11.945 1.41 12.075 1.75 ;
      RECT  12.465 1.41 12.595 1.75 ;
      RECT  12.99 1.21 13.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 13.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 13.2 0.05 ;
      RECT  0.06 0.05 0.19 0.36 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.34 0.05 1.465 0.36 ;
      RECT  1.87 0.05 2.0 0.36 ;
      RECT  11.945 0.05 12.075 0.38 ;
      RECT  12.465 0.05 12.595 0.38 ;
      RECT  8.63 0.05 8.76 0.385 ;
      RECT  4.97 0.05 5.1 0.39 ;
      RECT  5.51 0.05 5.62 0.39 ;
      RECT  6.01 0.05 6.14 0.39 ;
      RECT  9.15 0.05 9.28 0.39 ;
      RECT  9.67 0.05 9.8 0.39 ;
      RECT  7.315 0.05 7.445 0.41 ;
      RECT  4.455 0.05 4.575 0.59 ;
      RECT  6.54 0.05 6.655 0.59 ;
      RECT  11.43 0.05 11.55 0.59 ;
      RECT  12.99 0.05 13.11 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 13.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.915 0.14 3.53 0.23 ;
      RECT  2.915 0.23 3.035 0.505 ;
      RECT  3.425 0.23 3.53 1.045 ;
      RECT  2.37 0.505 3.035 0.625 ;
      RECT  2.37 0.625 2.46 0.78 ;
      RECT  1.335 0.78 2.46 0.87 ;
      RECT  1.335 0.87 1.425 1.015 ;
      RECT  0.3 1.015 1.425 1.135 ;
      RECT  3.425 1.045 3.83 1.135 ;
      RECT  3.74 1.135 3.83 1.245 ;
      RECT  3.74 1.245 4.12 1.35 ;
      RECT  3.685 0.14 4.31 0.23 ;
      RECT  3.685 0.23 3.805 0.345 ;
      RECT  4.21 0.23 4.31 1.465 ;
      RECT  3.14 1.465 4.31 1.585 ;
      RECT  7.58 0.14 8.28 0.23 ;
      RECT  7.58 0.23 7.7 0.55 ;
      RECT  7.06 0.375 7.18 0.55 ;
      RECT  7.06 0.55 7.7 0.64 ;
      RECT  2.135 0.215 2.8 0.335 ;
      RECT  2.135 0.335 2.255 0.45 ;
      RECT  1.63 0.315 1.72 0.45 ;
      RECT  1.63 0.45 2.255 0.54 ;
      RECT  10.07 0.215 10.78 0.335 ;
      RECT  10.66 0.335 10.78 0.62 ;
      RECT  10.66 0.62 11.3 0.71 ;
      RECT  11.18 0.24 11.3 0.62 ;
      RECT  11.18 0.71 11.3 0.76 ;
      RECT  11.18 0.76 12.61 0.87 ;
      RECT  11.18 0.87 11.3 1.48 ;
      RECT  10.08 1.48 11.3 1.585 ;
      RECT  6.81 0.19 6.925 0.43 ;
      RECT  6.835 0.43 6.925 0.815 ;
      RECT  6.835 0.815 7.5 0.925 ;
      RECT  6.835 0.925 6.925 1.32 ;
      RECT  6.81 1.32 6.925 1.54 ;
      RECT  8.035 0.35 8.24 0.45 ;
      RECT  8.035 0.45 8.125 0.92 ;
      RECT  7.82 0.92 8.125 1.03 ;
      RECT  4.72 0.315 4.83 0.51 ;
      RECT  4.72 0.51 5.05 0.6 ;
      RECT  4.95 0.6 5.05 1.19 ;
      RECT  4.72 1.19 5.05 1.285 ;
      RECT  4.72 1.285 4.835 1.49 ;
      RECT  8.375 0.39 8.495 0.525 ;
      RECT  8.375 0.525 9.245 0.615 ;
      RECT  8.895 0.29 9.015 0.525 ;
      RECT  9.155 0.615 9.245 0.77 ;
      RECT  9.155 0.77 9.75 0.88 ;
      RECT  9.155 0.88 9.245 1.24 ;
      RECT  8.39 1.24 9.245 1.28 ;
      RECT  8.39 1.28 10.545 1.33 ;
      RECT  9.155 1.33 10.545 1.39 ;
      RECT  8.39 1.33 8.495 1.46 ;
      RECT  10.905 0.17 11.04 0.53 ;
      RECT  9.36 0.5 10.535 0.62 ;
      RECT  10.445 0.62 10.535 0.8 ;
      RECT  9.84 0.62 9.93 1.05 ;
      RECT  10.445 0.8 11.09 0.89 ;
      RECT  11.0 0.89 11.09 1.23 ;
      RECT  9.36 1.05 10.11 1.17 ;
      RECT  10.86 1.23 11.09 1.35 ;
      RECT  3.18 0.32 3.285 0.715 ;
      RECT  3.04 0.715 3.285 0.82 ;
      RECT  5.14 0.51 5.24 0.8 ;
      RECT  5.14 0.8 6.16 0.91 ;
      RECT  8.215 0.785 9.04 0.895 ;
      RECT  8.215 0.895 8.305 1.12 ;
      RECT  7.84 0.32 7.945 0.73 ;
      RECT  7.61 0.73 7.945 0.82 ;
      RECT  7.61 0.82 7.71 1.12 ;
      RECT  7.32 1.12 8.305 1.21 ;
      RECT  7.32 1.21 7.44 1.49 ;
      RECT  7.84 1.21 7.96 1.49 ;
      RECT  10.02 0.75 10.355 0.9 ;
      RECT  3.62 0.47 3.72 0.95 ;
      RECT  3.95 0.365 4.05 1.13 ;
      RECT  6.54 0.78 6.745 1.13 ;
      RECT  1.585 1.015 2.83 1.135 ;
      RECT  3.235 0.91 3.335 1.225 ;
      RECT  3.235 1.225 3.6 1.25 ;
      RECT  0.325 0.31 0.445 0.45 ;
      RECT  0.12 0.45 0.965 0.54 ;
      RECT  0.845 0.31 0.965 0.45 ;
      RECT  0.12 0.54 0.21 1.25 ;
      RECT  0.12 1.25 3.6 1.35 ;
      LAYER M2 ;
      RECT  3.39 0.35 8.215 0.45 ;
      RECT  8.87 0.35 11.045 0.45 ;
      RECT  3.14 0.55 5.28 0.65 ;
      RECT  3.58 0.75 10.335 0.85 ;
      RECT  3.195 0.95 6.68 1.05 ;
      LAYER V1 ;
      RECT  3.43 0.35 3.53 0.45 ;
      RECT  8.075 0.35 8.175 0.45 ;
      RECT  8.91 0.35 9.01 0.45 ;
      RECT  10.905 0.35 11.005 0.45 ;
      RECT  3.18 0.55 3.28 0.65 ;
      RECT  4.21 0.55 4.31 0.65 ;
      RECT  5.14 0.55 5.24 0.65 ;
      RECT  3.62 0.75 3.72 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
      RECT  10.06 0.75 10.16 0.85 ;
      RECT  3.235 0.95 3.335 1.05 ;
      RECT  3.95 0.95 4.05 1.05 ;
      RECT  6.54 0.95 6.64 1.05 ;
  END
END SEN_ADDF_D_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_0P5
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_0P5
  CLASS CORE ;
  FOREIGN SEN_ADDF_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.67 3.315 0.84 ;
      RECT  3.15 0.84 3.25 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1275 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.27 0.71 0.545 0.88 ;
      RECT  3.42 0.51 3.56 0.83 ;
      RECT  2.32 0.55 2.67 0.56 ;
      RECT  2.205 0.56 2.67 0.65 ;
      RECT  1.165 0.55 1.62 0.665 ;
      LAYER M2 ;
      RECT  0.35 0.55 3.59 0.65 ;
      RECT  0.35 0.65 0.45 0.75 ;
      RECT  0.27 0.75 0.45 0.85 ;
      LAYER V1 ;
      RECT  0.31 0.75 0.41 0.85 ;
      RECT  3.45 0.55 3.55 0.65 ;
      RECT  2.53 0.55 2.63 0.65 ;
      RECT  1.275 0.55 1.375 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1275 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.055 0.75 ;
      RECT  1.97 0.75 3.055 0.85 ;
      RECT  2.75 0.85 3.055 0.89 ;
      RECT  0.695 0.71 0.885 0.97 ;
      LAYER M2 ;
      RECT  0.705 0.75 2.15 0.85 ;
      LAYER V1 ;
      RECT  2.01 0.75 2.11 0.85 ;
      RECT  0.745 0.75 0.845 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.555 0.265 1.675 0.355 ;
      RECT  1.555 0.355 1.85 0.455 ;
      RECT  1.75 0.455 1.85 1.11 ;
      RECT  1.55 1.11 1.85 1.29 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.83 0.29 3.955 0.46 ;
      RECT  3.855 0.46 3.955 1.11 ;
      RECT  3.75 1.11 3.955 1.29 ;
      RECT  3.75 1.29 3.85 1.49 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.24 0.445 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  1.29 1.17 1.415 1.75 ;
      RECT  1.805 1.39 1.925 1.75 ;
      RECT  2.355 1.18 2.475 1.75 ;
      RECT  3.545 1.18 3.65 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  3.52 0.05 3.69 0.2 ;
      RECT  2.32 0.05 2.49 0.25 ;
      RECT  1.78 0.05 1.95 0.265 ;
      RECT  0.3 0.05 0.47 0.355 ;
      RECT  1.295 0.05 1.415 0.375 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.09 0.25 2.18 0.34 ;
      RECT  2.09 0.34 2.72 0.43 ;
      RECT  2.63 0.25 2.72 0.34 ;
      RECT  0.82 0.24 1.065 0.36 ;
      RECT  0.975 0.36 1.065 0.825 ;
      RECT  0.975 0.825 1.545 0.915 ;
      RECT  0.975 0.915 1.065 1.225 ;
      RECT  0.86 1.225 1.065 1.49 ;
      RECT  2.85 0.33 3.74 0.42 ;
      RECT  3.65 0.42 3.74 0.93 ;
      RECT  3.355 0.93 3.74 1.02 ;
      RECT  3.355 1.02 3.445 1.225 ;
      RECT  2.85 1.075 3.06 1.2 ;
      RECT  2.97 1.2 3.06 1.225 ;
      RECT  2.97 1.225 3.445 1.315 ;
      RECT  0.065 0.26 0.185 0.445 ;
      RECT  0.065 0.445 0.705 0.545 ;
      RECT  0.585 0.25 0.705 0.445 ;
      RECT  2.075 1.0 2.735 1.09 ;
      RECT  2.075 1.09 2.195 1.215 ;
      RECT  2.61 1.09 2.735 1.22 ;
      RECT  0.065 1.06 0.695 1.15 ;
      RECT  0.59 1.15 0.695 1.325 ;
      RECT  0.065 1.15 0.185 1.35 ;
      RECT  2.59 1.31 2.88 1.56 ;
      LAYER M2 ;
      RECT  0.86 1.35 2.73 1.45 ;
      LAYER V1 ;
      RECT  0.9 1.35 1.0 1.45 ;
      RECT  2.59 1.35 2.69 1.45 ;
  END
END SEN_ADDF_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_1
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_1
  CLASS CORE ;
  FOREIGN SEN_ADDF_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.89 0.755 2.99 1.01 ;
      RECT  2.85 1.01 2.99 1.2 ;
      RECT  1.72 0.63 1.82 1.09 ;
      RECT  0.985 0.8 1.085 1.22 ;
      RECT  0.35 0.71 0.65 0.9 ;
      RECT  0.55 0.9 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 3.03 1.05 ;
      LAYER V1 ;
      RECT  2.89 0.95 2.99 1.05 ;
      RECT  1.72 0.95 1.82 1.05 ;
      RECT  0.985 0.95 1.085 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1413 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.1 0.72 3.2 1.29 ;
      RECT  1.23 0.78 1.33 1.29 ;
      RECT  0.15 0.91 0.25 1.11 ;
      RECT  0.15 1.11 0.45 1.29 ;
      LAYER M2 ;
      RECT  0.31 1.15 3.24 1.25 ;
      LAYER V1 ;
      RECT  3.1 1.15 3.2 1.25 ;
      RECT  1.23 1.15 1.33 1.25 ;
      RECT  0.35 1.15 0.45 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1413 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.68 0.52 2.78 0.94 ;
      RECT  1.91 0.69 2.21 0.895 ;
      RECT  0.75 0.7 0.865 1.09 ;
      LAYER M2 ;
      RECT  0.71 0.75 2.82 0.85 ;
      LAYER V1 ;
      RECT  2.68 0.75 2.78 0.85 ;
      RECT  1.91 0.75 2.01 0.85 ;
      RECT  2.11 0.75 2.21 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1086 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.495 0.245 3.65 0.425 ;
      RECT  3.55 0.425 3.65 1.11 ;
      RECT  3.43 1.11 3.65 1.2 ;
    END
    ANTENNADIFFAREA 0.177 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.51 4.14 0.69 ;
      RECT  3.95 0.69 4.05 0.995 ;
      RECT  3.95 0.995 4.145 1.175 ;
      RECT  3.95 1.175 4.05 1.29 ;
    END
    ANTENNADIFFAREA 0.149 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.6 0.48 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  1.31 1.6 1.48 1.75 ;
      RECT  1.875 1.54 1.995 1.75 ;
      RECT  3.18 1.56 3.35 1.75 ;
      RECT  3.74 1.47 3.91 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  1.84 0.05 2.01 0.305 ;
      RECT  0.33 0.05 0.46 0.39 ;
      RECT  1.33 0.05 1.46 0.39 ;
      RECT  3.215 0.05 3.34 0.4 ;
      RECT  3.755 0.05 3.86 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.32 0.16 3.125 0.25 ;
      RECT  3.035 0.25 3.125 0.535 ;
      RECT  2.32 0.25 2.41 1.18 ;
      RECT  3.035 0.535 3.435 0.625 ;
      RECT  3.325 0.625 3.435 0.94 ;
      RECT  0.84 0.3 1.195 0.42 ;
      RECT  1.105 0.42 1.195 0.6 ;
      RECT  1.105 0.6 1.53 0.69 ;
      RECT  1.44 0.69 1.53 1.18 ;
      RECT  1.44 1.18 2.41 1.27 ;
      RECT  1.44 1.27 1.53 1.395 ;
      RECT  0.84 1.395 1.53 1.485 ;
      RECT  2.13 0.35 2.23 0.4 ;
      RECT  1.575 0.4 2.23 0.52 ;
      RECT  0.065 0.22 0.185 0.495 ;
      RECT  0.065 0.495 0.725 0.59 ;
      RECT  0.605 0.22 0.725 0.495 ;
      RECT  3.755 0.71 3.845 1.29 ;
      RECT  3.3 1.29 3.845 1.38 ;
      RECT  2.5 0.36 2.59 1.38 ;
      RECT  2.5 1.38 3.39 1.47 ;
      RECT  1.62 1.36 2.32 1.45 ;
      RECT  1.62 1.45 1.725 1.58 ;
      RECT  0.065 1.41 0.75 1.5 ;
      RECT  0.065 1.5 0.185 1.59 ;
  END
END SEN_ADDF_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_2
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_2
  CLASS CORE ;
  FOREIGN SEN_ADDF_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.13 0.635 2.45 0.725 ;
      RECT  2.35 0.725 2.45 1.07 ;
      RECT  1.13 0.725 1.25 1.245 ;
      RECT  2.35 1.07 4.34 1.16 ;
      RECT  4.25 0.77 4.34 1.07 ;
      RECT  0.515 0.71 0.65 1.245 ;
      RECT  0.515 1.245 1.25 1.335 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2802 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.645 0.96 5.245 1.055 ;
      RECT  5.155 1.055 5.245 1.15 ;
      RECT  4.645 1.055 4.745 1.32 ;
      RECT  1.35 0.835 1.88 0.925 ;
      RECT  1.35 0.925 1.45 1.3 ;
      RECT  0.15 0.7 0.25 1.32 ;
      LAYER M2 ;
      RECT  0.11 1.15 4.785 1.25 ;
      LAYER V1 ;
      RECT  4.645 1.15 4.745 1.25 ;
      RECT  1.35 1.15 1.45 1.25 ;
      RECT  0.15 1.15 0.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2802 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.905 0.75 4.12 0.97 ;
      RECT  2.68 0.7 2.99 0.9 ;
      RECT  0.75 0.705 0.85 1.14 ;
      LAYER M2 ;
      RECT  0.71 0.75 4.085 0.85 ;
      LAYER V1 ;
      RECT  3.945 0.75 4.045 0.85 ;
      RECT  2.68 0.75 2.78 0.85 ;
      RECT  2.885 0.75 2.985 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.216 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 5.95 0.69 ;
      RECT  5.75 0.69 5.85 1.05 ;
      RECT  5.75 1.05 6.0 1.17 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.51 6.655 0.69 ;
      RECT  6.55 0.69 6.655 1.11 ;
      RECT  6.35 1.11 6.655 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.34 1.61 0.51 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.445 1.43 1.575 1.75 ;
      RECT  1.975 1.455 2.105 1.75 ;
      RECT  2.515 1.455 2.645 1.75 ;
      RECT  3.045 1.44 3.175 1.75 ;
      RECT  5.025 1.48 5.195 1.75 ;
      RECT  5.545 1.48 5.715 1.75 ;
      RECT  6.065 1.495 6.235 1.75 ;
      RECT  6.605 1.41 6.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  1.955 0.05 2.125 0.185 ;
      RECT  2.495 0.05 2.665 0.185 ;
      RECT  3.035 0.05 3.205 0.185 ;
      RECT  1.445 0.05 1.575 0.365 ;
      RECT  5.565 0.05 5.705 0.385 ;
      RECT  0.36 0.05 0.49 0.39 ;
      RECT  6.605 0.05 6.735 0.39 ;
      RECT  6.09 0.05 6.21 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.855 0.14 5.455 0.23 ;
      RECT  3.855 0.23 3.945 0.39 ;
      RECT  5.365 0.23 5.455 0.5 ;
      RECT  3.475 0.39 3.945 0.455 ;
      RECT  0.94 0.455 3.945 0.48 ;
      RECT  0.94 0.48 3.565 0.545 ;
      RECT  5.365 0.5 5.64 0.59 ;
      RECT  3.1 0.545 3.19 0.87 ;
      RECT  0.94 0.545 1.04 1.155 ;
      RECT  5.55 0.59 5.64 0.92 ;
      RECT  3.1 0.87 3.745 0.96 ;
      RECT  3.295 0.16 3.76 0.25 ;
      RECT  3.295 0.25 3.385 0.275 ;
      RECT  1.685 0.275 3.385 0.365 ;
      RECT  4.15 0.32 5.065 0.41 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 0.83 0.59 ;
      RECT  5.185 0.38 5.275 0.515 ;
      RECT  4.61 0.515 5.275 0.605 ;
      RECT  6.155 0.795 6.45 0.895 ;
      RECT  6.155 0.895 6.245 1.295 ;
      RECT  3.655 0.57 4.52 0.635 ;
      RECT  3.28 0.635 4.52 0.66 ;
      RECT  3.28 0.66 3.745 0.725 ;
      RECT  4.43 0.66 4.52 0.74 ;
      RECT  4.43 0.74 5.45 0.83 ;
      RECT  5.36 0.83 5.45 1.04 ;
      RECT  4.43 0.83 4.52 1.3 ;
      RECT  5.36 1.04 5.595 1.13 ;
      RECT  5.505 1.13 5.595 1.295 ;
      RECT  5.505 1.295 6.245 1.385 ;
      RECT  3.85 1.3 4.52 1.39 ;
      RECT  3.85 1.39 3.98 1.48 ;
      RECT  3.27 1.48 3.98 1.57 ;
      RECT  4.84 1.24 5.415 1.33 ;
      RECT  5.325 1.33 5.415 1.5 ;
      RECT  1.66 1.25 3.74 1.35 ;
      RECT  3.57 1.35 3.74 1.39 ;
      RECT  0.065 1.43 0.84 1.52 ;
      RECT  0.065 1.52 0.185 1.635 ;
      RECT  4.09 1.48 4.78 1.57 ;
  END
END SEN_ADDF_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_4
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_4
  CLASS CORE ;
  FOREIGN SEN_ADDF_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.77 0.9 ;
      RECT  7.15 0.9 7.25 0.95 ;
      RECT  7.04 0.95 7.25 1.05 ;
      RECT  2.15 0.54 3.5 0.63 ;
      RECT  3.41 0.63 3.5 0.745 ;
      RECT  2.15 0.63 2.25 1.09 ;
      RECT  3.41 0.745 4.765 0.855 ;
      RECT  0.75 0.7 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
      LAYER M2 ;
      RECT  0.91 0.95 7.25 1.05 ;
      LAYER V1 ;
      RECT  7.11 0.95 7.21 1.05 ;
      RECT  2.15 0.95 2.25 1.05 ;
      RECT  0.95 0.95 1.05 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5529 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.35 0.7 8.65 0.89 ;
      RECT  8.55 0.89 8.65 1.0 ;
      RECT  8.55 1.0 8.72 1.09 ;
      RECT  8.62 1.09 8.72 1.31 ;
      RECT  2.945 0.79 3.32 0.89 ;
      RECT  3.225 0.89 3.32 1.025 ;
      RECT  3.225 1.025 3.36 1.125 ;
      RECT  3.26 1.125 3.36 1.305 ;
      RECT  0.15 0.7 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.29 ;
      LAYER M2 ;
      RECT  0.11 1.15 8.76 1.25 ;
      LAYER V1 ;
      RECT  8.62 1.15 8.72 1.25 ;
      RECT  3.26 1.15 3.36 1.25 ;
      RECT  0.15 1.15 0.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5529 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.7 0.74 7.045 0.85 ;
      RECT  6.7 0.85 6.8 1.1 ;
      RECT  5.045 0.7 5.54 0.9 ;
      RECT  1.35 0.7 1.65 0.9 ;
      RECT  1.35 0.9 1.45 1.1 ;
      LAYER M2 ;
      RECT  1.415 0.75 7.045 0.85 ;
      LAYER V1 ;
      RECT  6.87 0.75 6.97 0.85 ;
      RECT  5.235 0.75 5.335 0.85 ;
      RECT  5.435 0.75 5.535 0.85 ;
      RECT  1.455 0.75 1.555 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4245 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.55 0.495 9.65 0.51 ;
      RECT  9.0 0.51 9.65 0.69 ;
      RECT  9.55 0.69 9.65 1.135 ;
      RECT  8.93 1.135 9.65 1.225 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.025 0.51 10.65 0.69 ;
      RECT  10.55 0.69 10.65 1.11 ;
      RECT  10.025 1.11 10.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 11.0 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  2.68 1.59 2.85 1.75 ;
      RECT  3.3 1.59 3.47 1.75 ;
      RECT  3.88 1.435 4.01 1.75 ;
      RECT  4.4 1.435 4.53 1.75 ;
      RECT  4.92 1.435 5.05 1.75 ;
      RECT  5.44 1.435 5.57 1.75 ;
      RECT  8.035 1.615 8.205 1.75 ;
      RECT  8.66 1.615 8.83 1.75 ;
      RECT  9.22 1.495 9.39 1.75 ;
      RECT  9.74 1.495 9.91 1.75 ;
      RECT  10.28 1.435 10.41 1.75 ;
      RECT  10.805 1.21 10.925 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      RECT  5.46 0.05 5.63 0.215 ;
      RECT  2.72 0.05 2.855 0.225 ;
      RECT  3.88 0.05 4.01 0.35 ;
      RECT  4.4 0.05 4.53 0.35 ;
      RECT  4.92 0.05 5.05 0.35 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  8.12 0.05 8.25 0.36 ;
      RECT  8.68 0.05 8.81 0.36 ;
      RECT  10.28 0.05 10.41 0.36 ;
      RECT  9.24 0.05 9.37 0.385 ;
      RECT  3.32 0.05 3.45 0.43 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  9.765 0.05 9.885 0.59 ;
      RECT  10.805 0.05 10.925 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  5.785 0.16 6.425 0.25 ;
      RECT  5.785 0.25 5.905 0.305 ;
      RECT  6.305 0.25 6.425 0.38 ;
      RECT  5.185 0.305 5.905 0.395 ;
      RECT  5.185 0.395 5.305 0.44 ;
      RECT  3.6 0.44 5.305 0.56 ;
      RECT  6.77 0.25 8.01 0.345 ;
      RECT  2.11 0.36 3.19 0.45 ;
      RECT  0.3 0.45 1.76 0.56 ;
      RECT  7.54 0.465 8.56 0.57 ;
      RECT  5.87 0.51 5.97 0.735 ;
      RECT  5.87 0.735 6.38 0.74 ;
      RECT  5.67 0.74 6.38 0.835 ;
      RECT  5.67 0.835 5.765 1.01 ;
      RECT  3.45 1.01 5.765 1.1 ;
      RECT  3.45 1.1 3.54 1.41 ;
      RECT  2.405 1.41 3.54 1.5 ;
      RECT  2.405 1.5 2.525 1.55 ;
      RECT  1.355 0.16 2.6 0.25 ;
      RECT  1.355 0.25 1.475 0.36 ;
      RECT  1.875 0.25 1.995 1.55 ;
      RECT  1.355 1.44 1.475 1.55 ;
      RECT  1.355 1.55 2.525 1.64 ;
      RECT  8.75 0.5 8.85 0.79 ;
      RECT  8.75 0.79 9.44 0.89 ;
      RECT  9.81 0.79 10.44 0.89 ;
      RECT  9.81 0.89 9.9 1.315 ;
      RECT  8.995 1.315 9.9 1.405 ;
      RECT  8.995 1.405 9.085 1.435 ;
      RECT  6.06 0.36 6.15 0.47 ;
      RECT  6.06 0.47 7.26 0.56 ;
      RECT  6.52 0.56 6.61 1.095 ;
      RECT  5.94 1.095 6.61 1.21 ;
      RECT  6.49 1.21 6.61 1.435 ;
      RECT  6.49 1.435 9.085 1.525 ;
      RECT  7.365 1.03 8.0 1.12 ;
      RECT  7.365 1.12 7.455 1.23 ;
      RECT  6.74 1.23 7.455 1.32 ;
      RECT  3.63 1.21 5.83 1.305 ;
      RECT  3.63 1.305 3.745 1.43 ;
      RECT  5.7 1.305 5.83 1.45 ;
      RECT  5.7 1.45 6.4 1.545 ;
      RECT  2.11 1.23 3.17 1.32 ;
      RECT  7.545 1.23 8.53 1.32 ;
      RECT  0.34 1.24 1.775 1.35 ;
      RECT  0.34 1.35 0.445 1.46 ;
      LAYER M2 ;
      RECT  5.83 0.55 8.95 0.65 ;
      LAYER V1 ;
      RECT  5.87 0.55 5.97 0.65 ;
      RECT  8.75 0.55 8.85 0.65 ;
  END
END SEN_ADDF_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_P1_1
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_P1_1
  CLASS CORE ;
  FOREIGN SEN_ADDF_P1_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.265 0.71 1.25 0.8 ;
      RECT  0.265 0.8 0.45 1.09 ;
      RECT  1.14 0.8 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.89 0.885 1.09 ;
      RECT  0.55 1.09 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.93 0.8 5.05 1.18 ;
      RECT  4.38 0.8 4.61 0.91 ;
      RECT  4.38 0.91 4.48 1.095 ;
      RECT  3.335 0.875 3.435 1.49 ;
      LAYER M2 ;
      RECT  3.295 0.95 5.07 1.05 ;
      LAYER V1 ;
      RECT  4.93 0.95 5.03 1.05 ;
      RECT  4.38 0.95 4.48 1.05 ;
      RECT  3.335 0.95 3.435 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0816 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 2.865 0.63 ;
      RECT  2.55 0.63 2.65 1.015 ;
      RECT  2.55 1.015 2.78 1.135 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.31 5.91 0.49 ;
      RECT  5.805 0.49 5.91 1.31 ;
      RECT  5.75 1.31 5.91 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.77 1.18 0.915 1.35 ;
      RECT  0.825 1.35 0.915 1.75 ;
      RECT  0.06 1.4 0.19 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  1.285 1.445 1.415 1.75 ;
      RECT  1.875 1.45 2.005 1.75 ;
      RECT  2.335 1.465 2.505 1.75 ;
      RECT  4.105 1.425 4.235 1.75 ;
      RECT  5.415 1.63 5.585 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  5.295 0.05 5.465 0.17 ;
      RECT  1.93 0.05 2.045 0.225 ;
      RECT  2.415 0.05 2.545 0.23 ;
      RECT  0.06 0.05 0.19 0.36 ;
      RECT  0.605 0.05 0.735 0.36 ;
      RECT  4.03 0.05 4.16 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.885 0.14 1.84 0.23 ;
      RECT  1.75 0.23 1.84 0.32 ;
      RECT  0.885 0.23 0.985 0.45 ;
      RECT  1.75 0.32 3.61 0.41 ;
      RECT  3.49 0.41 3.61 0.5 ;
      RECT  1.94 0.41 2.03 0.79 ;
      RECT  0.085 0.45 0.985 0.57 ;
      RECT  3.49 0.5 3.615 0.68 ;
      RECT  0.085 0.57 0.175 1.2 ;
      RECT  3.525 0.68 3.615 1.42 ;
      RECT  1.94 0.79 2.245 0.9 ;
      RECT  0.085 1.2 0.45 1.3 ;
      RECT  0.35 1.3 0.45 1.465 ;
      RECT  3.525 1.42 3.765 1.54 ;
      RECT  0.35 1.465 0.73 1.585 ;
      RECT  2.945 0.14 3.83 0.23 ;
      RECT  3.705 0.23 3.83 1.185 ;
      RECT  3.705 1.185 4.66 1.275 ;
      RECT  4.57 1.08 4.66 1.185 ;
      RECT  3.855 1.275 3.97 1.63 ;
      RECT  4.82 0.26 5.61 0.35 ;
      RECT  5.52 0.35 5.61 0.575 ;
      RECT  5.52 0.575 5.715 0.665 ;
      RECT  5.625 0.665 5.715 1.015 ;
      RECT  5.52 1.015 5.715 1.105 ;
      RECT  5.52 1.105 5.61 1.45 ;
      RECT  5.11 1.45 5.61 1.54 ;
      RECT  5.11 1.54 5.215 1.64 ;
      RECT  1.34 0.33 1.66 0.44 ;
      RECT  1.56 0.44 1.66 1.155 ;
      RECT  4.565 0.28 4.685 0.44 ;
      RECT  4.565 0.44 5.43 0.53 ;
      RECT  5.34 0.53 5.43 0.755 ;
      RECT  5.34 0.755 5.535 0.925 ;
      RECT  5.34 0.925 5.43 1.27 ;
      RECT  4.93 1.27 5.43 1.36 ;
      RECT  4.93 1.36 5.02 1.56 ;
      RECT  4.68 1.56 5.02 1.66 ;
      RECT  2.13 0.5 2.25 0.58 ;
      RECT  2.13 0.58 2.425 0.67 ;
      RECT  2.335 0.67 2.425 1.04 ;
      RECT  1.755 0.695 1.85 1.04 ;
      RECT  1.755 1.04 2.425 1.16 ;
      RECT  4.31 0.28 4.42 0.62 ;
      RECT  4.31 0.62 5.25 0.71 ;
      RECT  5.15 0.71 5.25 0.94 ;
      RECT  4.75 0.71 4.84 1.365 ;
      RECT  4.325 1.365 4.84 1.47 ;
      RECT  3.155 0.54 3.39 0.66 ;
      RECT  3.155 0.66 3.245 0.915 ;
      RECT  3.105 0.915 3.245 1.095 ;
      RECT  3.135 1.095 3.245 1.595 ;
      RECT  2.955 0.5 3.055 0.75 ;
      RECT  2.89 0.75 3.055 0.84 ;
      RECT  2.89 0.84 2.98 1.265 ;
      RECT  1.11 0.53 1.46 0.62 ;
      RECT  1.36 0.62 1.46 0.75 ;
      RECT  1.36 0.75 1.47 0.92 ;
      RECT  1.36 0.92 1.46 1.235 ;
      RECT  1.005 1.235 1.46 1.265 ;
      RECT  1.005 1.265 2.98 1.355 ;
      RECT  2.86 1.355 2.98 1.6 ;
      RECT  3.96 0.51 4.06 0.8 ;
      RECT  3.96 0.8 4.29 0.905 ;
      LAYER M2 ;
      RECT  1.52 0.55 4.1 0.65 ;
      LAYER V1 ;
      RECT  1.56 0.55 1.66 0.65 ;
      RECT  3.96 0.55 4.06 0.65 ;
  END
END SEN_ADDF_P1_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_P1_2
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_P1_2
  CLASS CORE ;
  FOREIGN SEN_ADDF_P1_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.93 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
      LAYER M2 ;
      RECT  0.31 0.75 2.07 0.85 ;
      LAYER V1 ;
      RECT  1.93 0.75 2.03 0.85 ;
      RECT  0.35 0.75 0.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.42 0.8 7.52 1.025 ;
      RECT  7.42 1.025 7.935 1.115 ;
      RECT  7.835 0.8 7.935 1.025 ;
      RECT  5.425 0.895 5.535 1.28 ;
      LAYER M2 ;
      RECT  5.385 0.95 7.56 1.05 ;
      LAYER V1 ;
      RECT  7.42 0.95 7.52 1.05 ;
      RECT  5.425 0.95 5.525 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.31 4.67 1.145 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.15 0.31 9.26 1.3 ;
    END
    ANTENNADIFFAREA 0.218 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.4 0.45 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  1.34 1.4 1.46 1.75 ;
      RECT  1.85 1.43 1.98 1.75 ;
      RECT  2.38 1.43 2.51 1.75 ;
      RECT  2.995 1.43 3.125 1.75 ;
      RECT  3.595 1.43 3.725 1.75 ;
      RECT  4.205 1.43 4.335 1.75 ;
      RECT  4.82 1.43 4.95 1.75 ;
      RECT  6.35 1.345 6.48 1.75 ;
      RECT  6.91 1.44 7.04 1.75 ;
      RECT  8.385 1.455 8.495 1.75 ;
      RECT  8.895 1.24 9.015 1.75 ;
      RECT  9.415 1.21 9.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  8.01 0.05 8.18 0.17 ;
      RECT  4.86 0.05 4.99 0.225 ;
      RECT  6.435 0.05 6.565 0.26 ;
      RECT  3.78 0.05 3.905 0.365 ;
      RECT  1.62 0.05 1.74 0.38 ;
      RECT  6.965 0.05 7.095 0.38 ;
      RECT  3.335 0.05 3.465 0.39 ;
      RECT  0.58 0.05 0.71 0.4 ;
      RECT  8.89 0.05 9.015 0.4 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.105 0.05 1.225 0.59 ;
      RECT  4.305 0.05 4.425 0.59 ;
      RECT  9.415 0.05 9.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  5.33 0.14 6.285 0.23 ;
      RECT  6.11 0.23 6.285 0.42 ;
      RECT  6.11 0.42 6.2 1.01 ;
      RECT  6.11 1.01 7.15 1.1 ;
      RECT  7.06 0.87 7.15 1.01 ;
      RECT  6.11 1.1 6.2 1.275 ;
      RECT  6.06 1.275 6.2 1.505 ;
      RECT  2.575 0.16 3.2 0.25 ;
      RECT  2.575 0.25 2.68 0.39 ;
      RECT  3.08 0.25 3.2 0.535 ;
      RECT  3.08 0.535 3.77 0.655 ;
      RECT  7.715 0.26 8.8 0.35 ;
      RECT  8.71 0.35 8.8 0.6 ;
      RECT  8.71 0.6 9.06 0.69 ;
      RECT  8.97 0.69 9.06 1.06 ;
      RECT  8.685 1.06 9.06 1.15 ;
      RECT  8.685 1.15 8.775 1.245 ;
      RECT  8.205 1.245 8.775 1.365 ;
      RECT  8.205 1.365 8.295 1.44 ;
      RECT  8.0 1.44 8.295 1.56 ;
      RECT  4.005 0.24 4.215 0.36 ;
      RECT  4.125 0.36 4.215 1.02 ;
      RECT  3.29 0.785 3.68 0.895 ;
      RECT  3.59 0.895 3.68 1.02 ;
      RECT  3.59 1.02 4.215 1.14 ;
      RECT  4.76 0.32 5.755 0.41 ;
      RECT  4.76 0.41 5.26 0.445 ;
      RECT  5.635 0.41 5.755 0.715 ;
      RECT  4.76 0.445 4.85 0.955 ;
      RECT  5.245 0.715 5.755 0.805 ;
      RECT  5.245 0.805 5.335 1.37 ;
      RECT  5.245 1.37 5.395 1.57 ;
      RECT  5.245 1.57 5.91 1.66 ;
      RECT  5.805 1.35 5.91 1.57 ;
      RECT  6.38 0.35 6.575 0.45 ;
      RECT  6.485 0.45 6.575 0.795 ;
      RECT  6.485 0.795 6.86 0.905 ;
      RECT  2.785 0.35 2.965 0.505 ;
      RECT  2.865 0.505 2.965 1.02 ;
      RECT  2.615 1.02 3.5 1.14 ;
      RECT  7.455 0.44 8.595 0.53 ;
      RECT  8.505 0.53 8.595 0.785 ;
      RECT  8.505 0.785 8.88 0.895 ;
      RECT  8.505 0.895 8.595 1.065 ;
      RECT  8.025 1.065 8.595 1.155 ;
      RECT  8.025 1.155 8.115 1.21 ;
      RECT  7.72 1.21 8.115 1.3 ;
      RECT  7.72 1.3 7.84 1.57 ;
      RECT  7.165 1.44 7.285 1.57 ;
      RECT  7.165 1.57 7.84 1.66 ;
      RECT  5.35 0.5 5.52 0.535 ;
      RECT  5.01 0.535 5.52 0.625 ;
      RECT  5.01 0.625 5.13 1.235 ;
      RECT  1.83 0.23 2.485 0.35 ;
      RECT  2.375 0.35 2.485 0.785 ;
      RECT  2.375 0.785 2.775 0.895 ;
      RECT  2.375 0.895 2.485 1.215 ;
      RECT  1.555 1.215 2.485 1.235 ;
      RECT  1.555 1.235 5.13 1.34 ;
      RECT  1.325 0.47 2.26 0.59 ;
      RECT  6.67 0.47 7.365 0.59 ;
      RECT  7.24 0.59 7.365 0.62 ;
      RECT  7.24 0.62 8.15 0.71 ;
      RECT  8.06 0.71 8.15 0.785 ;
      RECT  7.24 0.71 7.33 1.21 ;
      RECT  8.06 0.785 8.415 0.895 ;
      RECT  7.24 1.21 7.57 1.235 ;
      RECT  6.6 1.235 7.57 1.35 ;
      RECT  7.4 1.35 7.57 1.48 ;
      RECT  0.285 0.49 0.965 0.61 ;
      RECT  0.845 0.61 0.965 1.21 ;
      RECT  3.935 0.51 4.035 0.785 ;
      RECT  3.83 0.785 4.035 0.895 ;
      RECT  5.9 0.505 6.02 1.0 ;
      RECT  5.625 1.0 6.02 1.09 ;
      RECT  5.625 1.09 5.715 1.37 ;
      RECT  5.505 1.37 5.715 1.48 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.585 1.3 0.705 1.44 ;
      RECT  0.585 1.44 1.25 1.56 ;
      LAYER M2 ;
      RECT  2.785 0.35 6.56 0.45 ;
      RECT  0.825 0.55 6.04 0.65 ;
      LAYER V1 ;
      RECT  2.825 0.35 2.925 0.45 ;
      RECT  6.42 0.35 6.52 0.45 ;
      RECT  0.865 0.55 0.965 0.65 ;
      RECT  3.935 0.55 4.035 0.65 ;
      RECT  5.9 0.55 6.0 0.65 ;
  END
END SEN_ADDF_P1_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_P1_3
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_P1_3
  CLASS CORE ;
  FOREIGN SEN_ADDF_P1_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 0.89 ;
      RECT  1.95 0.89 2.25 1.09 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 0.775 1.09 ;
      LAYER M2 ;
      RECT  0.435 0.95 2.29 1.05 ;
      LAYER V1 ;
      RECT  1.95 0.95 2.05 1.05 ;
      RECT  2.15 0.95 2.25 1.05 ;
      RECT  0.475 0.95 0.575 1.05 ;
      RECT  0.675 0.95 0.775 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.204 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.71 ;
      RECT  1.15 0.71 1.655 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.204 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.81 7.25 1.29 ;
      RECT  6.065 0.605 6.165 1.09 ;
      LAYER M2 ;
      RECT  6.025 0.95 7.29 1.05 ;
      LAYER V1 ;
      RECT  7.15 0.95 7.25 1.05 ;
      RECT  6.065 0.95 6.165 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1725 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.925 0.31 4.05 0.475 ;
      RECT  3.925 0.475 4.55 0.59 ;
      RECT  4.43 0.315 4.55 0.475 ;
      RECT  3.925 0.59 4.05 1.04 ;
      RECT  3.925 1.04 4.575 1.16 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.11 0.31 8.25 0.51 ;
      RECT  8.11 0.51 8.735 0.6 ;
      RECT  8.615 0.43 8.735 0.51 ;
      RECT  8.55 0.6 8.65 1.11 ;
      RECT  8.065 1.11 8.735 1.29 ;
    END
    ANTENNADIFFAREA 0.397 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.415 0.45 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  1.335 1.58 1.505 1.75 ;
      RECT  2.035 1.58 2.205 1.75 ;
      RECT  2.575 1.58 2.745 1.75 ;
      RECT  3.14 1.455 3.26 1.75 ;
      RECT  3.65 1.455 3.77 1.75 ;
      RECT  4.17 1.455 4.29 1.75 ;
      RECT  6.13 1.415 6.25 1.75 ;
      RECT  7.82 1.23 7.94 1.75 ;
      RECT  8.34 1.43 8.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  1.095 0.05 1.265 0.22 ;
      RECT  0.59 0.05 0.71 0.38 ;
      RECT  1.63 0.05 1.75 0.385 ;
      RECT  4.17 0.05 4.29 0.385 ;
      RECT  7.82 0.05 7.94 0.385 ;
      RECT  8.355 0.05 8.48 0.385 ;
      RECT  6.16 0.05 6.28 0.42 ;
      RECT  0.07 0.05 0.2 0.44 ;
      RECT  3.13 0.05 3.25 0.585 ;
      RECT  3.65 0.05 3.77 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.895 0.18 2.515 0.27 ;
      RECT  2.425 0.27 2.515 0.36 ;
      RECT  1.895 0.27 2.005 0.475 ;
      RECT  1.37 0.31 1.49 0.475 ;
      RECT  1.37 0.475 2.005 0.575 ;
      RECT  5.08 0.19 5.645 0.28 ;
      RECT  5.555 0.28 5.645 0.465 ;
      RECT  5.08 0.28 5.195 1.39 ;
      RECT  5.555 0.465 5.74 0.585 ;
      RECT  5.635 0.585 5.74 1.4 ;
      RECT  4.14 0.75 4.755 0.93 ;
      RECT  4.665 0.93 4.755 1.39 ;
      RECT  4.665 1.39 5.195 1.48 ;
      RECT  6.68 0.18 7.665 0.28 ;
      RECT  6.68 0.28 6.85 0.305 ;
      RECT  7.575 0.28 7.665 1.38 ;
      RECT  7.17 1.38 7.665 1.47 ;
      RECT  6.395 0.215 6.58 0.335 ;
      RECT  6.49 0.335 6.58 0.395 ;
      RECT  6.49 0.395 7.44 0.46 ;
      RECT  6.96 0.37 7.44 0.395 ;
      RECT  6.49 0.46 7.05 0.485 ;
      RECT  6.76 0.485 6.85 1.36 ;
      RECT  6.365 1.36 6.85 1.48 ;
      RECT  6.755 1.48 6.85 1.56 ;
      RECT  6.755 1.56 7.525 1.66 ;
      RECT  2.165 0.36 2.255 0.45 ;
      RECT  2.165 0.45 2.585 0.54 ;
      RECT  2.48 0.54 2.585 0.805 ;
      RECT  2.48 0.805 2.795 1.09 ;
      RECT  2.48 1.09 2.58 1.205 ;
      RECT  1.605 1.205 2.58 1.31 ;
      RECT  4.655 0.34 4.945 0.46 ;
      RECT  4.845 0.46 4.945 1.3 ;
      RECT  2.675 0.315 2.765 0.51 ;
      RECT  2.675 0.51 2.975 0.69 ;
      RECT  2.885 0.69 2.975 1.185 ;
      RECT  7.305 0.55 7.485 0.575 ;
      RECT  6.94 0.575 7.485 0.665 ;
      RECT  6.94 0.665 7.03 1.385 ;
      RECT  3.38 0.315 3.495 0.69 ;
      RECT  3.38 0.69 3.47 0.795 ;
      RECT  3.065 0.795 3.47 0.905 ;
      RECT  3.365 0.905 3.47 1.055 ;
      RECT  3.365 1.055 3.535 1.185 ;
      RECT  7.92 0.51 8.02 0.785 ;
      RECT  7.92 0.785 8.395 0.895 ;
      RECT  6.285 0.51 6.395 0.925 ;
      RECT  3.56 0.78 3.715 0.95 ;
      RECT  3.625 0.95 3.715 1.275 ;
      RECT  2.91 1.275 4.535 1.365 ;
      RECT  2.91 1.365 3.0 1.4 ;
      RECT  4.445 1.365 4.535 1.57 ;
      RECT  0.33 0.21 0.45 0.47 ;
      RECT  0.33 0.47 0.97 0.56 ;
      RECT  0.865 0.21 0.97 0.47 ;
      RECT  0.865 0.56 0.97 1.025 ;
      RECT  0.865 1.025 1.49 1.115 ;
      RECT  1.4 1.115 1.49 1.4 ;
      RECT  0.865 1.115 0.97 1.48 ;
      RECT  1.4 1.4 3.0 1.49 ;
      RECT  4.445 1.57 5.465 1.66 ;
      RECT  5.35 0.45 5.465 1.57 ;
      RECT  6.5 0.82 6.67 0.99 ;
      RECT  6.5 0.99 6.59 1.18 ;
      RECT  5.735 0.14 6.005 0.31 ;
      RECT  5.885 0.31 6.005 0.53 ;
      RECT  5.885 0.53 5.975 1.18 ;
      RECT  5.885 1.18 6.59 1.27 ;
      RECT  5.885 1.27 5.975 1.495 ;
      RECT  5.555 1.495 5.975 1.66 ;
      RECT  0.07 1.18 0.71 1.295 ;
      RECT  0.07 1.295 0.19 1.485 ;
      RECT  0.585 1.295 0.71 1.57 ;
      RECT  0.585 1.57 1.23 1.66 ;
      RECT  1.11 1.315 1.23 1.57 ;
      LAYER M2 ;
      RECT  2.635 0.55 6.425 0.65 ;
      RECT  7.305 0.55 8.06 0.65 ;
      RECT  2.455 0.95 4.985 1.05 ;
      LAYER V1 ;
      RECT  2.675 0.55 2.775 0.65 ;
      RECT  2.875 0.55 2.975 0.65 ;
      RECT  6.285 0.55 6.385 0.65 ;
      RECT  7.345 0.55 7.445 0.65 ;
      RECT  7.92 0.55 8.02 0.65 ;
      RECT  2.495 0.95 2.595 1.05 ;
      RECT  2.695 0.95 2.795 1.05 ;
      RECT  4.845 0.95 4.945 1.05 ;
  END
END SEN_ADDF_P1_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDF_P1_4
#      Description : "Full adder"
#      Equation    : S=(A^B)^CI:CO=(A&B)|(A&CI)|(B&CI)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDF_P1_4
  CLASS CORE ;
  FOREIGN SEN_ADDF_P1_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.605 0.71 4.25 0.89 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
      LAYER M2 ;
      RECT  0.71 0.75 3.745 0.85 ;
      LAYER V1 ;
      RECT  3.605 0.75 3.705 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.79 ;
      RECT  1.55 0.79 3.25 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 ;
  END B
  PIN CI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  13.035 0.71 14.055 0.89 ;
      RECT  13.945 0.89 14.055 1.09 ;
      RECT  10.95 0.685 11.45 0.89 ;
      LAYER M2 ;
      RECT  11.31 0.75 13.215 0.85 ;
      LAYER V1 ;
      RECT  13.075 0.75 13.175 0.85 ;
      RECT  11.35 0.75 11.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.327 ;
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.95 0.31 9.05 0.51 ;
      RECT  8.35 0.51 9.05 0.69 ;
      RECT  8.35 0.69 8.455 1.04 ;
      RECT  8.35 1.04 9.04 1.16 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  15.925 0.475 16.65 0.595 ;
      RECT  16.55 0.595 16.65 1.11 ;
      RECT  15.95 1.11 16.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 17.0 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  2.565 1.465 2.735 1.75 ;
      RECT  3.085 1.465 3.255 1.75 ;
      RECT  3.53 1.465 3.7 1.75 ;
      RECT  4.055 1.465 4.225 1.75 ;
      RECT  4.575 1.465 4.745 1.75 ;
      RECT  5.095 1.465 5.265 1.75 ;
      RECT  5.615 1.465 5.785 1.75 ;
      RECT  6.06 1.465 6.23 1.75 ;
      RECT  6.58 1.465 6.75 1.75 ;
      RECT  7.02 1.465 7.195 1.75 ;
      RECT  7.545 1.465 7.715 1.75 ;
      RECT  8.065 1.465 8.235 1.75 ;
      RECT  8.585 1.465 8.755 1.75 ;
      RECT  9.105 1.465 9.275 1.75 ;
      RECT  11.56 1.48 11.73 1.75 ;
      RECT  12.08 1.48 12.25 1.75 ;
      RECT  12.6 1.48 12.77 1.75 ;
      RECT  14.655 1.4 14.785 1.75 ;
      RECT  15.175 1.4 15.305 1.75 ;
      RECT  15.69 1.2 15.81 1.75 ;
      RECT  16.205 1.4 16.335 1.75 ;
      RECT  16.76 1.21 16.88 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 17.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
      RECT  14.65 1.75 14.75 1.85 ;
      RECT  15.25 1.75 15.35 1.85 ;
      RECT  15.85 1.75 15.95 1.85 ;
      RECT  16.45 1.75 16.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 17.0 0.05 ;
      RECT  5.875 0.05 6.045 0.305 ;
      RECT  6.395 0.05 6.565 0.305 ;
      RECT  11.015 0.05 11.185 0.305 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.1 0.05 1.23 0.385 ;
      RECT  1.62 0.05 1.75 0.385 ;
      RECT  2.14 0.05 2.27 0.385 ;
      RECT  7.505 0.05 7.635 0.385 ;
      RECT  8.605 0.05 8.735 0.385 ;
      RECT  16.205 0.05 16.335 0.385 ;
      RECT  11.58 0.05 11.71 0.39 ;
      RECT  2.585 0.05 2.715 0.4 ;
      RECT  3.105 0.05 3.235 0.4 ;
      RECT  6.985 0.05 7.115 0.4 ;
      RECT  9.235 0.05 9.365 0.4 ;
      RECT  12.1 0.05 12.23 0.4 ;
      RECT  12.62 0.05 12.735 0.4 ;
      RECT  14.655 0.05 14.785 0.4 ;
      RECT  15.175 0.05 15.305 0.4 ;
      RECT  15.685 0.05 15.815 0.4 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  8.06 0.05 8.18 0.59 ;
      RECT  16.75 0.05 16.87 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 17.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
      RECT  14.65 -0.05 14.75 0.05 ;
      RECT  15.25 -0.05 15.35 0.05 ;
      RECT  15.85 -0.05 15.95 0.05 ;
      RECT  16.45 -0.05 16.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.41 0.17 4.52 0.27 ;
      RECT  3.37 0.27 4.52 0.39 ;
      RECT  3.37 0.39 3.49 0.525 ;
      RECT  2.34 0.46 2.45 0.525 ;
      RECT  2.34 0.525 3.49 0.645 ;
      RECT  9.57 0.21 10.78 0.305 ;
      RECT  9.57 0.305 10.21 0.32 ;
      RECT  9.57 0.32 9.69 0.505 ;
      RECT  10.09 0.32 10.21 0.61 ;
      RECT  9.14 0.505 9.69 0.605 ;
      RECT  9.14 0.605 9.24 0.785 ;
      RECT  10.09 0.61 10.435 0.7 ;
      RECT  10.315 0.7 10.435 1.48 ;
      RECT  8.545 0.785 9.24 0.895 ;
      RECT  9.715 1.48 10.995 1.6 ;
      RECT  4.61 0.24 5.76 0.36 ;
      RECT  5.64 0.36 5.76 0.395 ;
      RECT  4.61 0.36 4.72 0.66 ;
      RECT  5.64 0.395 6.8 0.515 ;
      RECT  6.68 0.185 6.8 0.395 ;
      RECT  12.825 0.24 13.5 0.36 ;
      RECT  12.825 0.36 12.93 0.54 ;
      RECT  11.845 0.4 11.965 0.54 ;
      RECT  11.845 0.54 12.93 0.66 ;
      RECT  12.81 0.66 12.93 1.06 ;
      RECT  11.79 1.06 13.455 1.18 ;
      RECT  13.335 1.18 13.455 1.32 ;
      RECT  13.8 0.24 14.52 0.36 ;
      RECT  14.41 0.36 14.52 0.505 ;
      RECT  14.41 0.505 15.585 0.625 ;
      RECT  15.48 0.625 15.585 1.165 ;
      RECT  14.41 0.625 14.52 1.465 ;
      RECT  14.87 1.165 15.585 1.285 ;
      RECT  13.9 1.465 14.52 1.585 ;
      RECT  10.75 0.395 11.485 0.5 ;
      RECT  10.75 0.5 10.85 1.085 ;
      RECT  10.75 1.085 11.445 1.175 ;
      RECT  10.99 1.08 11.16 1.085 ;
      RECT  11.325 1.175 11.445 1.27 ;
      RECT  11.325 1.27 12.975 1.39 ;
      RECT  10.31 0.405 10.66 0.52 ;
      RECT  10.55 0.52 10.66 1.27 ;
      RECT  10.55 1.27 11.215 1.39 ;
      RECT  11.095 1.39 11.215 1.48 ;
      RECT  13.03 0.455 14.32 0.575 ;
      RECT  14.22 0.575 14.32 1.185 ;
      RECT  13.655 1.185 14.32 1.305 ;
      RECT  13.655 1.305 13.775 1.44 ;
      RECT  13.05 1.44 13.775 1.56 ;
      RECT  4.835 0.465 5.525 0.585 ;
      RECT  5.435 0.585 5.525 1.05 ;
      RECT  4.81 1.05 6.985 1.17 ;
      RECT  6.88 0.91 6.985 1.05 ;
      RECT  7.25 0.475 7.93 0.595 ;
      RECT  7.25 0.595 7.37 0.605 ;
      RECT  6.555 0.605 7.37 0.695 ;
      RECT  6.555 0.695 6.645 0.78 ;
      RECT  7.25 0.695 7.37 1.05 ;
      RECT  6.085 0.78 6.645 0.895 ;
      RECT  7.25 1.05 7.985 1.17 ;
      RECT  3.59 0.5 4.51 0.62 ;
      RECT  4.41 0.62 4.51 0.75 ;
      RECT  4.41 0.75 5.34 0.895 ;
      RECT  4.41 0.895 4.51 1.05 ;
      RECT  2.28 1.05 4.51 1.17 ;
      RECT  9.83 0.41 9.94 0.75 ;
      RECT  9.33 0.75 9.94 0.85 ;
      RECT  9.83 0.85 9.94 1.27 ;
      RECT  9.44 1.27 10.18 1.39 ;
      RECT  15.675 0.51 15.775 0.785 ;
      RECT  15.675 0.785 16.44 0.895 ;
      RECT  11.595 0.79 12.405 0.89 ;
      RECT  11.595 0.89 11.695 1.09 ;
      RECT  7.475 0.795 8.185 0.895 ;
      RECT  8.095 0.895 8.185 1.26 ;
      RECT  0.285 0.475 2.045 0.595 ;
      RECT  1.34 0.595 1.43 1.26 ;
      RECT  1.34 1.26 8.185 1.285 ;
      RECT  1.34 1.285 9.25 1.375 ;
      RECT  9.15 1.09 9.25 1.285 ;
      RECT  14.61 0.78 15.23 0.9 ;
      RECT  14.61 0.9 14.71 1.29 ;
      RECT  10.03 0.79 10.145 1.18 ;
      RECT  0.065 1.205 1.225 1.325 ;
      RECT  0.065 1.325 0.185 1.43 ;
      RECT  1.105 1.325 1.225 1.465 ;
      RECT  1.105 1.465 2.32 1.585 ;
      LAYER M2 ;
      RECT  14.18 0.55 15.815 0.65 ;
      RECT  5.16 0.75 9.51 0.85 ;
      RECT  9.75 0.75 11.145 0.85 ;
      RECT  9.75 0.85 9.85 0.95 ;
      RECT  11.045 0.85 11.145 0.95 ;
      RECT  6.845 0.95 9.85 1.05 ;
      RECT  11.045 0.95 11.735 1.05 ;
      RECT  9.995 0.95 10.89 1.05 ;
      RECT  9.11 1.15 10.69 1.25 ;
      RECT  13.305 1.15 14.75 1.25 ;
      LAYER V1 ;
      RECT  14.22 0.55 14.32 0.65 ;
      RECT  15.675 0.55 15.775 0.65 ;
      RECT  5.2 0.75 5.3 0.85 ;
      RECT  9.37 0.75 9.47 0.85 ;
      RECT  6.885 0.95 6.985 1.05 ;
      RECT  10.035 0.95 10.135 1.05 ;
      RECT  10.75 0.95 10.85 1.05 ;
      RECT  11.595 0.95 11.695 1.05 ;
      RECT  9.15 1.15 9.25 1.25 ;
      RECT  10.55 1.15 10.65 1.25 ;
      RECT  13.345 1.15 13.445 1.25 ;
      RECT  14.61 1.15 14.71 1.25 ;
  END
END SEN_ADDF_P1_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_0P5
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_0P5
  CLASS CORE ;
  FOREIGN SEN_ADDH_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 0.85 ;
      RECT  0.905 0.85 1.85 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0684 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.84 0.685 1.08 ;
      RECT  0.55 1.08 2.05 1.17 ;
      RECT  1.95 0.65 2.05 1.08 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0684 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.425 0.21 2.525 0.91 ;
      RECT  2.35 0.91 2.525 1.52 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.12 0.21 0.25 1.53 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.44 0.49 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.14 1.44 1.27 1.75 ;
      RECT  1.63 1.33 1.76 1.75 ;
      RECT  2.15 1.44 2.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.87 0.05 1.0 0.28 ;
      RECT  2.15 0.05 2.28 0.38 ;
      RECT  0.36 0.05 0.49 0.44 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.275 0.17 1.695 0.215 ;
      RECT  1.275 0.215 2.06 0.28 ;
      RECT  1.58 0.28 2.06 0.335 ;
      RECT  1.97 0.335 2.06 0.47 ;
      RECT  1.97 0.47 2.335 0.56 ;
      RECT  2.15 0.56 2.335 0.715 ;
      RECT  2.15 0.715 2.24 1.26 ;
      RECT  1.895 1.26 2.24 1.35 ;
      RECT  1.895 1.35 2.015 1.57 ;
      RECT  0.625 0.24 0.745 0.37 ;
      RECT  0.625 0.37 1.25 0.485 ;
      RECT  1.16 0.485 1.25 0.54 ;
      RECT  1.42 0.43 1.51 0.63 ;
      RECT  0.34 0.63 1.51 0.72 ;
      RECT  0.34 0.72 0.43 1.26 ;
      RECT  0.34 1.26 1.525 1.35 ;
      RECT  1.405 1.35 1.525 1.51 ;
      RECT  0.865 1.35 0.985 1.61 ;
  END
END SEN_ADDH_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_1
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_1
  CLASS CORE ;
  FOREIGN SEN_ADDH_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 1.65 0.9 ;
      LAYER M2 ;
      RECT  1.1 0.75 1.7 0.85 ;
      LAYER V1 ;
      RECT  1.25 0.75 1.35 0.85 ;
      RECT  1.45 0.75 1.55 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0792 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.66 1.01 ;
      RECT  0.55 1.01 1.85 1.1 ;
      RECT  1.75 0.9 1.85 1.01 ;
      RECT  0.55 1.1 0.66 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0792 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.305 2.53 0.49 ;
      RECT  2.35 0.49 2.45 1.31 ;
      RECT  2.35 1.31 2.53 1.49 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.31 0.25 0.49 ;
      RECT  0.15 0.49 0.25 1.31 ;
      RECT  0.065 1.31 0.25 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.355 1.61 0.525 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.355 1.61 1.525 1.75 ;
      RECT  2.06 1.61 2.23 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.865 0.05 0.995 0.39 ;
      RECT  2.12 0.05 2.25 0.39 ;
      RECT  0.34 0.05 0.46 0.57 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.55 0.225 2.03 0.345 ;
      RECT  1.94 0.345 2.03 0.5 ;
      RECT  1.94 0.5 2.26 0.59 ;
      RECT  2.16 0.59 2.26 1.41 ;
      RECT  1.175 1.41 2.26 1.5 ;
      RECT  1.175 1.5 1.265 1.545 ;
      RECT  1.065 1.545 1.265 1.65 ;
      RECT  0.61 0.35 0.73 0.51 ;
      RECT  0.61 0.51 1.22 0.6 ;
      RECT  1.095 0.39 1.22 0.51 ;
      RECT  1.33 0.46 1.85 0.55 ;
      RECT  1.75 0.55 1.85 0.7 ;
      RECT  1.75 0.7 2.05 0.79 ;
      RECT  1.95 0.79 2.05 1.21 ;
      RECT  0.87 1.21 2.05 1.3 ;
      RECT  0.87 1.3 0.96 1.41 ;
      RECT  0.34 0.725 0.43 1.41 ;
      RECT  0.34 1.41 0.96 1.5 ;
  END
END SEN_ADDH_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_2
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_2
  CLASS CORE ;
  FOREIGN SEN_ADDH_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.45 0.82 ;
      RECT  1.55 0.82 3.0 0.89 ;
      RECT  2.35 0.89 3.0 0.92 ;
      LAYER M2 ;
      RECT  1.9 0.75 2.5 0.85 ;
      LAYER V1 ;
      RECT  2.05 0.75 2.15 0.85 ;
      RECT  2.25 0.75 2.35 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.156 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.82 3.525 0.92 ;
      RECT  3.15 0.92 3.25 1.075 ;
      RECT  0.95 0.71 1.05 0.91 ;
      RECT  0.95 0.91 1.45 1.0 ;
      RECT  0.95 1.0 2.25 1.075 ;
      RECT  0.95 1.075 3.25 1.1 ;
      RECT  2.15 1.1 3.25 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.156 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.145 0.5 4.25 1.5 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.31 0.31 0.45 0.49 ;
      RECT  0.35 0.49 0.45 1.31 ;
      RECT  0.31 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.09 1.61 1.26 1.75 ;
      RECT  2.165 1.53 2.295 1.75 ;
      RECT  2.73 1.63 2.9 1.75 ;
      RECT  3.38 1.63 3.55 1.75 ;
      RECT  3.8 1.63 3.97 1.75 ;
      RECT  4.415 1.21 4.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  3.335 0.05 3.505 0.185 ;
      RECT  1.08 0.05 1.25 0.305 ;
      RECT  1.62 0.05 1.745 0.36 ;
      RECT  3.875 0.05 4.005 0.365 ;
      RECT  0.585 0.05 0.705 0.545 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  4.415 0.05 4.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.835 0.16 2.455 0.25 ;
      RECT  2.34 0.25 2.455 0.425 ;
      RECT  1.835 0.25 1.94 0.505 ;
      RECT  0.795 0.4 1.51 0.505 ;
      RECT  0.795 0.505 1.94 0.52 ;
      RECT  1.42 0.52 1.94 0.595 ;
      RECT  2.545 0.275 3.785 0.365 ;
      RECT  2.08 0.36 2.2 0.515 ;
      RECT  2.08 0.515 2.65 0.605 ;
      RECT  2.55 0.605 2.65 0.64 ;
      RECT  2.55 0.64 3.8 0.73 ;
      RECT  3.71 0.73 3.8 1.255 ;
      RECT  0.54 0.73 0.63 1.21 ;
      RECT  0.54 1.21 2.025 1.255 ;
      RECT  0.54 1.255 3.8 1.3 ;
      RECT  1.86 1.3 3.8 1.345 ;
      RECT  2.78 0.455 4.045 0.545 ;
      RECT  3.955 0.545 4.045 1.45 ;
      RECT  2.51 1.45 4.045 1.54 ;
      RECT  2.51 1.54 2.6 1.55 ;
      RECT  2.385 1.55 2.6 1.64 ;
      RECT  0.8 1.41 1.77 1.5 ;
  END
END SEN_ADDH_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_4
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_4
  CLASS CORE ;
  FOREIGN SEN_ADDH_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 3.45 0.82 ;
      RECT  2.35 0.82 4.435 0.89 ;
      RECT  3.35 0.89 4.435 0.915 ;
      LAYER M2 ;
      RECT  2.9 0.75 3.5 0.85 ;
      LAYER V1 ;
      RECT  3.05 0.75 3.15 0.85 ;
      RECT  3.25 0.75 3.35 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3114 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.82 5.25 0.92 ;
      RECT  4.75 0.92 4.85 1.09 ;
      RECT  1.35 0.71 1.45 0.9 ;
      RECT  1.35 0.9 2.25 1.0 ;
      RECT  1.35 1.0 3.25 1.09 ;
      RECT  3.15 1.09 4.85 1.18 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3114 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.835 0.51 6.45 0.69 ;
      RECT  6.35 0.69 6.45 1.1 ;
      RECT  5.835 1.1 6.45 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.97 0.69 ;
      RECT  0.35 0.69 0.45 1.11 ;
      RECT  0.35 1.11 0.97 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  0.595 1.43 0.725 1.75 ;
      RECT  1.175 1.415 1.305 1.75 ;
      RECT  1.815 1.6 1.985 1.75 ;
      RECT  3.385 1.505 3.515 1.75 ;
      RECT  4.035 1.63 4.205 1.75 ;
      RECT  4.705 1.63 4.875 1.75 ;
      RECT  5.42 1.63 5.59 1.75 ;
      RECT  6.075 1.425 6.205 1.75 ;
      RECT  6.615 1.21 6.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  5.005 0.05 5.175 0.185 ;
      RECT  1.635 0.05 1.765 0.345 ;
      RECT  2.155 0.05 2.285 0.345 ;
      RECT  5.555 0.05 5.685 0.365 ;
      RECT  2.675 0.05 2.81 0.37 ;
      RECT  0.595 0.05 0.725 0.39 ;
      RECT  6.075 0.05 6.205 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.12 0.05 1.24 0.59 ;
      RECT  6.615 0.05 6.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.94 0.2 3.64 0.32 ;
      RECT  2.94 0.32 3.06 0.5 ;
      RECT  1.35 0.44 2.565 0.5 ;
      RECT  1.35 0.5 3.06 0.56 ;
      RECT  2.475 0.56 3.06 0.59 ;
      RECT  4.215 0.275 5.445 0.365 ;
      RECT  3.98 0.32 4.1 0.455 ;
      RECT  3.98 0.455 5.74 0.545 ;
      RECT  5.65 0.545 5.74 0.785 ;
      RECT  5.65 0.785 6.235 0.895 ;
      RECT  5.65 0.895 5.74 1.45 ;
      RECT  3.8 1.45 5.74 1.54 ;
      RECT  3.8 1.54 3.895 1.55 ;
      RECT  3.665 1.55 3.895 1.64 ;
      RECT  3.175 0.44 3.87 0.56 ;
      RECT  3.78 0.56 3.87 0.64 ;
      RECT  3.78 0.64 5.46 0.73 ;
      RECT  5.36 0.73 5.46 1.27 ;
      RECT  0.55 0.79 1.15 0.89 ;
      RECT  1.06 0.89 1.15 1.2 ;
      RECT  1.06 1.2 3.04 1.27 ;
      RECT  1.06 1.27 5.46 1.29 ;
      RECT  2.905 1.29 5.46 1.36 ;
      RECT  1.45 1.4 2.82 1.49 ;
  END
END SEN_ADDH_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_D_1
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_D_1
  CLASS CORE ;
  FOREIGN SEN_ADDH_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.77 0.71 1.305 0.915 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0921 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.11 0.51 2.25 0.89 ;
      RECT  2.11 0.89 2.2 1.26 ;
      RECT  0.95 1.26 2.2 1.35 ;
      RECT  0.95 1.35 1.25 1.49 ;
      RECT  2.11 1.35 2.2 1.57 ;
      RECT  2.11 1.57 3.155 1.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1059 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.63 0.19 1.735 0.455 ;
      RECT  1.63 0.455 1.85 0.545 ;
      RECT  1.75 0.545 1.85 0.99 ;
      RECT  1.63 0.99 1.85 1.09 ;
      RECT  1.63 1.09 1.735 1.16 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.37 0.14 3.05 0.24 ;
      RECT  2.925 0.24 3.05 0.8 ;
      RECT  2.795 0.8 3.05 0.89 ;
      RECT  2.795 0.89 2.885 1.35 ;
      RECT  2.3 1.29 2.405 1.35 ;
      RECT  2.3 1.35 2.97 1.46 ;
    END
    ANTENNADIFFAREA 0.234 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.77 1.03 0.98 1.15 ;
      RECT  0.77 1.15 0.86 1.75 ;
      RECT  0.065 1.435 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  1.365 1.44 1.485 1.75 ;
      RECT  1.875 1.44 1.995 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.85 0.05 0.94 0.36 ;
      RECT  1.875 0.05 1.995 0.36 ;
      RECT  0.335 0.05 0.435 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.16 0.19 2.25 0.33 ;
      RECT  2.16 0.33 2.445 0.42 ;
      RECT  2.355 0.42 2.445 0.78 ;
      RECT  2.355 0.78 2.495 0.95 ;
      RECT  2.355 0.95 2.445 1.0 ;
      RECT  2.29 1.0 2.445 1.17 ;
      RECT  1.38 0.21 1.535 0.38 ;
      RECT  1.445 0.38 1.535 0.77 ;
      RECT  1.445 0.77 1.615 0.86 ;
      RECT  1.445 0.86 1.535 1.04 ;
      RECT  1.07 1.04 1.535 1.16 ;
      RECT  2.615 0.35 2.81 0.465 ;
      RECT  2.615 0.465 2.705 1.04 ;
      RECT  2.57 1.04 2.705 1.21 ;
      RECT  0.58 0.305 0.68 0.785 ;
      RECT  0.275 0.785 0.68 0.895 ;
      RECT  0.575 0.895 0.68 1.415 ;
      RECT  3.185 0.36 3.305 1.13 ;
      RECT  3.045 1.13 3.305 1.25 ;
      RECT  0.065 0.315 0.185 1.15 ;
      RECT  0.065 1.15 0.445 1.25 ;
      RECT  0.325 1.25 0.445 1.33 ;
      LAYER M2 ;
      RECT  0.54 0.35 2.81 0.45 ;
      RECT  0.215 1.15 3.295 1.25 ;
      LAYER V1 ;
      RECT  0.58 0.35 0.68 0.45 ;
      RECT  2.67 0.35 2.77 0.45 ;
      RECT  0.255 1.15 0.355 1.25 ;
      RECT  3.155 1.15 3.255 1.25 ;
  END
END SEN_ADDH_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_D_2
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_D_2
  CLASS CORE ;
  FOREIGN SEN_ADDH_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.935 0.71 1.71 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1845 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.495 0.51 2.595 0.71 ;
      RECT  2.35 0.71 2.595 0.91 ;
      RECT  2.35 0.91 2.45 1.26 ;
      RECT  1.35 1.26 2.795 1.35 ;
      RECT  1.35 1.35 1.45 1.485 ;
      RECT  2.695 1.35 2.795 1.57 ;
      RECT  1.285 1.485 1.45 1.655 ;
      RECT  2.695 1.57 4.135 1.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2034 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.1 0.51 2.26 0.69 ;
      RECT  2.15 0.69 2.26 0.99 ;
      RECT  2.1 0.99 2.26 1.16 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.23 4.34 0.32 ;
      RECT  3.75 0.32 3.85 0.415 ;
      RECT  3.115 0.415 3.85 0.52 ;
      RECT  3.75 0.52 3.85 1.37 ;
      RECT  3.75 1.37 4.345 1.38 ;
      RECT  4.225 1.29 4.345 1.37 ;
      RECT  3.14 1.23 3.26 1.38 ;
      RECT  3.14 1.38 4.345 1.47 ;
    END
    ANTENNADIFFAREA 0.428 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.105 1.24 1.22 1.41 ;
      RECT  1.105 1.41 1.195 1.75 ;
      RECT  0.075 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.595 1.24 0.715 1.75 ;
      RECT  1.73 1.44 1.85 1.75 ;
      RECT  2.36 1.44 2.475 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.595 0.05 0.715 0.36 ;
      RECT  1.115 0.05 1.235 0.36 ;
      RECT  1.84 0.05 1.96 0.36 ;
      RECT  2.36 0.05 2.48 0.36 ;
      RECT  0.075 0.05 0.185 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.88 0.19 3.545 0.325 ;
      RECT  2.88 0.325 2.995 0.635 ;
      RECT  2.88 0.635 3.59 0.725 ;
      RECT  3.5 0.725 3.59 1.05 ;
      RECT  2.895 1.05 3.59 1.14 ;
      RECT  3.375 1.14 3.59 1.225 ;
      RECT  2.895 1.14 3.0 1.335 ;
      RECT  2.645 0.19 2.775 0.36 ;
      RECT  2.685 0.36 2.775 0.815 ;
      RECT  2.685 0.815 3.39 0.925 ;
      RECT  2.685 0.925 2.775 1.0 ;
      RECT  2.645 1.0 2.775 1.17 ;
      RECT  1.345 0.31 1.455 0.45 ;
      RECT  0.655 0.45 1.455 0.57 ;
      RECT  0.655 0.57 0.745 0.785 ;
      RECT  0.455 0.785 0.745 0.895 ;
      RECT  0.655 0.895 0.745 1.0 ;
      RECT  0.655 1.0 0.975 1.09 ;
      RECT  0.855 1.09 0.975 1.17 ;
      RECT  0.275 0.45 0.48 0.57 ;
      RECT  0.275 0.57 0.365 1.14 ;
      RECT  0.275 1.14 0.49 1.26 ;
      RECT  1.61 0.5 2.005 0.62 ;
      RECT  1.915 0.62 2.005 1.015 ;
      RECT  1.35 1.015 2.005 1.135 ;
      RECT  3.94 0.41 4.055 1.065 ;
      RECT  3.94 1.065 4.125 1.25 ;
      LAYER M2 ;
      RECT  1.31 0.35 3.035 0.45 ;
      RECT  0.31 1.15 4.125 1.25 ;
      LAYER V1 ;
      RECT  1.35 0.35 1.45 0.45 ;
      RECT  2.895 0.35 2.995 0.45 ;
      RECT  0.35 1.15 0.45 1.25 ;
      RECT  3.985 1.15 4.085 1.25 ;
  END
END SEN_ADDH_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_D_3
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_D_3
  CLASS CORE ;
  FOREIGN SEN_ADDH_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.71 ;
      RECT  1.15 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.276 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.935 0.51 4.05 0.73 ;
      RECT  3.935 0.73 4.11 0.9 ;
      RECT  3.935 0.9 4.045 1.275 ;
      RECT  2.735 0.91 2.845 1.215 ;
      RECT  2.735 1.215 3.25 1.275 ;
      RECT  2.735 1.275 4.25 1.305 ;
      RECT  3.15 1.305 4.25 1.365 ;
      RECT  3.15 1.365 3.25 1.49 ;
      RECT  4.15 1.365 4.25 1.57 ;
      RECT  4.15 1.57 6.2 1.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3042 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.125 0.3 3.25 0.47 ;
      RECT  3.125 0.47 3.8 0.595 ;
      RECT  3.55 0.595 3.65 1.0 ;
      RECT  3.075 1.0 3.83 1.125 ;
    END
    ANTENNADIFFAREA 0.369 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.185 6.52 0.305 ;
      RECT  4.35 0.305 5.45 0.315 ;
      RECT  6.43 0.305 6.52 0.36 ;
      RECT  4.35 0.315 4.44 0.36 ;
      RECT  5.345 0.315 5.45 1.35 ;
      RECT  4.69 1.35 6.52 1.46 ;
      RECT  6.43 1.22 6.52 1.35 ;
    END
    ANTENNADIFFAREA 0.623 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.36 1.41 1.49 1.75 ;
      RECT  2.13 1.395 2.26 1.75 ;
      RECT  2.66 1.575 2.79 1.75 ;
      RECT  3.37 1.455 3.54 1.75 ;
      RECT  3.89 1.455 4.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  0.84 0.05 0.97 0.36 ;
      RECT  1.36 0.05 1.49 0.36 ;
      RECT  3.885 0.05 4.015 0.36 ;
      RECT  3.365 0.05 3.495 0.38 ;
      RECT  2.68 0.05 2.8 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.82 0.2 2.54 0.32 ;
      RECT  6.13 0.415 6.3 0.45 ;
      RECT  5.61 0.45 6.3 0.56 ;
      RECT  5.61 0.56 5.7 1.145 ;
      RECT  5.61 1.145 6.3 1.255 ;
      RECT  4.54 0.405 5.235 0.525 ;
      RECT  5.13 0.525 5.235 1.14 ;
      RECT  4.48 1.14 5.235 1.26 ;
      RECT  4.48 1.26 4.6 1.42 ;
      RECT  4.16 0.465 4.26 0.54 ;
      RECT  4.16 0.54 4.365 0.635 ;
      RECT  4.275 0.635 4.365 0.83 ;
      RECT  4.275 0.83 4.99 0.94 ;
      RECT  4.275 0.94 4.365 1.015 ;
      RECT  4.19 1.015 4.365 1.185 ;
      RECT  0.065 0.46 0.73 0.585 ;
      RECT  0.065 0.585 0.185 1.145 ;
      RECT  0.065 1.145 0.735 1.265 ;
      RECT  0.825 0.475 1.77 0.595 ;
      RECT  0.825 0.595 0.925 0.785 ;
      RECT  0.3 0.785 0.925 0.895 ;
      RECT  0.825 0.895 0.925 1.075 ;
      RECT  0.825 1.075 1.74 1.195 ;
      RECT  1.63 1.195 1.74 1.38 ;
      RECT  2.15 0.41 2.255 0.73 ;
      RECT  2.15 0.73 3.46 0.82 ;
      RECT  3.275 0.82 3.46 0.87 ;
      RECT  2.15 0.82 2.24 1.205 ;
      RECT  1.875 1.205 2.515 1.295 ;
      RECT  2.395 1.295 2.515 1.395 ;
      RECT  1.875 1.295 1.995 1.47 ;
      RECT  2.395 1.395 3.055 1.485 ;
      RECT  2.935 1.485 3.055 1.59 ;
      LAYER M2 ;
      RECT  0.785 0.95 5.27 1.05 ;
      RECT  0.51 1.15 5.995 1.25 ;
      LAYER V1 ;
      RECT  0.825 0.95 0.925 1.05 ;
      RECT  5.13 0.95 5.23 1.05 ;
      RECT  0.55 1.15 0.65 1.25 ;
      RECT  5.84 1.15 5.94 1.25 ;
  END
END SEN_ADDH_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_D_4
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_D_4
  CLASS CORE ;
  FOREIGN SEN_ADDH_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 0.91 ;
      RECT  1.95 0.91 2.45 1.09 ;
      RECT  2.35 0.71 2.45 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.369 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 5.085 0.89 ;
      RECT  4.55 0.89 4.65 1.29 ;
      RECT  4.55 1.29 5.25 1.3 ;
      RECT  3.085 0.94 3.45 1.05 ;
      RECT  3.35 1.05 3.45 1.3 ;
      RECT  3.35 1.3 5.25 1.39 ;
      RECT  4.35 1.39 4.45 1.49 ;
      RECT  5.15 1.39 5.25 1.57 ;
      RECT  5.15 1.57 7.13 1.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4068 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.415 4.44 0.475 ;
      RECT  3.79 0.475 4.44 0.595 ;
      RECT  4.15 0.595 4.25 1.04 ;
      RECT  3.79 1.04 4.45 1.16 ;
      RECT  4.335 1.16 4.45 1.21 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.605 0.2 7.855 0.32 ;
      RECT  6.685 0.32 7.855 0.335 ;
      RECT  6.685 0.335 6.85 0.71 ;
      RECT  6.55 0.71 6.85 0.89 ;
      RECT  6.55 0.89 6.71 1.35 ;
      RECT  5.41 1.35 6.71 1.355 ;
      RECT  5.41 1.355 7.74 1.48 ;
    END
    ANTENNADIFFAREA 0.767 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.0 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  1.645 1.44 1.775 1.75 ;
      RECT  2.26 1.18 2.38 1.75 ;
      RECT  2.845 1.435 2.975 1.75 ;
      RECT  3.47 1.48 3.64 1.75 ;
      RECT  4.05 1.48 4.22 1.75 ;
      RECT  4.57 1.48 4.74 1.75 ;
      RECT  4.875 1.61 5.045 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      RECT  5.1 0.05 5.27 0.325 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  4.07 0.05 4.2 0.36 ;
      RECT  3.105 0.05 3.235 0.39 ;
      RECT  3.55 0.05 3.68 0.39 ;
      RECT  4.59 0.05 4.72 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  2.16 0.05 2.25 0.69 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.345 0.19 2.965 0.285 ;
      RECT  2.345 0.285 2.435 0.36 ;
      RECT  2.86 0.285 2.965 0.56 ;
      RECT  2.86 0.56 3.515 0.65 ;
      RECT  5.37 0.31 5.515 0.41 ;
      RECT  5.37 0.41 6.555 0.53 ;
      RECT  6.35 0.53 6.45 1.14 ;
      RECT  5.685 1.14 6.45 1.26 ;
      RECT  4.865 0.25 4.985 0.415 ;
      RECT  4.865 0.415 5.265 0.505 ;
      RECT  5.175 0.505 5.265 0.89 ;
      RECT  5.175 0.89 6.25 1.0 ;
      RECT  5.175 1.0 5.265 1.04 ;
      RECT  4.84 1.04 5.265 1.16 ;
      RECT  1.87 0.29 2.0 0.475 ;
      RECT  1.155 0.475 2.0 0.595 ;
      RECT  1.155 0.595 1.245 0.785 ;
      RECT  0.565 0.785 1.245 0.895 ;
      RECT  1.155 0.895 1.245 1.23 ;
      RECT  1.155 1.23 2.03 1.35 ;
      RECT  1.91 1.35 2.03 1.49 ;
      RECT  0.325 0.475 0.99 0.595 ;
      RECT  0.325 0.595 0.445 1.14 ;
      RECT  0.325 1.14 0.99 1.26 ;
      RECT  6.945 0.45 7.88 0.62 ;
      RECT  7.79 0.62 7.88 1.085 ;
      RECT  7.79 1.085 7.945 1.13 ;
      RECT  6.8 1.075 6.905 1.13 ;
      RECT  6.8 1.13 7.945 1.265 ;
      RECT  2.59 0.45 2.71 0.74 ;
      RECT  2.59 0.74 4.04 0.845 ;
      RECT  2.59 0.845 2.71 1.235 ;
      RECT  2.59 1.235 3.23 1.345 ;
      RECT  3.11 1.345 3.23 1.46 ;
      LAYER M2 ;
      RECT  1.83 0.35 5.54 0.45 ;
      RECT  0.62 1.15 7.2 1.25 ;
      LAYER V1 ;
      RECT  1.885 0.35 1.985 0.45 ;
      RECT  5.4 0.35 5.5 0.45 ;
      RECT  0.66 1.15 0.76 1.25 ;
      RECT  7.06 1.15 7.16 1.25 ;
  END
END SEN_ADDH_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ADDH_D_6
#      Description : "Half adder"
#      Equation    : S=A^B:CO=A&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ADDH_D_6
  CLASS CORE ;
  FOREIGN SEN_ADDH_D_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 0.71 ;
      RECT  2.15 0.71 3.25 0.76 ;
      RECT  2.15 0.76 3.825 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5535 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.51 6.85 0.71 ;
      RECT  6.75 0.71 7.495 0.85 ;
      RECT  6.75 0.85 7.185 0.915 ;
      RECT  6.75 0.915 6.845 1.25 ;
      RECT  4.485 0.94 5.245 1.05 ;
      RECT  5.155 1.05 5.245 1.25 ;
      RECT  5.155 1.25 6.845 1.34 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6102 ;
  END B
  PIN CO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.44 0.37 5.56 0.475 ;
      RECT  5.44 0.475 6.65 0.59 ;
      RECT  6.55 0.31 6.65 0.475 ;
      RECT  6.35 0.59 6.45 0.99 ;
      RECT  5.455 0.99 6.585 1.16 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END CO
  PIN S
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.465 0.21 10.73 0.345 ;
      RECT  10.55 0.345 10.73 0.4 ;
      RECT  10.55 0.4 10.68 1.49 ;
      RECT  9.545 1.48 9.715 1.49 ;
      RECT  7.97 1.49 10.68 1.62 ;
    END
    ANTENNADIFFAREA 1.135 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 10.8 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.625 1.24 1.745 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.18 1.435 3.31 1.75 ;
      RECT  3.625 1.43 3.755 1.75 ;
      RECT  4.145 1.43 4.275 1.75 ;
      RECT  4.665 1.43 4.795 1.75 ;
      RECT  5.175 1.43 5.305 1.75 ;
      RECT  5.695 1.44 5.825 1.75 ;
      RECT  6.215 1.44 6.345 1.75 ;
      RECT  6.735 1.44 6.865 1.75 ;
      RECT  7.285 1.41 7.415 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      RECT  4.405 0.05 4.535 0.345 ;
      RECT  2.14 0.05 2.27 0.35 ;
      RECT  2.66 0.05 2.79 0.35 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  3.18 0.05 3.31 0.36 ;
      RECT  5.695 0.05 5.825 0.36 ;
      RECT  6.215 0.05 6.345 0.36 ;
      RECT  7.255 0.05 7.365 0.36 ;
      RECT  6.74 0.05 6.865 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.07 0.05 5.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.58 0.215 4.26 0.335 ;
      RECT  4.16 0.335 4.26 0.475 ;
      RECT  4.16 0.475 4.85 0.575 ;
      RECT  7.0 0.3 7.12 0.45 ;
      RECT  7.0 0.45 7.675 0.54 ;
      RECT  7.585 0.54 7.675 0.71 ;
      RECT  7.585 0.71 8.07 0.89 ;
      RECT  7.585 0.89 7.675 0.95 ;
      RECT  7.275 0.95 7.675 1.025 ;
      RECT  6.975 1.025 7.675 1.04 ;
      RECT  6.975 1.04 7.365 1.145 ;
      RECT  7.765 0.45 8.935 0.57 ;
      RECT  7.765 0.57 8.3 0.62 ;
      RECT  8.21 0.62 8.3 1.13 ;
      RECT  7.48 1.13 8.3 1.22 ;
      RECT  7.48 1.22 7.66 1.25 ;
      RECT  0.34 0.475 1.54 0.595 ;
      RECT  0.34 0.595 0.47 1.045 ;
      RECT  0.34 1.045 1.535 1.165 ;
      RECT  1.86 0.44 3.045 0.61 ;
      RECT  1.86 0.61 1.99 0.735 ;
      RECT  0.705 0.735 1.99 0.87 ;
      RECT  1.86 0.87 1.99 1.03 ;
      RECT  1.86 1.03 3.03 1.16 ;
      RECT  2.93 1.16 3.03 1.29 ;
      RECT  9.025 0.45 10.455 0.62 ;
      RECT  9.025 0.62 9.155 0.91 ;
      RECT  8.455 0.91 9.155 1.04 ;
      RECT  8.455 1.04 8.595 1.28 ;
      RECT  8.455 1.28 8.92 1.31 ;
      RECT  7.735 1.31 8.92 1.4 ;
      RECT  7.735 1.4 7.855 1.54 ;
      RECT  3.345 0.555 4.035 0.65 ;
      RECT  3.945 0.65 4.035 0.73 ;
      RECT  3.945 0.73 6.175 0.82 ;
      RECT  4.275 0.82 6.175 0.845 ;
      RECT  4.275 0.845 4.365 1.17 ;
      RECT  3.345 1.17 5.035 1.34 ;
      RECT  4.945 1.34 5.035 1.43 ;
      RECT  9.51 0.71 10.3 0.9 ;
      RECT  9.01 1.15 9.19 1.18 ;
      RECT  9.01 1.18 10.46 1.35 ;
      LAYER M2 ;
      RECT  7.69 0.75 9.85 0.85 ;
      RECT  0.325 0.95 8.62 1.05 ;
      RECT  2.89 1.15 9.19 1.25 ;
      LAYER V1 ;
      RECT  7.73 0.75 7.83 0.85 ;
      RECT  7.93 0.75 8.03 0.85 ;
      RECT  9.51 0.75 9.61 0.85 ;
      RECT  9.71 0.75 9.81 0.85 ;
      RECT  0.37 0.95 0.47 1.05 ;
      RECT  8.475 0.95 8.575 1.05 ;
      RECT  2.93 1.15 3.03 1.25 ;
      RECT  7.52 1.15 7.62 1.25 ;
      RECT  9.05 1.15 9.15 1.25 ;
  END
END SEN_ADDH_D_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_1
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_1
  CLASS CORE ;
  FOREIGN SEN_AN2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.22 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.63 1.39 0.77 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.63 0.05 0.77 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.3 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.19 0.18 0.3 ;
      RECT  0.08 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 0.5 ;
      RECT  0.34 0.5 0.85 0.59 ;
      RECT  0.75 0.59 0.85 1.21 ;
      RECT  0.34 1.21 0.85 1.3 ;
      RECT  0.34 1.3 0.455 1.46 ;
  END
END SEN_AN2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_12
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_12
  CLASS CORE ;
  FOREIGN SEN_AN2_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.85 0.91 ;
      RECT  0.55 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5616 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 4.25 0.91 ;
      RECT  2.75 0.91 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5616 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.23 0.19 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.59 1.45 0.71 1.75 ;
      RECT  1.11 1.45 1.23 1.75 ;
      RECT  1.63 1.45 1.75 1.75 ;
      RECT  2.15 1.45 2.27 1.75 ;
      RECT  2.665 1.45 2.795 1.75 ;
      RECT  3.19 1.45 3.31 1.75 ;
      RECT  3.71 1.45 3.83 1.75 ;
      RECT  4.23 1.45 4.35 1.75 ;
      RECT  4.75 1.45 4.87 1.75 ;
      RECT  5.28 1.42 5.4 1.75 ;
      RECT  5.82 1.42 5.94 1.75 ;
      RECT  6.36 1.415 6.48 1.75 ;
      RECT  6.895 1.42 7.025 1.75 ;
      RECT  7.44 1.415 7.56 1.75 ;
      RECT  7.99 1.21 8.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  2.685 0.05 2.79 0.35 ;
      RECT  3.19 0.05 3.31 0.35 ;
      RECT  3.71 0.05 3.83 0.35 ;
      RECT  4.23 0.05 4.35 0.35 ;
      RECT  5.28 0.05 5.4 0.35 ;
      RECT  5.82 0.05 5.94 0.35 ;
      RECT  6.36 0.05 6.48 0.35 ;
      RECT  6.9 0.05 7.02 0.35 ;
      RECT  7.44 0.05 7.56 0.35 ;
      RECT  4.75 0.05 4.87 0.59 ;
      RECT  7.99 0.05 8.11 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.985 0.44 7.855 0.56 ;
      RECT  6.075 0.56 7.06 0.61 ;
      RECT  6.81 0.61 7.06 1.11 ;
      RECT  4.95 1.11 7.85 1.29 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.865 0.185 2.595 0.24 ;
      RECT  0.305 0.24 2.595 0.355 ;
      RECT  2.385 0.355 2.595 0.44 ;
      RECT  2.385 0.44 4.635 0.56 ;
      RECT  2.385 0.56 3.05 0.61 ;
      RECT  4.63 0.755 6.71 0.89 ;
      RECT  4.63 0.89 5.8 0.965 ;
      RECT  4.63 0.965 4.84 1.15 ;
      RECT  2.94 1.15 4.84 1.18 ;
      RECT  0.045 0.445 2.295 0.56 ;
      RECT  1.09 0.56 2.295 0.615 ;
      RECT  2.085 0.615 2.295 1.15 ;
      RECT  1.37 1.15 2.65 1.18 ;
      RECT  1.37 1.18 4.84 1.24 ;
      RECT  0.305 1.24 4.84 1.36 ;
  END
END SEN_AN2_12
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_2
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_2
  CLASS CORE ;
  FOREIGN SEN_AN2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.175 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.575 1.43 0.695 1.75 ;
      RECT  1.195 1.43 1.315 1.75 ;
      RECT  1.815 1.2 1.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.295 0.05 1.415 0.36 ;
      RECT  0.835 0.05 0.955 0.41 ;
      RECT  1.815 0.05 1.935 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.66 1.29 ;
    END
    ANTENNADIFFAREA 0.228 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.17 0.695 0.26 ;
      RECT  0.055 0.26 0.175 0.39 ;
      RECT  0.575 0.26 0.695 0.5 ;
      RECT  0.575 0.5 1.22 0.59 ;
      RECT  1.09 0.42 1.22 0.5 ;
      RECT  1.165 0.75 1.46 0.93 ;
      RECT  1.165 0.93 1.265 1.22 ;
      RECT  0.315 0.36 0.435 0.56 ;
      RECT  0.34 0.56 0.435 1.22 ;
      RECT  0.34 1.22 1.265 1.34 ;
      RECT  0.34 1.34 0.435 1.41 ;
      RECT  0.315 1.41 0.435 1.61 ;
  END
END SEN_AN2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_3
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_3
  CLASS CORE ;
  FOREIGN SEN_AN2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.56 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1404 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1404 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.24 1.225 0.36 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.85 1.45 0.97 1.75 ;
      RECT  1.5 1.45 1.62 1.75 ;
      RECT  2.15 1.43 2.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.11 0.05 1.23 0.35 ;
      RECT  2.15 0.05 2.27 0.37 ;
      RECT  1.63 0.05 1.75 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.89 0.51 2.535 0.69 ;
      RECT  2.35 0.69 2.45 1.11 ;
      RECT  1.89 1.11 2.535 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.305 0.24 0.975 0.36 ;
      RECT  0.85 0.36 0.975 0.44 ;
      RECT  0.85 0.44 1.515 0.56 ;
      RECT  1.56 0.79 2.26 0.89 ;
      RECT  1.56 0.89 1.65 1.24 ;
      RECT  0.045 0.45 0.75 0.555 ;
      RECT  0.65 0.555 0.75 1.24 ;
      RECT  0.565 1.24 1.65 1.36 ;
  END
END SEN_AN2_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_4
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_4
  CLASS CORE ;
  FOREIGN SEN_AN2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.7 1.65 0.91 ;
      RECT  1.15 0.91 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1869 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1869 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.45 0.445 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.845 1.45 0.965 1.75 ;
      RECT  1.365 1.45 1.485 1.75 ;
      RECT  2.11 1.225 2.23 1.75 ;
      RECT  2.69 1.415 2.815 1.75 ;
      RECT  3.215 1.2 3.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.325 0.05 0.445 0.35 ;
      RECT  0.845 0.05 0.965 0.35 ;
      RECT  2.695 0.05 2.815 0.37 ;
      RECT  2.165 0.05 2.285 0.6 ;
      RECT  3.215 0.05 3.335 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.435 0.51 3.06 0.69 ;
      RECT  2.95 0.69 3.06 1.11 ;
      RECT  2.43 1.11 3.06 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.34 0.24 2.015 0.35 ;
      RECT  1.895 0.35 2.015 0.79 ;
      RECT  1.895 0.79 2.86 0.89 ;
      RECT  1.895 0.89 2.015 1.24 ;
      RECT  0.065 1.24 2.015 1.36 ;
      RECT  0.065 1.36 0.185 1.41 ;
      RECT  0.065 0.37 0.19 0.44 ;
      RECT  0.065 0.44 1.77 0.56 ;
  END
END SEN_AN2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_6
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_6
  CLASS CORE ;
  FOREIGN SEN_AN2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 1.05 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.7 2.25 0.89 ;
      RECT  1.55 0.89 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.24 1.21 0.36 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.84 1.45 0.96 1.75 ;
      RECT  1.46 1.45 1.58 1.75 ;
      RECT  2.145 1.45 2.265 1.75 ;
      RECT  2.665 1.2 2.785 1.75 ;
      RECT  3.18 1.44 3.31 1.75 ;
      RECT  3.7 1.43 3.83 1.75 ;
      RECT  4.225 1.425 4.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  3.18 0.05 3.31 0.35 ;
      RECT  3.705 0.05 3.83 0.35 ;
      RECT  4.225 0.05 4.345 0.37 ;
      RECT  2.66 0.05 2.79 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.9 0.44 4.075 0.56 ;
      RECT  3.945 0.56 4.075 1.11 ;
      RECT  2.925 1.11 4.075 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.24 1.485 0.36 ;
      RECT  1.365 0.36 1.485 0.44 ;
      RECT  1.365 0.44 2.55 0.56 ;
      RECT  2.46 0.79 3.72 0.89 ;
      RECT  2.46 0.89 2.55 1.24 ;
      RECT  0.065 0.37 0.19 0.48 ;
      RECT  0.065 0.48 1.26 0.59 ;
      RECT  1.15 0.59 1.26 1.24 ;
      RECT  0.52 1.24 2.55 1.36 ;
  END
END SEN_AN2_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_8
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_8
  CLASS CORE ;
  FOREIGN SEN_AN2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.45 0.91 ;
      RECT  0.35 0.91 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3729 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.7 2.45 0.91 ;
      RECT  2.35 0.91 3.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3729 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.59 1.455 0.71 1.75 ;
      RECT  1.11 1.455 1.23 1.75 ;
      RECT  1.63 1.455 1.75 1.75 ;
      RECT  1.975 1.455 2.095 1.75 ;
      RECT  2.495 1.455 2.615 1.75 ;
      RECT  3.015 1.455 3.135 1.75 ;
      RECT  3.535 1.23 3.655 1.75 ;
      RECT  4.05 1.44 4.18 1.75 ;
      RECT  4.57 1.43 4.7 1.75 ;
      RECT  5.095 1.43 5.215 1.75 ;
      RECT  5.615 1.21 5.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  1.935 0.05 2.105 0.305 ;
      RECT  2.495 0.05 2.615 0.35 ;
      RECT  3.015 0.05 3.135 0.35 ;
      RECT  4.05 0.05 4.18 0.35 ;
      RECT  4.575 0.05 4.7 0.35 ;
      RECT  5.095 0.05 5.215 0.35 ;
      RECT  3.53 0.05 3.66 0.585 ;
      RECT  5.615 0.05 5.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.77 0.44 5.5 0.56 ;
      RECT  3.77 0.56 5.26 0.57 ;
      RECT  5.09 0.57 5.26 1.11 ;
      RECT  3.75 1.11 5.475 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.345 0.205 1.71 0.24 ;
      RECT  0.305 0.24 1.71 0.36 ;
      RECT  1.56 0.36 1.71 0.41 ;
      RECT  1.56 0.41 2.38 0.44 ;
      RECT  1.56 0.44 3.42 0.56 ;
      RECT  3.29 0.775 4.96 0.905 ;
      RECT  3.29 0.905 3.42 1.235 ;
      RECT  0.045 0.45 1.305 0.56 ;
      RECT  1.155 0.56 1.305 0.65 ;
      RECT  1.155 0.65 1.78 0.76 ;
      RECT  1.155 0.76 1.305 1.235 ;
      RECT  1.155 1.235 3.42 1.24 ;
      RECT  0.305 1.24 3.42 1.365 ;
  END
END SEN_AN2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_16
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_16
  CLASS CORE ;
  FOREIGN SEN_AN2_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.47 6.85 0.97 ;
      RECT  5.75 0.51 5.85 0.96 ;
      RECT  4.75 0.51 4.85 0.96 ;
      RECT  3.55 0.51 3.65 0.96 ;
      RECT  2.55 0.47 2.65 0.96 ;
      RECT  1.55 0.47 1.65 0.96 ;
      RECT  0.55 0.47 0.65 0.96 ;
      LAYER M2 ;
      RECT  0.51 0.55 6.89 0.65 ;
      LAYER V1 ;
      RECT  6.75 0.55 6.85 0.65 ;
      RECT  5.75 0.55 5.85 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.55 0.55 3.65 0.65 ;
      RECT  2.55 0.55 2.65 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7476 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.07 0.71 7.18 1.1 ;
      RECT  6.15 0.71 6.45 0.89 ;
      RECT  5.15 0.71 5.455 0.89 ;
      RECT  3.95 0.71 4.25 0.89 ;
      RECT  2.95 0.71 3.25 0.89 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.145 0.71 0.455 0.89 ;
      LAYER M2 ;
      RECT  0.11 0.75 7.215 0.85 ;
      LAYER V1 ;
      RECT  7.075 0.75 7.175 0.85 ;
      RECT  6.15 0.75 6.25 0.85 ;
      RECT  6.35 0.75 6.45 0.85 ;
      RECT  5.15 0.75 5.25 0.85 ;
      RECT  5.355 0.75 5.455 0.85 ;
      RECT  3.95 0.75 4.05 0.85 ;
      RECT  4.15 0.75 4.25 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  3.15 0.75 3.25 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  0.95 0.75 1.05 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  0.15 0.75 0.25 0.85 ;
      RECT  0.355 0.75 0.455 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7476 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.965 1.41 1.095 1.75 ;
      RECT  0.0 1.75 11.6 1.85 ;
      RECT  1.51 1.41 1.64 1.75 ;
      RECT  2.03 1.41 2.16 1.75 ;
      RECT  2.55 1.41 2.68 1.75 ;
      RECT  3.07 1.41 3.2 1.75 ;
      RECT  3.59 1.41 3.72 1.75 ;
      RECT  4.11 1.41 4.24 1.75 ;
      RECT  4.63 1.41 4.76 1.75 ;
      RECT  5.15 1.41 5.28 1.75 ;
      RECT  5.67 1.41 5.8 1.75 ;
      RECT  6.22 1.41 6.35 1.75 ;
      RECT  7.21 1.41 7.34 1.75 ;
      RECT  7.77 1.41 7.9 1.75 ;
      RECT  8.29 1.41 8.42 1.75 ;
      RECT  8.81 1.41 8.94 1.75 ;
      RECT  9.33 1.41 9.46 1.75 ;
      RECT  9.85 1.41 9.965 1.75 ;
      RECT  10.37 1.41 10.5 1.75 ;
      RECT  10.89 1.41 11.02 1.75 ;
      RECT  11.415 1.21 11.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.6 0.05 ;
      RECT  7.77 0.05 7.9 0.385 ;
      RECT  8.29 0.05 8.42 0.385 ;
      RECT  9.33 0.05 9.46 0.385 ;
      RECT  10.37 0.05 10.5 0.385 ;
      RECT  10.89 0.05 11.02 0.385 ;
      RECT  7.24 0.05 7.37 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  0.995 0.05 1.115 0.59 ;
      RECT  2.035 0.05 2.155 0.59 ;
      RECT  3.075 0.05 3.195 0.59 ;
      RECT  4.115 0.05 4.235 0.59 ;
      RECT  5.155 0.05 5.275 0.59 ;
      RECT  6.195 0.05 6.315 0.59 ;
      RECT  8.815 0.05 8.935 0.59 ;
      RECT  9.855 0.05 9.975 0.59 ;
      RECT  11.415 0.05 11.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.09 0.475 11.3 0.595 ;
      RECT  10.35 0.595 10.45 1.11 ;
      RECT  9.045 0.475 9.74 0.595 ;
      RECT  9.15 0.595 9.25 1.11 ;
      RECT  7.49 0.475 8.7 0.595 ;
      RECT  8.35 0.595 8.45 1.11 ;
      RECT  7.515 1.11 11.275 1.29 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.54 0.24 7.12 0.36 ;
      RECT  7.0 0.36 7.12 0.49 ;
      RECT  6.54 0.36 6.66 1.085 ;
      RECT  7.0 0.49 7.395 0.61 ;
      RECT  7.275 0.61 7.395 0.71 ;
      RECT  7.275 0.71 8.185 0.96 ;
      RECT  7.275 0.96 7.405 1.19 ;
      RECT  5.55 0.24 5.85 0.36 ;
      RECT  5.55 0.36 5.65 1.085 ;
      RECT  5.55 1.085 6.66 1.115 ;
      RECT  4.55 0.24 4.81 0.36 ;
      RECT  4.55 0.36 4.65 1.115 ;
      RECT  4.55 1.115 6.66 1.145 ;
      RECT  3.54 0.24 3.85 0.36 ;
      RECT  3.75 0.36 3.85 1.145 ;
      RECT  3.75 1.145 6.66 1.17 ;
      RECT  2.5 0.24 2.85 0.36 ;
      RECT  2.75 0.36 2.85 1.17 ;
      RECT  2.75 1.17 6.66 1.19 ;
      RECT  2.75 1.19 7.405 1.2 ;
      RECT  1.46 0.24 1.85 0.36 ;
      RECT  1.75 0.36 1.85 1.2 ;
      RECT  0.47 0.24 0.85 0.36 ;
      RECT  0.75 0.36 0.85 1.2 ;
      RECT  0.75 1.2 7.405 1.32 ;
      RECT  8.55 0.71 9.05 0.89 ;
      RECT  9.35 0.71 10.05 0.89 ;
      RECT  10.55 0.71 11.25 0.89 ;
      LAYER M2 ;
      RECT  7.61 0.75 11.19 0.85 ;
      LAYER V1 ;
      RECT  7.65 0.75 7.75 0.85 ;
      RECT  7.85 0.75 7.95 0.85 ;
      RECT  8.05 0.75 8.15 0.85 ;
      RECT  8.65 0.75 8.75 0.85 ;
      RECT  8.85 0.75 8.95 0.85 ;
      RECT  9.45 0.75 9.55 0.85 ;
      RECT  9.65 0.75 9.75 0.85 ;
      RECT  9.85 0.75 9.95 0.85 ;
      RECT  10.65 0.75 10.75 0.85 ;
      RECT  10.85 0.75 10.95 0.85 ;
      RECT  11.05 0.75 11.15 0.85 ;
  END
END SEN_AN2_16
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_24
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_24
  CLASS CORE ;
  FOREIGN SEN_AN2_24 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.24 0.51 10.34 0.93 ;
      RECT  9.35 0.47 9.45 0.91 ;
      RECT  8.15 0.49 8.25 0.93 ;
      RECT  7.15 0.49 7.25 0.95 ;
      RECT  6.15 0.49 6.25 0.95 ;
      RECT  5.15 0.49 5.25 0.95 ;
      RECT  4.145 0.49 4.245 0.95 ;
      RECT  2.95 0.47 3.05 0.95 ;
      RECT  1.95 0.47 2.05 0.95 ;
      RECT  0.95 0.47 1.05 0.95 ;
      RECT  0.15 0.49 0.25 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.55 10.38 0.65 ;
      LAYER V1 ;
      RECT  10.24 0.55 10.34 0.65 ;
      RECT  9.35 0.55 9.45 0.65 ;
      RECT  8.15 0.55 8.25 0.65 ;
      RECT  7.15 0.55 7.25 0.65 ;
      RECT  6.15 0.55 6.25 0.65 ;
      RECT  5.15 0.55 5.25 0.65 ;
      RECT  4.145 0.55 4.245 0.65 ;
      RECT  2.95 0.55 3.05 0.65 ;
      RECT  1.95 0.55 2.05 0.65 ;
      RECT  0.95 0.55 1.05 0.65 ;
      RECT  0.15 0.55 0.25 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1214 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.53 0.71 10.65 1.07 ;
      RECT  9.55 0.71 9.85 0.89 ;
      RECT  8.75 0.71 9.05 0.89 ;
      RECT  7.55 0.71 7.85 0.89 ;
      RECT  6.55 0.71 6.85 0.89 ;
      RECT  5.55 0.71 5.855 0.89 ;
      RECT  4.55 0.71 4.85 0.89 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  2.35 0.71 2.65 0.89 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  0.55 0.71 0.855 0.89 ;
      LAYER M2 ;
      RECT  0.51 0.75 10.69 0.85 ;
      LAYER V1 ;
      RECT  10.55 0.75 10.65 0.85 ;
      RECT  9.55 0.75 9.65 0.85 ;
      RECT  9.75 0.75 9.85 0.85 ;
      RECT  8.75 0.75 8.85 0.85 ;
      RECT  8.95 0.75 9.05 0.85 ;
      RECT  7.55 0.75 7.65 0.85 ;
      RECT  7.75 0.75 7.85 0.85 ;
      RECT  6.55 0.75 6.65 0.85 ;
      RECT  6.75 0.75 6.85 0.85 ;
      RECT  5.55 0.75 5.65 0.85 ;
      RECT  5.755 0.75 5.855 0.85 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.35 0.75 2.45 0.85 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
      RECT  0.755 0.75 0.855 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1214 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.47 1.41 1.6 1.75 ;
      RECT  0.0 1.75 17.2 1.85 ;
      RECT  1.99 1.41 2.12 1.75 ;
      RECT  2.51 1.41 2.64 1.75 ;
      RECT  3.03 1.41 3.16 1.75 ;
      RECT  3.55 1.41 3.68 1.75 ;
      RECT  4.07 1.41 4.2 1.75 ;
      RECT  4.59 1.41 4.72 1.75 ;
      RECT  5.11 1.41 5.24 1.75 ;
      RECT  5.63 1.41 5.76 1.75 ;
      RECT  6.15 1.41 6.28 1.75 ;
      RECT  6.67 1.41 6.8 1.75 ;
      RECT  7.19 1.41 7.32 1.75 ;
      RECT  7.71 1.41 7.84 1.75 ;
      RECT  8.23 1.41 8.36 1.75 ;
      RECT  8.75 1.41 8.88 1.75 ;
      RECT  9.27 1.41 9.4 1.75 ;
      RECT  10.7 1.41 10.83 1.75 ;
      RECT  11.275 1.41 11.405 1.75 ;
      RECT  11.795 1.41 11.925 1.75 ;
      RECT  12.315 1.41 12.445 1.75 ;
      RECT  12.835 1.41 12.965 1.75 ;
      RECT  13.355 1.41 13.485 1.75 ;
      RECT  13.875 1.41 14.005 1.75 ;
      RECT  14.395 1.41 14.525 1.75 ;
      RECT  14.915 1.41 15.045 1.75 ;
      RECT  15.435 1.41 15.565 1.75 ;
      RECT  15.95 1.41 16.085 1.75 ;
      RECT  16.47 1.41 16.605 1.75 ;
      RECT  17.0 1.21 17.12 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 17.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
      RECT  11.85 1.75 11.95 1.85 ;
      RECT  12.45 1.75 12.55 1.85 ;
      RECT  13.05 1.75 13.15 1.85 ;
      RECT  13.65 1.75 13.75 1.85 ;
      RECT  14.25 1.75 14.35 1.85 ;
      RECT  14.85 1.75 14.95 1.85 ;
      RECT  15.45 1.75 15.55 1.85 ;
      RECT  16.05 1.75 16.15 1.85 ;
      RECT  16.65 1.75 16.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 17.2 0.05 ;
      RECT  10.725 0.05 10.855 0.37 ;
      RECT  11.275 0.05 11.405 0.385 ;
      RECT  11.795 0.05 11.925 0.385 ;
      RECT  12.835 0.05 12.965 0.385 ;
      RECT  13.875 0.05 14.005 0.385 ;
      RECT  14.915 0.05 15.045 0.385 ;
      RECT  15.955 0.05 16.085 0.385 ;
      RECT  16.475 0.05 16.605 0.385 ;
      RECT  0.54 0.05 0.66 0.59 ;
      RECT  1.475 0.05 1.595 0.59 ;
      RECT  2.515 0.05 2.635 0.59 ;
      RECT  3.555 0.05 3.675 0.59 ;
      RECT  4.595 0.05 4.715 0.59 ;
      RECT  5.635 0.05 5.755 0.59 ;
      RECT  6.675 0.05 6.795 0.59 ;
      RECT  7.715 0.05 7.835 0.59 ;
      RECT  8.755 0.05 8.875 0.59 ;
      RECT  9.74 0.05 9.86 0.59 ;
      RECT  12.32 0.05 12.44 0.59 ;
      RECT  13.36 0.05 13.48 0.59 ;
      RECT  14.4 0.05 14.52 0.59 ;
      RECT  15.44 0.05 15.56 0.59 ;
      RECT  17.0 0.05 17.12 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 17.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
      RECT  11.85 -0.05 11.95 0.05 ;
      RECT  12.45 -0.05 12.55 0.05 ;
      RECT  13.05 -0.05 13.15 0.05 ;
      RECT  13.65 -0.05 13.75 0.05 ;
      RECT  14.25 -0.05 14.35 0.05 ;
      RECT  14.85 -0.05 14.95 0.05 ;
      RECT  15.45 -0.05 15.55 0.05 ;
      RECT  16.05 -0.05 16.15 0.05 ;
      RECT  16.65 -0.05 16.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  15.675 0.475 16.885 0.595 ;
      RECT  15.94 0.595 16.065 1.11 ;
      RECT  14.635 0.475 15.325 0.595 ;
      RECT  14.95 0.595 15.05 1.11 ;
      RECT  13.595 0.475 14.285 0.595 ;
      RECT  13.75 0.595 13.85 1.11 ;
      RECT  12.55 0.475 13.245 0.595 ;
      RECT  12.55 0.595 12.65 1.11 ;
      RECT  10.995 0.475 12.205 0.595 ;
      RECT  11.74 0.595 11.87 1.11 ;
      RECT  11.02 1.11 16.905 1.29 ;
    END
    ANTENNADIFFAREA 2.592 ;
  END X
  OBS
      LAYER M1 ;
      RECT  9.975 0.22 10.6 0.38 ;
      RECT  10.44 0.38 10.6 0.46 ;
      RECT  9.975 0.38 10.135 1.0 ;
      RECT  10.44 0.46 10.9 0.62 ;
      RECT  10.74 0.62 10.9 0.71 ;
      RECT  10.74 0.71 11.65 0.95 ;
      RECT  10.74 0.95 10.9 1.16 ;
      RECT  9.15 0.24 9.45 0.36 ;
      RECT  9.15 0.36 9.25 1.0 ;
      RECT  9.15 1.0 10.135 1.025 ;
      RECT  8.18 0.24 8.445 0.36 ;
      RECT  8.345 0.36 8.445 1.025 ;
      RECT  8.345 1.025 10.135 1.055 ;
      RECT  7.14 0.24 7.45 0.36 ;
      RECT  7.35 0.36 7.45 1.055 ;
      RECT  7.35 1.055 10.135 1.085 ;
      RECT  6.1 0.24 6.45 0.36 ;
      RECT  6.35 0.36 6.45 1.085 ;
      RECT  6.35 1.085 10.135 1.115 ;
      RECT  4.95 0.24 5.29 0.36 ;
      RECT  4.95 0.36 5.05 1.115 ;
      RECT  4.95 1.115 10.135 1.145 ;
      RECT  3.95 0.24 4.25 0.36 ;
      RECT  3.95 0.36 4.05 1.145 ;
      RECT  3.95 1.145 10.135 1.16 ;
      RECT  3.95 1.16 10.9 1.17 ;
      RECT  2.98 0.24 3.25 0.36 ;
      RECT  3.15 0.36 3.25 1.17 ;
      RECT  3.15 1.17 10.9 1.2 ;
      RECT  1.94 0.24 2.25 0.36 ;
      RECT  2.15 0.36 2.25 1.2 ;
      RECT  0.95 0.24 1.25 0.36 ;
      RECT  1.15 0.36 1.25 1.2 ;
      RECT  1.15 1.2 10.9 1.23 ;
      RECT  0.075 0.17 0.195 0.27 ;
      RECT  0.075 0.27 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.23 ;
      RECT  0.35 1.23 10.9 1.32 ;
      RECT  11.96 0.71 12.45 0.89 ;
      RECT  12.75 0.71 13.45 0.89 ;
      RECT  14.15 0.71 14.85 0.89 ;
      RECT  15.15 0.71 15.65 0.89 ;
      RECT  16.165 0.71 16.85 0.89 ;
      LAYER M2 ;
      RECT  10.81 0.75 16.79 0.85 ;
      LAYER V1 ;
      RECT  10.85 0.75 10.95 0.85 ;
      RECT  11.05 0.75 11.15 0.85 ;
      RECT  11.25 0.75 11.35 0.85 ;
      RECT  11.45 0.75 11.55 0.85 ;
      RECT  12.05 0.75 12.15 0.85 ;
      RECT  12.25 0.75 12.35 0.85 ;
      RECT  12.85 0.75 12.95 0.85 ;
      RECT  13.05 0.75 13.15 0.85 ;
      RECT  13.25 0.75 13.35 0.85 ;
      RECT  14.25 0.75 14.35 0.85 ;
      RECT  14.45 0.75 14.55 0.85 ;
      RECT  14.65 0.75 14.75 0.85 ;
      RECT  15.25 0.75 15.35 0.85 ;
      RECT  15.45 0.75 15.55 0.85 ;
      RECT  16.25 0.75 16.35 0.85 ;
      RECT  16.45 0.75 16.55 0.85 ;
      RECT  16.65 0.75 16.75 0.85 ;
  END
END SEN_AN2_24
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_DG_1
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_DG_1
  CLASS CORE ;
  FOREIGN SEN_AN2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.41 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.62 1.41 0.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.62 0.05 0.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.31 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.17 0.19 0.3 ;
      RECT  0.07 0.3 0.45 0.39 ;
      RECT  0.36 0.39 0.45 0.5 ;
      RECT  0.36 0.5 0.85 0.59 ;
      RECT  0.75 0.59 0.85 1.21 ;
      RECT  0.34 1.21 0.85 1.3 ;
      RECT  0.34 1.3 0.455 1.61 ;
  END
END SEN_AN2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_DG_16
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_DG_16
  CLASS CORE ;
  FOREIGN SEN_AN2_DG_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  0.595 1.42 0.725 1.75 ;
      RECT  1.115 1.42 1.245 1.75 ;
      RECT  1.635 1.42 1.765 1.75 ;
      RECT  2.28 1.21 2.4 1.75 ;
      RECT  2.89 1.415 3.02 1.75 ;
      RECT  3.41 1.415 3.54 1.75 ;
      RECT  3.93 1.415 4.06 1.75 ;
      RECT  4.45 1.415 4.58 1.75 ;
      RECT  4.97 1.415 5.1 1.75 ;
      RECT  5.49 1.415 5.62 1.75 ;
      RECT  6.01 1.415 6.14 1.75 ;
      RECT  6.555 1.395 6.685 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  0.34 0.05 0.46 0.365 ;
      RECT  0.86 0.05 0.98 0.365 ;
      RECT  2.63 0.05 2.76 0.39 ;
      RECT  3.15 0.05 3.28 0.39 ;
      RECT  3.67 0.05 3.8 0.39 ;
      RECT  4.19 0.05 4.32 0.39 ;
      RECT  4.71 0.05 4.84 0.39 ;
      RECT  5.23 0.05 5.36 0.39 ;
      RECT  5.75 0.05 5.88 0.39 ;
      RECT  6.27 0.05 6.4 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.335 0.5 6.67 0.69 ;
      RECT  2.335 0.69 5.45 0.7 ;
      RECT  5.13 0.7 5.45 1.11 ;
      RECT  2.55 1.11 6.48 1.31 ;
    END
    ANTENNADIFFAREA 1.776 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.115 0.22 2.33 0.34 ;
      RECT  1.115 0.34 1.245 0.46 ;
      RECT  0.08 0.37 0.2 0.46 ;
      RECT  0.08 0.46 1.245 0.59 ;
      RECT  1.34 0.475 2.055 0.595 ;
      RECT  1.96 0.595 2.055 0.795 ;
      RECT  1.96 0.795 4.98 0.885 ;
      RECT  1.96 0.885 2.055 1.21 ;
      RECT  0.315 1.21 2.055 1.33 ;
  END
END SEN_AN2_DG_16
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_DG_2
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_DG_2
  CLASS CORE ;
  FOREIGN SEN_AN2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.18 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.58 1.41 0.7 1.75 ;
      RECT  1.17 1.21 1.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.58 0.05 0.7 0.39 ;
      RECT  1.17 0.05 1.27 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.83 0.24 1.05 0.36 ;
      RECT  0.95 0.36 1.05 1.24 ;
      RECT  0.81 1.24 1.05 1.36 ;
    END
    ANTENNADIFFAREA 0.26 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.2 0.19 0.33 ;
      RECT  0.07 0.33 0.445 0.42 ;
      RECT  0.355 0.42 0.445 0.48 ;
      RECT  0.355 0.48 0.845 0.57 ;
      RECT  0.755 0.57 0.845 1.055 ;
      RECT  0.55 1.055 0.845 1.145 ;
      RECT  0.55 1.145 0.65 1.21 ;
      RECT  0.32 1.21 0.65 1.31 ;
      RECT  0.32 1.31 0.44 1.54 ;
  END
END SEN_AN2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_DG_3
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_DG_3
  CLASS CORE ;
  FOREIGN SEN_AN2_DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.18 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.58 1.42 0.7 1.75 ;
      RECT  1.12 1.445 1.24 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  1.14 0.05 1.26 0.39 ;
      RECT  0.58 0.05 0.7 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.815 0.255 1.05 0.345 ;
      RECT  0.95 0.345 1.05 0.51 ;
      RECT  0.95 0.51 1.51 0.69 ;
      RECT  1.35 0.69 1.45 1.235 ;
      RECT  0.815 1.235 1.545 1.355 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.06 0.17 0.18 0.3 ;
      RECT  0.06 0.3 0.445 0.39 ;
      RECT  0.355 0.39 0.445 0.53 ;
      RECT  0.355 0.53 0.845 0.62 ;
      RECT  0.755 0.62 0.845 0.785 ;
      RECT  0.755 0.785 1.24 0.895 ;
      RECT  0.755 0.895 0.845 1.055 ;
      RECT  0.55 1.055 0.845 1.145 ;
      RECT  0.55 1.145 0.65 1.21 ;
      RECT  0.295 1.21 0.65 1.33 ;
  END
END SEN_AN2_DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_DG_4
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_DG_4
  CLASS CORE ;
  FOREIGN SEN_AN2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.9 ;
      RECT  0.35 0.9 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.575 1.41 0.705 1.75 ;
      RECT  1.095 1.435 1.225 1.75 ;
      RECT  1.615 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.58 0.05 0.7 0.39 ;
      RECT  1.115 0.05 1.215 0.39 ;
      RECT  1.62 0.05 1.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.815 0.255 1.025 0.345 ;
      RECT  0.935 0.345 1.025 0.48 ;
      RECT  0.935 0.48 1.505 0.59 ;
      RECT  1.35 0.59 1.45 1.22 ;
      RECT  1.35 1.22 1.505 1.225 ;
      RECT  0.815 1.225 1.505 1.345 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.06 0.17 0.18 0.3 ;
      RECT  0.06 0.3 0.445 0.39 ;
      RECT  0.355 0.39 0.445 0.48 ;
      RECT  0.355 0.48 0.845 0.57 ;
      RECT  0.755 0.57 0.845 0.785 ;
      RECT  0.755 0.785 1.24 0.895 ;
      RECT  0.755 0.895 0.845 1.045 ;
      RECT  0.55 1.045 0.845 1.135 ;
      RECT  0.55 1.135 0.65 1.21 ;
      RECT  0.295 1.21 0.65 1.32 ;
  END
END SEN_AN2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_DG_8
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_DG_8
  CLASS CORE ;
  FOREIGN SEN_AN2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.945 0.89 ;
      RECT  0.75 0.89 0.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.595 1.42 0.725 1.75 ;
      RECT  1.24 1.21 1.36 1.75 ;
      RECT  1.84 1.415 1.99 1.75 ;
      RECT  2.36 1.415 2.51 1.75 ;
      RECT  2.88 1.415 3.03 1.75 ;
      RECT  3.415 1.21 3.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.34 0.05 0.46 0.37 ;
      RECT  1.58 0.05 1.725 0.385 ;
      RECT  2.1 0.05 2.25 0.385 ;
      RECT  2.615 0.05 2.77 0.385 ;
      RECT  3.14 0.05 3.29 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.295 0.51 3.54 0.69 ;
      RECT  2.68 0.69 2.85 1.11 ;
      RECT  1.54 1.11 3.3 1.29 ;
    END
    ANTENNADIFFAREA 0.912 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.595 0.23 1.29 0.345 ;
      RECT  0.595 0.345 0.725 0.46 ;
      RECT  0.08 0.37 0.2 0.46 ;
      RECT  0.08 0.46 0.725 0.59 ;
      RECT  0.82 0.48 1.135 0.6 ;
      RECT  1.04 0.6 1.135 0.785 ;
      RECT  1.04 0.785 2.555 0.895 ;
      RECT  1.04 0.895 1.135 1.21 ;
      RECT  0.315 1.21 1.135 1.33 ;
  END
END SEN_AN2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_S_0P5
#      Description : "2-Input AND, symmetric rise/fall"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_S_0P5
  CLASS CORE ;
  FOREIGN SEN_AN2_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0201 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0201 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.41 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.62 1.41 0.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.62 0.05 0.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.22 1.05 1.55 ;
    END
    ANTENNADIFFAREA 0.108 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.17 0.19 0.28 ;
      RECT  0.07 0.28 0.43 0.39 ;
      RECT  0.34 0.39 0.43 0.48 ;
      RECT  0.34 0.48 0.85 0.57 ;
      RECT  0.75 0.57 0.85 1.21 ;
      RECT  0.34 1.21 0.85 1.3 ;
      RECT  0.34 1.3 0.455 1.63 ;
  END
END SEN_AN2_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_S_1
#      Description : "2-Input AND, symmetric rise/fall"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_S_1
  CLASS CORE ;
  FOREIGN SEN_AN2_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.41 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.615 1.41 0.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.615 0.05 0.745 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.31 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.17 0.2 0.27 ;
      RECT  0.08 0.27 0.43 0.39 ;
      RECT  0.34 0.39 0.43 0.48 ;
      RECT  0.34 0.48 0.85 0.57 ;
      RECT  0.75 0.57 0.85 1.23 ;
      RECT  0.34 1.23 0.85 1.32 ;
      RECT  0.34 1.32 0.455 1.59 ;
  END
END SEN_AN2_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_S_16
#      Description : "2-Input AND, symmetric rise/fall"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_S_16
  CLASS CORE ;
  FOREIGN SEN_AN2_S_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  0.75 0.91 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4932 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 3.85 0.91 ;
      RECT  2.75 0.91 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4932 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  1.62 1.44 1.75 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  2.66 1.44 2.79 1.75 ;
      RECT  3.18 1.44 3.31 1.75 ;
      RECT  3.7 1.44 3.83 1.75 ;
      RECT  4.35 1.21 4.47 1.75 ;
      RECT  4.97 1.41 5.1 1.75 ;
      RECT  5.49 1.41 5.62 1.75 ;
      RECT  6.01 1.41 6.14 1.75 ;
      RECT  6.53 1.41 6.66 1.75 ;
      RECT  7.05 1.41 7.18 1.75 ;
      RECT  7.57 1.41 7.7 1.75 ;
      RECT  8.09 1.41 8.22 1.75 ;
      RECT  8.615 1.21 8.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  4.95 0.05 5.12 0.325 ;
      RECT  5.47 0.05 5.64 0.325 ;
      RECT  5.99 0.05 6.16 0.325 ;
      RECT  6.51 0.05 6.68 0.325 ;
      RECT  7.03 0.05 7.2 0.325 ;
      RECT  7.55 0.05 7.72 0.325 ;
      RECT  8.095 0.05 8.215 0.37 ;
      RECT  2.405 0.05 2.53 0.38 ;
      RECT  2.92 0.05 3.05 0.38 ;
      RECT  3.44 0.05 3.57 0.38 ;
      RECT  3.96 0.05 4.09 0.38 ;
      RECT  4.46 0.05 4.575 0.59 ;
      RECT  8.615 0.05 8.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.69 0.415 7.65 0.51 ;
      RECT  4.69 0.51 8.5 0.545 ;
      RECT  6.24 0.545 8.5 0.635 ;
      RECT  7.33 0.635 8.5 0.69 ;
      RECT  7.33 0.69 7.65 1.07 ;
      RECT  6.245 1.07 7.65 1.11 ;
      RECT  4.69 1.11 8.5 1.29 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.605 0.195 2.29 0.235 ;
      RECT  0.065 0.235 2.29 0.365 ;
      RECT  0.065 0.365 0.185 0.46 ;
      RECT  2.08 0.365 2.29 0.48 ;
      RECT  2.08 0.48 4.37 0.61 ;
      RECT  2.08 0.61 2.81 0.65 ;
      RECT  4.1 0.765 7.225 0.91 ;
      RECT  4.1 0.91 4.24 1.215 ;
      RECT  0.3 0.455 1.99 0.585 ;
      RECT  1.86 0.585 1.99 1.205 ;
      RECT  0.3 1.205 1.99 1.215 ;
      RECT  0.3 1.215 4.24 1.345 ;
  END
END SEN_AN2_S_16
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_S_1P5
#      Description : "2-Input AND, symmetric rise/fall"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_S_1P5
  CLASS CORE ;
  FOREIGN SEN_AN2_S_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0498 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.95 ;
      RECT  0.35 0.95 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0498 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.585 1.39 0.71 1.75 ;
      RECT  1.14 1.21 1.25 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.585 0.05 0.715 0.39 ;
      RECT  1.14 0.05 1.25 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.825 0.24 1.05 0.36 ;
      RECT  0.95 0.36 1.05 1.255 ;
      RECT  0.825 1.255 1.05 1.375 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.17 0.19 0.3 ;
      RECT  0.07 0.3 0.445 0.39 ;
      RECT  0.355 0.39 0.445 0.48 ;
      RECT  0.355 0.48 0.845 0.57 ;
      RECT  0.755 0.57 0.845 1.055 ;
      RECT  0.55 1.055 0.845 1.145 ;
      RECT  0.55 1.145 0.65 1.21 ;
      RECT  0.33 1.21 0.65 1.3 ;
      RECT  0.33 1.3 0.45 1.48 ;
  END
END SEN_AN2_S_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_S_2
#      Description : "2-Input AND, symmetric rise/fall"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_S_2
  CLASS CORE ;
  FOREIGN SEN_AN2_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.7 1.05 0.9 ;
      RECT  0.75 0.9 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.38 0.185 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.64 1.415 0.79 1.75 ;
      RECT  1.245 1.4 1.395 1.75 ;
      RECT  1.82 1.41 1.94 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.755 0.05 0.905 0.23 ;
      RECT  1.29 0.05 1.435 0.39 ;
      RECT  1.82 0.05 1.94 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.85 0.69 ;
      RECT  1.75 0.69 1.85 1.11 ;
      RECT  1.55 1.11 1.85 1.295 ;
    END
    ANTENNADIFFAREA 0.232 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.325 0.19 0.445 0.32 ;
      RECT  0.325 0.32 1.16 0.41 ;
      RECT  1.04 0.19 1.16 0.32 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 1.44 0.59 ;
      RECT  1.35 0.59 1.44 0.785 ;
      RECT  1.35 0.785 1.64 0.895 ;
      RECT  1.35 0.895 1.44 1.21 ;
      RECT  0.325 1.21 1.44 1.3 ;
      RECT  0.325 1.3 0.445 1.54 ;
      RECT  0.975 1.3 1.095 1.54 ;
  END
END SEN_AN2_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_S_3
#      Description : "2-Input AND, symmetric rise/fall"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_S_3
  CLASS CORE ;
  FOREIGN SEN_AN2_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.75 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0984 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0984 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.575 1.46 0.745 1.75 ;
      RECT  1.09 1.465 1.27 1.75 ;
      RECT  1.37 1.21 1.49 1.75 ;
      RECT  1.885 1.41 2.015 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.33 0.05 0.465 0.37 ;
      RECT  1.885 0.05 2.015 0.39 ;
      RECT  1.37 0.05 1.49 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.615 0.51 2.265 0.69 ;
      RECT  2.15 0.69 2.265 1.11 ;
      RECT  1.61 1.11 2.265 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.595 0.235 1.28 0.36 ;
      RECT  0.595 0.36 0.725 0.46 ;
      RECT  0.08 0.37 0.2 0.46 ;
      RECT  0.08 0.46 0.725 0.59 ;
      RECT  0.82 0.465 1.255 0.59 ;
      RECT  1.16 0.59 1.255 0.795 ;
      RECT  1.16 0.795 2.03 0.885 ;
      RECT  1.16 0.885 1.255 1.26 ;
      RECT  0.315 1.26 1.255 1.37 ;
  END
END SEN_AN2_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_S_4
#      Description : "2-Input AND, symmetric rise/fall"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_S_4
  CLASS CORE ;
  FOREIGN SEN_AN2_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.6 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.45 0.91 ;
      RECT  0.95 0.91 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1608 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.23 0.19 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.61 1.45 0.73 1.75 ;
      RECT  1.13 1.45 1.25 1.75 ;
      RECT  1.74 1.225 1.86 1.75 ;
      RECT  2.255 1.415 2.38 1.75 ;
      RECT  2.78 1.21 2.9 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  1.13 0.05 1.25 0.35 ;
      RECT  2.26 0.05 2.38 0.37 ;
      RECT  2.78 0.05 2.9 0.59 ;
      RECT  1.695 0.05 1.815 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.66 0.69 ;
      RECT  2.55 0.69 2.66 1.11 ;
      RECT  1.95 1.11 2.66 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.32 0.24 0.99 0.355 ;
      RECT  0.87 0.355 0.99 0.44 ;
      RECT  0.87 0.44 1.57 0.56 ;
      RECT  1.55 0.79 2.425 0.89 ;
      RECT  1.55 0.89 1.65 1.24 ;
      RECT  0.09 0.34 0.21 0.445 ;
      RECT  0.09 0.445 0.78 0.56 ;
      RECT  0.69 0.56 0.78 1.24 ;
      RECT  0.325 1.24 1.65 1.36 ;
  END
END SEN_AN2_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_S_8
#      Description : "2-Input AND, symmetric rise/fall"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_S_8
  CLASS CORE ;
  FOREIGN SEN_AN2_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.45 0.91 ;
      RECT  0.35 0.91 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3207 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 0.91 ;
      RECT  1.75 0.91 2.495 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3207 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.455 0.45 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  0.85 1.455 0.97 1.75 ;
      RECT  1.37 1.455 1.49 1.75 ;
      RECT  1.89 1.455 2.01 1.75 ;
      RECT  2.41 1.455 2.53 1.75 ;
      RECT  2.975 1.21 3.095 1.75 ;
      RECT  3.55 1.44 3.68 1.75 ;
      RECT  4.1 1.43 4.23 1.75 ;
      RECT  4.655 1.43 4.775 1.75 ;
      RECT  5.21 1.21 5.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  1.89 0.05 2.01 0.35 ;
      RECT  2.41 0.05 2.53 0.35 ;
      RECT  3.55 0.05 3.68 0.35 ;
      RECT  4.105 0.05 4.23 0.35 ;
      RECT  4.655 0.05 4.775 0.35 ;
      RECT  2.97 0.05 3.095 0.585 ;
      RECT  5.21 0.05 5.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.225 0.44 5.075 0.56 ;
      RECT  3.225 0.56 4.86 0.57 ;
      RECT  4.69 0.57 4.86 1.11 ;
      RECT  3.28 1.11 5.05 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.24 1.765 0.36 ;
      RECT  1.615 0.36 1.765 0.44 ;
      RECT  0.08 0.36 0.19 0.46 ;
      RECT  1.615 0.44 2.85 0.56 ;
      RECT  2.71 0.775 4.56 0.905 ;
      RECT  2.71 0.905 2.84 1.235 ;
      RECT  0.3 0.45 1.515 0.56 ;
      RECT  1.365 0.56 1.515 1.235 ;
      RECT  1.365 1.235 2.84 1.24 ;
      RECT  0.07 1.24 2.84 1.365 ;
      RECT  0.07 1.365 0.19 1.46 ;
  END
END SEN_AN2_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_1P5
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_1P5
  CLASS CORE ;
  FOREIGN SEN_AN2_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0699 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.75 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0699 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.37 1.41 0.5 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.025 1.41 1.155 1.75 ;
      RECT  1.605 1.41 1.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.605 0.05 1.735 0.39 ;
      RECT  1.025 0.05 1.145 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.345 0.27 1.46 0.51 ;
      RECT  1.345 0.51 1.65 0.69 ;
      RECT  1.55 0.69 1.65 1.11 ;
      RECT  1.345 1.11 1.65 1.29 ;
      RECT  1.345 1.29 1.455 1.53 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.205 0.81 0.31 ;
      RECT  0.065 0.31 0.185 0.425 ;
      RECT  1.15 0.785 1.44 0.895 ;
      RECT  1.15 0.895 1.25 1.21 ;
      RECT  0.305 0.4 0.65 0.505 ;
      RECT  0.55 0.505 0.65 1.21 ;
      RECT  0.07 1.21 1.25 1.3 ;
      RECT  0.07 1.3 0.19 1.43 ;
      RECT  0.7 1.3 0.82 1.56 ;
  END
END SEN_AN2_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN2_5
#      Description : "2-Input AND"
#      Equation    : X=A1&A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN2_5
  CLASS CORE ;
  FOREIGN SEN_AN2_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 0.9 ;
      RECT  0.15 0.9 0.855 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2319 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.7 2.25 0.9 ;
      RECT  1.55 0.9 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2319 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.2 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.59 1.41 0.72 1.75 ;
      RECT  1.11 1.41 1.24 1.75 ;
      RECT  1.37 1.41 1.5 1.75 ;
      RECT  1.89 1.41 2.02 1.75 ;
      RECT  2.41 1.41 2.54 1.75 ;
      RECT  2.93 1.41 3.06 1.75 ;
      RECT  3.45 1.41 3.58 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  1.37 0.05 1.5 0.39 ;
      RECT  1.89 0.05 2.02 0.39 ;
      RECT  2.93 0.05 3.06 0.39 ;
      RECT  3.45 0.05 3.58 0.39 ;
      RECT  2.415 0.05 2.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.675 0.5 3.85 0.7 ;
      RECT  3.55 0.7 3.65 1.1 ;
      RECT  2.675 1.1 3.85 1.3 ;
    END
    ANTENNADIFFAREA 0.605 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.24 1.235 0.36 ;
      RECT  0.075 0.36 0.195 0.46 ;
      RECT  1.13 0.36 1.235 0.48 ;
      RECT  1.13 0.48 2.3 0.6 ;
      RECT  2.35 0.79 3.44 0.9 ;
      RECT  2.35 0.9 2.46 1.19 ;
      RECT  0.31 0.45 1.04 0.57 ;
      RECT  0.95 0.57 1.04 1.19 ;
      RECT  0.305 1.19 2.46 1.31 ;
  END
END SEN_AN2_5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_0P5
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_0P5
  CLASS CORE ;
  FOREIGN SEN_AN3_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0201 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0201 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.5 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0201 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.355 1.41 0.485 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.875 1.41 1.005 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.86 0.05 0.99 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.21 1.25 1.53 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.1 0.17 0.22 0.27 ;
      RECT  0.1 0.27 0.43 0.39 ;
      RECT  0.34 0.39 0.43 1.21 ;
      RECT  0.1 1.21 1.06 1.3 ;
      RECT  0.97 0.76 1.06 1.21 ;
      RECT  0.1 1.3 0.22 1.63 ;
      RECT  0.62 1.3 0.74 1.63 ;
  END
END SEN_AN3_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_1
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_1
  CLASS CORE ;
  FOREIGN SEN_AN3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0516 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.92 ;
      RECT  0.52 0.92 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0516 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.145 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0516 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.44 0.46 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.91 1.43 1.03 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.815 0.05 0.985 0.355 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.47 1.305 1.49 ;
    END
    ANTENNADIFFAREA 0.218 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.18 0.185 0.31 ;
      RECT  0.065 0.31 0.43 0.4 ;
      RECT  0.34 0.4 0.43 1.24 ;
      RECT  0.065 1.24 1.06 1.34 ;
      RECT  0.97 0.755 1.06 1.24 ;
      RECT  0.065 1.34 0.185 1.47 ;
  END
END SEN_AN3_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_2
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_2
  CLASS CORE ;
  FOREIGN SEN_AN3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1032 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.915 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1032 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.685 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1032 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.23 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.56 1.48 0.735 1.75 ;
      RECT  1.09 1.44 1.27 1.75 ;
      RECT  1.71 1.445 1.89 1.75 ;
      RECT  2.415 1.21 2.555 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.265 0.05 1.435 0.26 ;
      RECT  1.85 0.05 2.01 0.59 ;
      RECT  2.415 0.05 2.555 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.31 2.27 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.06 0.16 0.705 0.25 ;
      RECT  0.06 0.25 0.19 0.39 ;
      RECT  0.58 0.25 0.705 0.53 ;
      RECT  0.58 0.53 1.25 0.62 ;
      RECT  1.08 0.62 1.25 0.64 ;
      RECT  0.82 0.35 1.735 0.44 ;
      RECT  0.34 0.35 0.45 1.24 ;
      RECT  0.34 1.24 2.06 1.35 ;
      RECT  1.965 0.71 2.06 1.24 ;
      RECT  0.34 1.35 0.45 1.385 ;
  END
END SEN_AN3_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_4
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_4
  CLASS CORE ;
  FOREIGN SEN_AN3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.925 ;
      RECT  0.35 0.925 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2064 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.885 ;
      RECT  1.35 0.885 1.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2064 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.925 ;
      RECT  2.95 0.925 3.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2064 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.435 0.45 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.84 1.435 0.97 1.75 ;
      RECT  1.36 1.435 1.49 1.75 ;
      RECT  1.93 1.435 2.06 1.75 ;
      RECT  2.595 1.435 2.725 1.75 ;
      RECT  3.17 1.435 3.3 1.75 ;
      RECT  3.69 1.41 3.82 1.75 ;
      RECT  4.215 1.21 4.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  3.69 0.05 3.82 0.36 ;
      RECT  2.13 0.05 2.26 0.39 ;
      RECT  2.65 0.05 2.78 0.39 ;
      RECT  3.17 0.05 3.3 0.39 ;
      RECT  4.215 0.05 4.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 4.07 0.69 ;
      RECT  3.95 0.69 4.07 1.11 ;
      RECT  3.435 1.11 4.07 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.22 1.81 0.34 ;
      RECT  0.065 0.34 0.19 0.395 ;
      RECT  1.31 0.48 3.09 0.595 ;
      RECT  3.2 0.78 3.84 0.895 ;
      RECT  3.2 0.895 3.31 1.21 ;
      RECT  0.27 0.48 1.05 0.59 ;
      RECT  0.96 0.59 1.05 1.21 ;
      RECT  0.06 1.21 3.31 1.34 ;
      RECT  0.06 1.34 0.19 1.44 ;
  END
END SEN_AN3_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_16
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_16
  CLASS CORE ;
  FOREIGN SEN_AN3_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.75 0.47 11.85 1.025 ;
      RECT  10.15 0.47 10.25 1.025 ;
      RECT  8.55 0.48 8.65 1.02 ;
      RECT  6.95 0.48 7.05 1.02 ;
      RECT  5.55 0.47 5.65 1.025 ;
      RECT  3.95 0.47 4.05 1.065 ;
      RECT  2.35 0.47 2.45 1.025 ;
      RECT  0.75 0.51 0.85 1.05 ;
      LAYER M2 ;
      RECT  0.71 0.55 11.89 0.65 ;
      LAYER V1 ;
      RECT  11.75 0.55 11.85 0.65 ;
      RECT  10.15 0.55 10.25 0.65 ;
      RECT  8.55 0.55 8.65 0.65 ;
      RECT  6.95 0.55 7.05 0.65 ;
      RECT  5.55 0.55 5.65 0.65 ;
      RECT  3.95 0.55 4.05 0.65 ;
      RECT  2.35 0.55 2.45 0.65 ;
      RECT  0.75 0.55 0.85 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8535 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.95 0.71 12.25 0.985 ;
      RECT  11.35 0.67 11.45 1.09 ;
      RECT  10.55 0.71 10.85 0.985 ;
      RECT  9.75 0.71 10.05 0.985 ;
      RECT  8.95 0.71 9.25 0.985 ;
      RECT  8.155 0.71 8.455 0.985 ;
      RECT  7.35 0.71 7.65 0.985 ;
      RECT  6.55 0.71 6.85 0.985 ;
      RECT  5.75 0.71 6.05 0.985 ;
      RECT  4.95 0.71 5.25 0.985 ;
      RECT  4.35 0.71 4.65 0.985 ;
      RECT  3.55 0.71 3.85 0.985 ;
      RECT  2.75 0.71 3.05 0.985 ;
      RECT  1.95 0.71 2.25 0.985 ;
      RECT  1.15 0.71 1.45 0.985 ;
      RECT  0.35 0.71 0.65 0.985 ;
      LAYER M2 ;
      RECT  0.31 0.75 12.29 0.85 ;
      LAYER V1 ;
      RECT  11.95 0.75 12.05 0.85 ;
      RECT  12.15 0.75 12.25 0.85 ;
      RECT  11.35 0.75 11.45 0.85 ;
      RECT  10.55 0.75 10.65 0.85 ;
      RECT  10.75 0.75 10.85 0.85 ;
      RECT  9.75 0.75 9.85 0.85 ;
      RECT  9.95 0.75 10.05 0.85 ;
      RECT  8.95 0.75 9.05 0.85 ;
      RECT  9.15 0.75 9.25 0.85 ;
      RECT  8.155 0.75 8.255 0.85 ;
      RECT  8.355 0.75 8.455 0.85 ;
      RECT  7.35 0.75 7.45 0.85 ;
      RECT  7.55 0.75 7.65 0.85 ;
      RECT  6.55 0.75 6.65 0.85 ;
      RECT  6.75 0.75 6.85 0.85 ;
      RECT  5.75 0.75 5.85 0.85 ;
      RECT  5.95 0.75 6.05 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
      RECT  5.15 0.75 5.25 0.85 ;
      RECT  4.35 0.75 4.45 0.85 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
      RECT  0.35 0.75 0.45 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8535 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.35 0.71 12.47 1.09 ;
      RECT  10.95 0.91 11.25 1.09 ;
      RECT  9.35 0.88 9.65 1.09 ;
      RECT  7.75 0.885 8.05 1.09 ;
      RECT  6.15 0.885 6.45 1.09 ;
      RECT  4.75 0.675 4.85 1.1 ;
      RECT  3.15 0.885 3.45 1.09 ;
      RECT  1.55 0.885 1.85 1.09 ;
      RECT  0.15 0.675 0.25 1.095 ;
      LAYER M2 ;
      RECT  0.11 0.95 12.49 1.05 ;
      LAYER V1 ;
      RECT  12.35 0.95 12.45 1.05 ;
      RECT  10.95 0.95 11.05 1.05 ;
      RECT  11.15 0.95 11.25 1.05 ;
      RECT  9.35 0.95 9.45 1.05 ;
      RECT  9.55 0.95 9.65 1.05 ;
      RECT  7.75 0.95 7.85 1.05 ;
      RECT  7.95 0.95 8.05 1.05 ;
      RECT  6.15 0.95 6.25 1.05 ;
      RECT  6.35 0.95 6.45 1.05 ;
      RECT  4.75 0.95 4.85 1.05 ;
      RECT  3.15 0.95 3.25 1.05 ;
      RECT  3.35 0.95 3.45 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  1.75 0.95 1.85 1.05 ;
      RECT  0.15 0.95 0.25 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8535 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 17.0 1.85 ;
      RECT  0.56 1.45 0.73 1.75 ;
      RECT  1.08 1.45 1.25 1.75 ;
      RECT  1.6 1.45 1.77 1.75 ;
      RECT  2.12 1.45 2.29 1.75 ;
      RECT  2.64 1.45 2.81 1.75 ;
      RECT  3.16 1.45 3.33 1.75 ;
      RECT  3.68 1.45 3.85 1.75 ;
      RECT  4.2 1.45 4.37 1.75 ;
      RECT  4.72 1.45 4.89 1.75 ;
      RECT  5.24 1.45 5.41 1.75 ;
      RECT  5.76 1.45 5.93 1.75 ;
      RECT  6.28 1.45 6.45 1.75 ;
      RECT  6.8 1.45 6.97 1.75 ;
      RECT  7.32 1.45 7.49 1.75 ;
      RECT  7.84 1.45 8.01 1.75 ;
      RECT  8.36 1.45 8.53 1.75 ;
      RECT  8.88 1.45 9.05 1.75 ;
      RECT  9.4 1.45 9.57 1.75 ;
      RECT  9.92 1.45 10.09 1.75 ;
      RECT  10.44 1.45 10.61 1.75 ;
      RECT  10.96 1.45 11.13 1.75 ;
      RECT  11.48 1.45 11.65 1.75 ;
      RECT  12.0 1.45 12.17 1.75 ;
      RECT  12.52 1.45 12.69 1.75 ;
      RECT  13.06 1.39 13.19 1.75 ;
      RECT  13.58 1.39 13.71 1.75 ;
      RECT  14.1 1.39 14.23 1.75 ;
      RECT  14.62 1.39 14.75 1.75 ;
      RECT  15.14 1.39 15.27 1.75 ;
      RECT  15.66 1.39 15.79 1.75 ;
      RECT  16.195 1.39 16.325 1.75 ;
      RECT  16.76 1.21 16.88 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 17.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
      RECT  14.65 1.75 14.75 1.85 ;
      RECT  15.25 1.75 15.35 1.85 ;
      RECT  15.85 1.75 15.95 1.85 ;
      RECT  16.45 1.75 16.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 17.0 0.05 ;
      RECT  13.06 0.05 13.19 0.36 ;
      RECT  13.58 0.05 13.71 0.36 ;
      RECT  14.1 0.05 14.23 0.36 ;
      RECT  14.62 0.05 14.75 0.36 ;
      RECT  10.98 0.05 11.11 0.37 ;
      RECT  3.18 0.05 3.31 0.385 ;
      RECT  4.74 0.05 4.87 0.385 ;
      RECT  6.3 0.05 6.43 0.385 ;
      RECT  7.86 0.05 7.99 0.385 ;
      RECT  9.42 0.05 9.55 0.385 ;
      RECT  12.54 0.05 12.67 0.385 ;
      RECT  15.14 0.05 15.27 0.39 ;
      RECT  15.66 0.05 15.79 0.39 ;
      RECT  16.195 0.05 16.325 0.39 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  1.625 0.05 1.745 0.59 ;
      RECT  16.76 0.05 16.88 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 17.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
      RECT  14.65 -0.05 14.75 0.05 ;
      RECT  15.25 -0.05 15.35 0.05 ;
      RECT  15.85 -0.05 15.95 0.05 ;
      RECT  16.45 -0.05 16.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  12.78 0.45 15.05 0.51 ;
      RECT  12.78 0.51 16.65 0.61 ;
      RECT  14.74 0.61 16.65 0.69 ;
      RECT  14.74 0.69 15.06 1.11 ;
      RECT  12.805 1.11 16.65 1.29 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  11.54 0.235 12.265 0.36 ;
      RECT  11.54 0.36 11.66 0.46 ;
      RECT  12.14 0.36 12.265 0.495 ;
      RECT  9.75 0.24 10.45 0.36 ;
      RECT  10.35 0.36 10.45 0.46 ;
      RECT  9.75 0.36 9.85 0.475 ;
      RECT  10.35 0.46 11.66 0.575 ;
      RECT  8.15 0.24 8.85 0.36 ;
      RECT  8.75 0.36 8.85 0.475 ;
      RECT  8.15 0.36 8.25 0.485 ;
      RECT  8.75 0.475 9.85 0.575 ;
      RECT  6.55 0.24 7.25 0.36 ;
      RECT  6.55 0.36 6.65 0.485 ;
      RECT  7.15 0.36 7.25 0.485 ;
      RECT  5.35 0.24 6.05 0.36 ;
      RECT  5.35 0.36 5.45 0.485 ;
      RECT  5.95 0.36 6.05 0.485 ;
      RECT  3.55 0.24 4.25 0.36 ;
      RECT  3.55 0.36 3.65 0.485 ;
      RECT  4.15 0.36 4.25 0.485 ;
      RECT  2.35 0.24 2.65 0.36 ;
      RECT  2.55 0.36 2.65 0.485 ;
      RECT  2.55 0.485 3.65 0.585 ;
      RECT  4.15 0.485 5.45 0.585 ;
      RECT  5.95 0.485 6.65 0.585 ;
      RECT  7.15 0.485 8.25 0.585 ;
      RECT  12.14 0.495 12.685 0.62 ;
      RECT  8.75 0.575 8.85 1.18 ;
      RECT  10.35 0.575 10.45 1.18 ;
      RECT  11.54 0.575 11.66 1.18 ;
      RECT  2.55 0.585 2.65 1.18 ;
      RECT  5.35 0.585 5.45 1.18 ;
      RECT  4.15 0.585 4.25 1.19 ;
      RECT  7.15 0.585 7.25 1.18 ;
      RECT  12.56 0.62 12.685 0.72 ;
      RECT  12.56 0.72 14.6 0.97 ;
      RECT  12.56 0.97 12.685 1.18 ;
      RECT  0.79 0.24 1.05 0.36 ;
      RECT  0.95 0.36 1.05 1.18 ;
      RECT  0.95 1.18 2.65 1.19 ;
      RECT  5.35 1.18 12.685 1.19 ;
      RECT  0.95 1.19 3.03 1.195 ;
      RECT  3.46 1.19 12.685 1.195 ;
      RECT  0.95 1.195 12.685 1.24 ;
      RECT  0.3 1.24 12.685 1.36 ;
  END
END SEN_AN3_16
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_S_1
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_S_1
  CLASS CORE ;
  FOREIGN SEN_AN3_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0408 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.31 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0408 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0408 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.885 1.41 1.015 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.94 0.05 1.06 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.305 0.6 ;
      RECT  1.15 0.6 1.34 0.69 ;
      RECT  1.24 0.69 1.34 1.11 ;
      RECT  1.15 1.11 1.34 1.2 ;
      RECT  1.15 1.2 1.305 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.955 0.795 1.15 0.885 ;
      RECT  0.955 0.885 1.045 1.23 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 1.23 ;
      RECT  0.065 1.23 1.045 1.32 ;
      RECT  0.065 1.32 0.185 1.59 ;
      RECT  0.585 1.32 0.705 1.59 ;
  END
END SEN_AN3_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_S_2
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_S_2
  CLASS CORE ;
  FOREIGN SEN_AN3_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0774 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.7 1.05 1.13 ;
      RECT  0.85 1.13 1.05 1.22 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0774 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.45 1.21 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0774 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.41 0.205 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.58 1.49 0.75 1.75 ;
      RECT  1.1 1.49 1.27 1.75 ;
      RECT  1.62 1.49 1.79 1.75 ;
      RECT  2.185 1.21 2.305 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.13 0.05 1.26 0.355 ;
      RECT  1.645 0.05 1.765 0.59 ;
      RECT  2.185 0.05 2.305 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.92 0.31 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.085 0.17 0.725 0.28 ;
      RECT  0.085 0.28 0.205 0.39 ;
      RECT  0.605 0.28 0.725 0.39 ;
      RECT  0.825 0.445 1.54 0.555 ;
      RECT  0.36 0.41 0.45 1.31 ;
      RECT  0.36 1.31 1.83 1.4 ;
      RECT  1.73 0.725 1.83 1.31 ;
      RECT  0.36 1.4 0.465 1.595 ;
      RECT  0.865 1.4 0.985 1.595 ;
      RECT  1.385 1.4 1.505 1.595 ;
  END
END SEN_AN3_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_S_4
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_S_4
  CLASS CORE ;
  FOREIGN SEN_AN3_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 0.715 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1392 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 0.91 ;
      RECT  1.15 0.91 1.65 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1392 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.35 0.915 ;
      RECT  1.95 0.915 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1392 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.58 1.435 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  1.62 1.44 1.75 1.75 ;
      RECT  1.85 1.44 1.98 1.75 ;
      RECT  2.37 1.435 2.5 1.75 ;
      RECT  2.89 1.39 3.02 1.75 ;
      RECT  3.415 1.21 3.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  2.89 0.05 3.02 0.365 ;
      RECT  1.85 0.05 1.98 0.38 ;
      RECT  2.375 0.05 2.495 0.59 ;
      RECT  3.415 0.05 3.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.61 0.455 3.3 0.575 ;
      RECT  3.15 0.575 3.25 1.11 ;
      RECT  2.65 1.11 3.275 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 0.245 1.535 0.355 ;
      RECT  1.055 0.475 2.26 0.595 ;
      RECT  2.47 0.79 3.06 0.89 ;
      RECT  2.47 0.89 2.56 1.245 ;
      RECT  0.065 0.345 0.185 0.445 ;
      RECT  0.065 0.445 0.935 0.565 ;
      RECT  0.845 0.565 0.935 1.245 ;
      RECT  0.845 1.245 2.56 1.255 ;
      RECT  0.325 1.255 2.56 1.345 ;
      RECT  0.845 1.345 0.965 1.53 ;
      RECT  0.325 1.345 0.445 1.55 ;
      RECT  1.365 1.345 1.485 1.55 ;
  END
END SEN_AN3_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_S_8
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_S_8
  CLASS CORE ;
  FOREIGN SEN_AN3_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 0.98 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2754 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.91 ;
      RECT  1.75 0.91 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2754 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 3.65 0.91 ;
      RECT  2.95 0.91 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2754 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.43 0.45 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.84 1.43 0.97 1.75 ;
      RECT  1.36 1.43 1.49 1.75 ;
      RECT  1.88 1.43 2.01 1.75 ;
      RECT  2.4 1.43 2.53 1.75 ;
      RECT  2.92 1.43 3.05 1.75 ;
      RECT  3.44 1.43 3.57 1.75 ;
      RECT  3.965 1.21 4.085 1.75 ;
      RECT  4.48 1.415 4.61 1.75 ;
      RECT  5.0 1.415 5.13 1.75 ;
      RECT  5.52 1.415 5.65 1.75 ;
      RECT  6.08 1.21 6.2 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  4.48 0.05 4.61 0.365 ;
      RECT  5.0 0.05 5.13 0.365 ;
      RECT  5.52 0.05 5.65 0.365 ;
      RECT  2.92 0.05 3.05 0.385 ;
      RECT  3.44 0.05 3.57 0.385 ;
      RECT  3.965 0.05 4.085 0.59 ;
      RECT  6.08 0.05 6.2 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.2 0.455 5.96 0.575 ;
      RECT  4.2 0.575 5.65 0.585 ;
      RECT  5.48 0.585 5.65 1.11 ;
      RECT  4.225 1.11 5.905 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 0.24 2.575 0.36 ;
      RECT  1.575 0.475 3.875 0.595 ;
      RECT  3.745 0.775 5.39 0.905 ;
      RECT  3.745 0.905 3.875 1.21 ;
      RECT  0.065 0.345 0.185 0.455 ;
      RECT  0.065 0.455 1.25 0.575 ;
      RECT  1.12 0.575 1.25 1.21 ;
      RECT  1.12 1.21 3.875 1.25 ;
      RECT  0.065 1.25 3.875 1.34 ;
      RECT  0.585 1.34 0.705 1.49 ;
      RECT  1.105 1.34 1.225 1.49 ;
      RECT  1.625 1.34 1.745 1.49 ;
      RECT  2.145 1.34 2.265 1.49 ;
      RECT  3.705 1.34 3.875 1.49 ;
      RECT  0.065 1.34 0.185 1.5 ;
      RECT  2.665 1.34 2.785 1.5 ;
      RECT  3.185 1.34 3.305 1.5 ;
  END
END SEN_AN3_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3_8
#      Description : "3-Input AND"
#      Equation    : X=A1&A2&A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3_8
  CLASS CORE ;
  FOREIGN SEN_AN3_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  0.55 0.91 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4266 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.45 0.91 ;
      RECT  2.55 0.91 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4266 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.05 0.91 ;
      RECT  4.15 0.91 5.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4266 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.455 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.845 1.44 0.975 1.75 ;
      RECT  1.365 1.44 1.495 1.75 ;
      RECT  1.885 1.44 2.015 1.75 ;
      RECT  2.405 1.44 2.535 1.75 ;
      RECT  2.925 1.44 3.055 1.75 ;
      RECT  3.445 1.44 3.575 1.75 ;
      RECT  3.965 1.44 4.095 1.75 ;
      RECT  4.485 1.44 4.615 1.75 ;
      RECT  5.005 1.44 5.135 1.75 ;
      RECT  5.53 1.21 5.65 1.75 ;
      RECT  6.045 1.415 6.175 1.75 ;
      RECT  6.565 1.41 6.695 1.75 ;
      RECT  7.085 1.41 7.215 1.75 ;
      RECT  7.61 1.21 7.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  3.965 0.05 4.095 0.36 ;
      RECT  4.485 0.05 4.615 0.39 ;
      RECT  5.005 0.05 5.135 0.39 ;
      RECT  6.045 0.05 6.175 0.39 ;
      RECT  6.565 0.05 6.695 0.39 ;
      RECT  7.085 0.05 7.215 0.39 ;
      RECT  5.53 0.05 5.65 0.59 ;
      RECT  7.61 0.05 7.73 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.765 0.485 7.46 0.615 ;
      RECT  7.29 0.615 7.46 1.11 ;
      RECT  5.75 1.11 7.46 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.68 0.19 2.24 0.23 ;
      RECT  0.305 0.23 3.62 0.36 ;
      RECT  3.16 0.45 4.375 0.5 ;
      RECT  2.1 0.5 5.415 0.62 ;
      RECT  5.245 0.76 7.095 0.93 ;
      RECT  5.245 0.93 5.415 1.18 ;
      RECT  0.07 0.37 0.19 0.47 ;
      RECT  0.07 0.47 1.775 0.59 ;
      RECT  1.605 0.59 1.775 1.18 ;
      RECT  1.605 1.18 5.415 1.22 ;
      RECT  0.07 1.22 5.415 1.35 ;
      RECT  0.07 1.35 0.19 1.44 ;
  END
END SEN_AN3_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3B_0P5
#      Description : "3-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3B_0P5
  CLASS CORE ;
  FOREIGN SEN_AN3B_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.655 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.115 1.41 0.245 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.655 1.41 0.785 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.655 0.05 0.785 0.39 ;
      RECT  1.2 0.05 1.32 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.21 1.05 0.51 ;
      RECT  0.95 0.51 1.35 0.69 ;
      RECT  1.25 0.69 1.35 1.11 ;
      RECT  1.15 1.11 1.35 1.2 ;
      RECT  1.15 1.2 1.255 1.53 ;
    END
    ANTENNADIFFAREA 0.1 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.955 0.79 1.16 0.905 ;
      RECT  0.955 0.905 1.045 1.21 ;
      RECT  0.08 0.225 0.46 0.345 ;
      RECT  0.37 0.345 0.46 1.21 ;
      RECT  0.37 1.21 1.045 1.3 ;
      RECT  0.37 1.3 0.515 1.61 ;
  END
END SEN_AN3B_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3B_1
#      Description : "3-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3B_1
  CLASS CORE ;
  FOREIGN SEN_AN3B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0444 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.655 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0444 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.12 1.44 0.24 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.665 1.42 0.785 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.665 0.05 0.785 0.375 ;
      RECT  1.2 0.05 1.32 0.43 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.3 1.05 0.6 ;
      RECT  0.95 0.6 1.35 0.69 ;
      RECT  1.25 0.69 1.35 1.11 ;
      RECT  1.15 1.11 1.35 1.2 ;
      RECT  1.15 1.2 1.275 1.5 ;
    END
    ANTENNADIFFAREA 0.19 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.955 0.8 1.16 0.89 ;
      RECT  0.955 0.89 1.045 1.24 ;
      RECT  0.08 0.25 0.46 0.34 ;
      RECT  0.37 0.34 0.46 1.24 ;
      RECT  0.37 1.24 1.045 1.33 ;
      RECT  0.37 1.33 0.5 1.6 ;
  END
END SEN_AN3B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3B_2
#      Description : "3-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3B_2
  CLASS CORE ;
  FOREIGN SEN_AN3B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.4 0.185 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.59 1.44 0.71 1.75 ;
      RECT  1.11 1.44 1.23 1.75 ;
      RECT  1.605 1.495 1.775 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.85 0.05 0.97 0.345 ;
      RECT  1.36 0.05 1.48 0.38 ;
      RECT  1.89 0.05 2.01 0.385 ;
      RECT  2.415 0.05 2.535 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.59 0.475 2.45 0.595 ;
      RECT  2.35 0.595 2.45 1.11 ;
      RECT  1.87 1.11 2.535 1.21 ;
      RECT  2.15 1.21 2.535 1.29 ;
    END
    ANTENNADIFFAREA 0.38 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.215 0.71 0.305 ;
      RECT  0.59 0.305 0.71 0.435 ;
      RECT  0.065 0.305 0.19 0.45 ;
      RECT  0.59 0.435 1.255 0.56 ;
      RECT  1.555 0.79 2.26 0.88 ;
      RECT  1.555 0.88 1.645 1.05 ;
      RECT  1.14 1.05 1.645 1.14 ;
      RECT  1.14 1.14 1.23 1.23 ;
      RECT  0.34 0.415 0.445 0.585 ;
      RECT  0.34 0.585 0.43 1.23 ;
      RECT  0.34 1.23 1.23 1.35 ;
      RECT  0.34 1.35 0.45 1.44 ;
      RECT  1.345 1.3 2.0 1.38 ;
      RECT  1.345 1.38 2.3 1.405 ;
      RECT  1.91 1.405 2.3 1.5 ;
  END
END SEN_AN3B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3B_4
#      Description : "3-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3B_4
  CLASS CORE ;
  FOREIGN SEN_AN3B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.85 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1779 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1779 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.23 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.585 1.435 0.705 1.75 ;
      RECT  1.105 1.435 1.225 1.75 ;
      RECT  1.625 1.435 1.745 1.75 ;
      RECT  3.2 1.44 3.32 1.75 ;
      RECT  3.72 1.44 3.84 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.585 0.05 0.705 0.345 ;
      RECT  2.395 0.05 2.515 0.365 ;
      RECT  2.925 0.05 3.045 0.365 ;
      RECT  3.46 0.05 3.58 0.365 ;
      RECT  3.98 0.05 4.1 0.575 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  1.875 0.05 1.995 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.455 3.865 0.51 ;
      RECT  2.11 0.51 3.865 0.585 ;
      RECT  2.11 0.585 2.85 0.69 ;
      RECT  2.75 0.69 2.85 1.11 ;
      RECT  1.95 1.11 2.85 1.29 ;
    END
    ANTENNADIFFAREA 0.616 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.24 1.54 0.36 ;
      RECT  0.845 0.36 0.965 0.44 ;
      RECT  0.29 0.44 0.965 0.56 ;
      RECT  1.08 0.45 1.775 0.57 ;
      RECT  1.685 0.57 1.775 0.785 ;
      RECT  1.685 0.785 2.66 0.875 ;
      RECT  1.685 0.875 1.775 1.225 ;
      RECT  0.285 1.225 1.775 1.345 ;
      RECT  2.94 1.22 4.1 1.34 ;
      RECT  2.94 1.34 3.06 1.43 ;
      RECT  3.98 1.34 4.1 1.44 ;
      RECT  1.845 1.43 3.06 1.55 ;
  END
END SEN_AN3B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN3B_8
#      Description : "3-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN3B_8
  CLASS CORE ;
  FOREIGN SEN_AN3B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.05 0.89 ;
      RECT  5.95 0.89 6.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.234 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  0.585 1.42 0.715 1.75 ;
      RECT  1.105 1.42 1.235 1.75 ;
      RECT  1.625 1.42 1.755 1.75 ;
      RECT  2.145 1.42 2.275 1.75 ;
      RECT  4.735 1.43 4.865 1.75 ;
      RECT  5.255 1.43 5.385 1.75 ;
      RECT  5.775 1.43 5.905 1.75 ;
      RECT  6.295 1.43 6.425 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  2.915 0.05 3.045 0.365 ;
      RECT  3.435 0.05 3.565 0.365 ;
      RECT  3.955 0.05 4.085 0.365 ;
      RECT  4.475 0.05 4.605 0.365 ;
      RECT  4.995 0.05 5.125 0.365 ;
      RECT  5.515 0.05 5.645 0.365 ;
      RECT  6.035 0.05 6.165 0.365 ;
      RECT  0.325 0.05 0.455 0.38 ;
      RECT  0.845 0.05 0.975 0.38 ;
      RECT  2.4 0.05 2.52 0.59 ;
      RECT  6.58 0.05 6.7 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.635 0.455 6.47 0.585 ;
      RECT  4.15 0.585 4.86 0.69 ;
      RECT  4.15 0.69 4.325 1.11 ;
      RECT  2.55 1.11 4.325 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.11 0.24 2.295 0.36 ;
      RECT  1.11 0.36 1.23 0.47 ;
      RECT  0.07 0.37 0.19 0.47 ;
      RECT  0.07 0.47 1.23 0.59 ;
      RECT  1.345 0.46 2.245 0.58 ;
      RECT  2.155 0.58 2.245 0.785 ;
      RECT  2.155 0.785 3.91 0.895 ;
      RECT  2.155 0.895 2.245 1.21 ;
      RECT  0.28 1.21 2.245 1.33 ;
      RECT  4.455 1.21 6.72 1.34 ;
      RECT  4.455 1.34 4.625 1.395 ;
      RECT  3.92 1.395 4.625 1.435 ;
      RECT  2.365 1.435 4.625 1.545 ;
  END
END SEN_AN3B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_0P5
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_0P5
  CLASS CORE ;
  FOREIGN SEN_AN4_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0219 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0219 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.185 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0219 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.53 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0219 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.34 1.455 0.46 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.85 1.455 0.98 1.75 ;
      RECT  1.39 1.41 1.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.33 0.05 0.46 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.085 0.21 0.185 0.75 ;
      RECT  0.085 0.75 0.25 0.84 ;
      RECT  0.15 0.84 0.25 1.37 ;
      RECT  0.075 1.37 0.25 1.59 ;
    END
    ANTENNADIFFAREA 0.089 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.145 0.24 1.52 0.36 ;
      RECT  1.145 0.36 1.255 1.275 ;
      RECT  0.275 0.49 0.44 0.66 ;
      RECT  0.34 0.66 0.44 1.275 ;
      RECT  0.34 1.275 1.255 1.365 ;
      RECT  0.595 1.365 0.715 1.63 ;
      RECT  1.12 1.365 1.255 1.63 ;
  END
END SEN_AN4_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_1
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_1
  CLASS CORE ;
  FOREIGN SEN_AN4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.31 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0546 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.14 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0546 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.91 ;
      RECT  0.75 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0546 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.66 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0546 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.455 0.48 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.99 1.455 1.11 1.75 ;
      RECT  1.56 1.415 1.68 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.365 0.05 0.485 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.07 0.3 0.25 0.5 ;
      RECT  0.15 0.5 0.25 1.3 ;
      RECT  0.07 1.3 0.25 1.5 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.35 0.24 1.685 0.36 ;
      RECT  1.35 0.36 1.45 1.235 ;
      RECT  0.34 0.75 0.44 1.235 ;
      RECT  0.34 1.235 1.45 1.36 ;
  END
END SEN_AN4_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_1P5
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_1P5
  CLASS CORE ;
  FOREIGN SEN_AN4_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.5 1.45 1.18 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.075 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.415 1.48 0.585 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.065 1.48 1.235 1.75 ;
      RECT  1.64 1.48 1.82 1.75 ;
      RECT  2.2 1.21 2.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  1.66 0.05 1.78 0.58 ;
      RECT  2.2 0.05 2.32 0.58 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.05 1.49 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.54 0.25 0.76 0.35 ;
      RECT  0.54 0.35 0.63 0.5 ;
      RECT  0.075 0.27 0.175 0.5 ;
      RECT  0.075 0.5 0.63 0.59 ;
      RECT  1.55 0.745 1.86 0.855 ;
      RECT  1.55 0.855 1.65 1.28 ;
      RECT  1.165 0.25 1.55 0.35 ;
      RECT  1.165 0.35 1.255 1.28 ;
      RECT  0.08 1.28 1.65 1.38 ;
  END
END SEN_AN4_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_2
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_2
  CLASS CORE ;
  FOREIGN SEN_AN4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.15 0.91 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1092 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 0.91 ;
      RECT  0.75 0.91 1.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1092 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.905 ;
      RECT  1.55 0.905 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1092 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.67 2.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1092 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.175 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.575 1.455 0.695 1.75 ;
      RECT  1.225 1.45 1.345 1.75 ;
      RECT  1.875 1.455 1.995 1.75 ;
      RECT  2.56 1.21 2.68 1.75 ;
      RECT  3.215 1.21 3.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  2.135 0.05 2.255 0.345 ;
      RECT  2.645 0.05 2.765 0.59 ;
      RECT  3.215 0.05 3.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.31 3.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.215 1.24 0.335 ;
      RECT  0.055 0.335 0.175 0.39 ;
      RECT  1.33 0.215 1.995 0.335 ;
      RECT  1.875 0.335 1.995 0.44 ;
      RECT  1.875 0.44 2.54 0.56 ;
      RECT  0.81 0.44 1.765 0.56 ;
      RECT  2.35 0.795 2.86 0.885 ;
      RECT  2.35 0.885 2.44 1.24 ;
      RECT  0.29 0.44 0.65 0.56 ;
      RECT  0.55 0.56 0.65 1.24 ;
      RECT  0.29 1.24 2.44 1.36 ;
  END
END SEN_AN4_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_4
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_4
  CLASS CORE ;
  FOREIGN SEN_AN4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2181 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  1.35 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2181 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  2.15 0.91 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2181 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.7 3.65 0.89 ;
      RECT  3.15 0.89 3.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2181 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.43 0.18 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.575 1.45 0.695 1.75 ;
      RECT  1.14 1.45 1.26 1.75 ;
      RECT  1.705 1.45 1.825 1.75 ;
      RECT  2.225 1.45 2.345 1.75 ;
      RECT  2.745 1.45 2.865 1.75 ;
      RECT  3.465 1.45 3.585 1.75 ;
      RECT  3.985 1.2 4.105 1.75 ;
      RECT  4.505 1.43 4.625 1.75 ;
      RECT  5.025 1.425 5.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.945 0.05 3.065 0.36 ;
      RECT  3.465 0.05 3.585 0.36 ;
      RECT  4.505 0.05 4.625 0.385 ;
      RECT  5.025 0.05 5.145 0.385 ;
      RECT  3.985 0.05 4.105 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.245 0.51 4.875 0.69 ;
      RECT  4.75 0.69 4.875 1.11 ;
      RECT  4.245 1.11 4.875 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.215 1.265 0.335 ;
      RECT  0.055 0.335 0.175 0.385 ;
      RECT  1.145 0.335 1.265 0.445 ;
      RECT  1.145 0.445 1.88 0.56 ;
      RECT  1.42 0.24 2.66 0.355 ;
      RECT  2.17 0.45 3.87 0.56 ;
      RECT  2.74 0.56 2.865 0.84 ;
      RECT  3.78 0.785 4.59 0.895 ;
      RECT  3.78 0.895 3.87 1.24 ;
      RECT  0.29 0.44 1.05 0.56 ;
      RECT  0.96 0.56 1.05 1.24 ;
      RECT  0.29 1.24 3.87 1.36 ;
  END
END SEN_AN4_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_S_1
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_S_1
  CLASS CORE ;
  FOREIGN SEN_AN4_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.31 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.1 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.185 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.66 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.455 0.49 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.94 1.455 1.07 1.75 ;
      RECT  1.51 1.41 1.64 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.36 0.05 0.49 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.075 0.23 0.25 0.45 ;
      RECT  0.15 0.45 0.25 1.35 ;
      RECT  0.075 1.35 0.25 1.57 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.245 0.24 1.66 0.36 ;
      RECT  1.245 0.36 1.355 1.275 ;
      RECT  0.34 0.75 0.44 1.275 ;
      RECT  0.34 1.275 1.355 1.365 ;
      RECT  0.66 1.365 0.78 1.58 ;
      RECT  1.235 1.365 1.355 1.58 ;
  END
END SEN_AN4_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_S_1P5
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_S_1P5
  CLASS CORE ;
  FOREIGN SEN_AN4_S_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.67 1.45 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.46 1.075 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.215 1.48 0.385 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.82 1.48 0.99 1.75 ;
      RECT  1.34 1.48 1.51 1.75 ;
      RECT  1.705 1.455 1.815 1.75 ;
      RECT  2.215 1.215 2.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.3 0.05 0.47 0.33 ;
      RECT  1.68 0.05 1.8 0.37 ;
      RECT  2.215 0.05 2.335 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.065 1.49 ;
    END
    ANTENNADIFFAREA 0.176 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.33 0.185 0.43 ;
      RECT  0.065 0.43 0.73 0.55 ;
      RECT  1.34 0.46 1.64 0.58 ;
      RECT  1.54 0.58 1.64 0.745 ;
      RECT  1.54 0.745 1.86 0.855 ;
      RECT  1.54 0.855 1.64 1.27 ;
      RECT  0.545 1.27 1.64 1.39 ;
  END
END SEN_AN4_S_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_S_2
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_S_2
  CLASS CORE ;
  FOREIGN SEN_AN4_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.91 0.45 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 0.91 ;
      RECT  0.75 0.91 1.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.905 ;
      RECT  1.55 0.905 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.67 2.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.235 1.41 0.365 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  1.235 1.455 1.365 1.75 ;
      RECT  2.165 1.45 2.295 1.75 ;
      RECT  2.64 1.21 2.76 1.75 ;
      RECT  3.215 1.21 3.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  2.135 0.05 2.255 0.345 ;
      RECT  2.645 0.05 2.765 0.59 ;
      RECT  3.215 0.05 3.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.31 3.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.215 1.24 0.335 ;
      RECT  0.055 0.335 0.175 0.4 ;
      RECT  1.33 0.215 1.995 0.335 ;
      RECT  1.875 0.335 1.995 0.44 ;
      RECT  1.875 0.44 2.54 0.56 ;
      RECT  0.81 0.44 1.765 0.56 ;
      RECT  2.38 0.795 2.84 0.885 ;
      RECT  2.38 0.885 2.47 1.24 ;
      RECT  0.29 0.44 0.65 0.56 ;
      RECT  0.55 0.56 0.65 1.24 ;
      RECT  0.55 1.24 2.47 1.36 ;
  END
END SEN_AN4_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_S_4
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_S_4
  CLASS CORE ;
  FOREIGN SEN_AN4_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.25 0.91 ;
      RECT  2.75 0.91 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1572 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.14 0.71 2.25 0.91 ;
      RECT  1.75 0.91 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1572 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.15 0.91 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1572 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.35 0.91 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1572 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.585 1.48 0.755 1.75 ;
      RECT  1.105 1.48 1.275 1.75 ;
      RECT  1.625 1.48 1.795 1.75 ;
      RECT  2.145 1.48 2.315 1.75 ;
      RECT  2.685 1.48 2.855 1.75 ;
      RECT  3.225 1.48 3.395 1.75 ;
      RECT  3.52 1.21 3.64 1.75 ;
      RECT  4.035 1.4 4.165 1.75 ;
      RECT  4.58 1.21 4.7 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.605 0.05 0.735 0.345 ;
      RECT  4.035 0.05 4.165 0.35 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  3.52 0.05 3.64 0.59 ;
      RECT  4.58 0.05 4.7 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.755 0.44 4.47 0.56 ;
      RECT  4.15 0.56 4.25 1.11 ;
      RECT  3.75 1.11 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.08 0.23 1.77 0.35 ;
      RECT  1.65 0.35 1.77 0.44 ;
      RECT  1.65 0.44 2.34 0.56 ;
      RECT  1.86 0.23 3.14 0.35 ;
      RECT  0.325 0.44 1.56 0.56 ;
      RECT  3.34 0.785 4.06 0.895 ;
      RECT  3.34 0.895 3.43 1.3 ;
      RECT  2.55 0.44 3.42 0.56 ;
      RECT  2.55 0.56 2.65 1.3 ;
      RECT  0.34 1.3 3.43 1.39 ;
      RECT  0.34 1.39 0.46 1.54 ;
      RECT  0.87 1.39 0.99 1.54 ;
      RECT  1.39 1.39 1.51 1.54 ;
      RECT  1.91 1.39 2.03 1.54 ;
      RECT  2.44 1.39 2.56 1.54 ;
      RECT  2.97 1.39 3.09 1.54 ;
  END
END SEN_AN4_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_S_8
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_S_8
  CLASS CORE ;
  FOREIGN SEN_AN4_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.05 0.91 ;
      RECT  4.55 0.91 5.23 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3042 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.05 0.91 ;
      RECT  2.95 0.91 4.05 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3042 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 2.85 0.91 ;
      RECT  1.75 0.91 2.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3042 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 1.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3042 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.35 1.49 0.52 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.87 1.49 1.04 1.75 ;
      RECT  1.39 1.49 1.56 1.75 ;
      RECT  1.91 1.49 2.08 1.75 ;
      RECT  2.43 1.49 2.6 1.75 ;
      RECT  2.95 1.49 3.12 1.75 ;
      RECT  3.47 1.49 3.64 1.75 ;
      RECT  3.99 1.49 4.16 1.75 ;
      RECT  4.51 1.49 4.68 1.75 ;
      RECT  5.03 1.49 5.2 1.75 ;
      RECT  5.56 1.21 5.66 1.75 ;
      RECT  6.06 1.41 6.19 1.75 ;
      RECT  6.58 1.41 6.71 1.75 ;
      RECT  7.1 1.41 7.23 1.75 ;
      RECT  7.62 1.41 7.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  6.06 0.05 6.19 0.35 ;
      RECT  6.58 0.05 6.71 0.35 ;
      RECT  7.1 0.05 7.23 0.35 ;
      RECT  0.63 0.05 0.76 0.39 ;
      RECT  1.15 0.05 1.28 0.39 ;
      RECT  7.62 0.05 7.745 0.39 ;
      RECT  0.1 0.05 0.22 0.59 ;
      RECT  5.545 0.05 5.665 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.78 0.44 7.51 0.56 ;
      RECT  5.78 0.56 7.055 0.57 ;
      RECT  6.885 0.57 7.055 1.11 ;
      RECT  5.75 1.11 7.485 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.62 0.195 3.9 0.345 ;
      RECT  4.005 0.195 5.215 0.345 ;
      RECT  4.005 0.345 4.155 0.445 ;
      RECT  2.92 0.445 4.155 0.595 ;
      RECT  0.35 0.52 2.63 0.67 ;
      RECT  5.32 0.77 6.795 0.91 ;
      RECT  5.32 0.91 5.47 1.25 ;
      RECT  5.315 0.2 5.435 0.44 ;
      RECT  4.26 0.44 5.435 0.56 ;
      RECT  4.26 0.56 4.41 1.25 ;
      RECT  4.26 1.25 5.47 1.28 ;
      RECT  0.075 1.28 5.47 1.4 ;
      RECT  5.315 1.4 5.47 1.61 ;
  END
END SEN_AN4_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4_8
#      Description : "4-Input AND"
#      Equation    : X=A1&A2&A3&A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4_8
  CLASS CORE ;
  FOREIGN SEN_AN4_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  0.55 0.91 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4212 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.45 0.91 ;
      RECT  2.55 0.91 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4212 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.25 0.91 ;
      RECT  4.35 0.91 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4212 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.71 6.85 0.91 ;
      RECT  5.95 0.91 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4212 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  1.62 1.44 1.75 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  2.66 1.44 2.79 1.75 ;
      RECT  3.18 1.44 3.31 1.75 ;
      RECT  3.7 1.44 3.83 1.75 ;
      RECT  4.22 1.44 4.35 1.75 ;
      RECT  4.74 1.44 4.87 1.75 ;
      RECT  5.26 1.44 5.39 1.75 ;
      RECT  5.78 1.44 5.91 1.75 ;
      RECT  6.3 1.44 6.43 1.75 ;
      RECT  6.82 1.44 6.95 1.75 ;
      RECT  7.345 1.21 7.46 1.75 ;
      RECT  7.86 1.41 7.99 1.75 ;
      RECT  8.38 1.41 8.51 1.75 ;
      RECT  8.9 1.41 9.03 1.75 ;
      RECT  9.42 1.41 9.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  5.78 0.05 5.91 0.385 ;
      RECT  6.3 0.05 6.43 0.385 ;
      RECT  6.82 0.05 6.95 0.385 ;
      RECT  7.86 0.05 7.99 0.385 ;
      RECT  8.38 0.05 8.51 0.385 ;
      RECT  8.9 0.05 9.03 0.385 ;
      RECT  9.42 0.05 9.545 0.39 ;
      RECT  7.345 0.05 7.465 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.58 0.475 9.34 0.595 ;
      RECT  7.58 0.595 9.05 0.605 ;
      RECT  8.88 0.605 9.05 1.11 ;
      RECT  7.55 1.11 9.45 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.675 0.19 2.235 0.23 ;
      RECT  0.3 0.23 3.62 0.36 ;
      RECT  3.91 0.23 5.67 0.36 ;
      RECT  5.5 0.36 5.67 0.475 ;
      RECT  5.5 0.475 7.23 0.605 ;
      RECT  3.44 0.45 4.095 0.5 ;
      RECT  2.09 0.5 5.41 0.62 ;
      RECT  7.06 0.755 8.775 0.925 ;
      RECT  7.06 0.925 7.23 1.18 ;
      RECT  0.065 0.38 0.185 0.47 ;
      RECT  0.065 0.47 1.77 0.6 ;
      RECT  1.6 0.6 1.77 1.18 ;
      RECT  1.6 1.18 7.23 1.22 ;
      RECT  0.3 1.22 7.23 1.35 ;
  END
END SEN_AN4_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4B_0P5
#      Description : "4-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2&B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4B_0P5
  CLASS CORE ;
  FOREIGN SEN_AN4B_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.525 0.31 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.86 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.415 0.46 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.85 1.415 0.98 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.85 0.05 0.98 0.39 ;
      RECT  1.395 0.05 1.525 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.21 1.25 0.71 ;
      RECT  1.15 0.71 1.52 0.89 ;
      RECT  1.4 0.89 1.52 1.53 ;
    END
    ANTENNADIFFAREA 0.106 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.17 0.195 0.27 ;
      RECT  0.075 0.27 0.43 0.39 ;
      RECT  0.34 0.39 0.43 1.235 ;
      RECT  0.075 1.235 1.31 1.325 ;
      RECT  1.205 0.98 1.31 1.235 ;
      RECT  0.075 1.325 0.195 1.63 ;
      RECT  0.595 1.325 0.715 1.63 ;
  END
END SEN_AN4B_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4B_1
#      Description : "4-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2&B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4B_1
  CLASS CORE ;
  FOREIGN SEN_AN4B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.5 1.05 0.745 ;
      RECT  0.95 0.745 1.08 0.925 ;
      RECT  0.95 0.925 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.83 ;
      RECT  0.52 0.83 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.5 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.45 0.45 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.86 1.45 0.98 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  1.415 0.05 1.535 0.36 ;
      RECT  0.86 0.05 0.98 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.5 ;
      RECT  1.15 0.5 1.525 0.6 ;
      RECT  1.435 0.6 1.525 1.11 ;
      RECT  1.35 1.11 1.525 1.49 ;
    END
    ANTENNADIFFAREA 0.202 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.17 0.75 1.345 0.92 ;
      RECT  1.17 0.92 1.26 1.24 ;
      RECT  0.07 0.17 0.19 0.3 ;
      RECT  0.07 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 1.24 ;
      RECT  0.07 1.24 1.26 1.36 ;
      RECT  0.07 1.36 0.19 1.46 ;
  END
END SEN_AN4B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4B_2
#      Description : "4-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2&B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4B_2
  CLASS CORE ;
  FOREIGN SEN_AN4B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.7 2.85 0.9 ;
      RECT  2.75 0.9 2.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.7 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.7 1.05 0.91 ;
      RECT  0.75 0.91 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.45 0.91 ;
      RECT  1.35 0.91 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.59 1.43 0.71 1.75 ;
      RECT  1.105 1.43 1.235 1.75 ;
      RECT  1.63 1.425 1.75 1.75 ;
      RECT  2.67 1.45 2.79 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  2.41 0.05 2.53 0.35 ;
      RECT  1.36 0.05 1.48 0.37 ;
      RECT  2.96 0.05 3.08 0.59 ;
      RECT  1.89 0.05 2.01 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.3 2.255 0.44 ;
      RECT  2.15 0.44 2.85 0.56 ;
      RECT  2.35 0.56 2.45 1.025 ;
      RECT  2.115 1.025 2.45 1.145 ;
    END
    ANTENNADIFFAREA 0.308 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.24 1.255 0.35 ;
      RECT  0.075 0.35 0.18 0.46 ;
      RECT  0.79 0.46 1.765 0.58 ;
      RECT  1.91 0.78 2.22 0.89 ;
      RECT  1.91 0.89 2.01 1.21 ;
      RECT  0.29 0.44 0.65 0.56 ;
      RECT  0.55 0.56 0.65 1.21 ;
      RECT  0.305 1.21 2.01 1.33 ;
      RECT  2.405 1.24 3.1 1.36 ;
      RECT  2.405 1.36 2.535 1.44 ;
      RECT  1.865 1.44 2.535 1.56 ;
  END
END SEN_AN4B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4B_4
#      Description : "4-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2&B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4B_4
  CLASS CORE ;
  FOREIGN SEN_AN4B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.7 5.25 0.89 ;
      RECT  4.75 0.89 4.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.7 2.85 0.89 ;
      RECT  2.35 0.89 2.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2163 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  1.35 0.91 1.855 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2163 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2163 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.45 0.455 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.895 1.45 1.025 1.75 ;
      RECT  1.48 1.45 1.6 1.75 ;
      RECT  2.025 1.45 2.155 1.75 ;
      RECT  2.55 1.45 2.67 1.75 ;
      RECT  3.045 1.46 3.215 1.75 ;
      RECT  4.625 1.45 4.755 1.75 ;
      RECT  5.15 1.45 5.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.335 0.05 0.455 0.35 ;
      RECT  0.855 0.05 0.975 0.35 ;
      RECT  3.85 0.05 3.97 0.35 ;
      RECT  4.37 0.05 4.49 0.35 ;
      RECT  4.89 0.05 5.01 0.35 ;
      RECT  5.41 0.05 5.53 0.59 ;
      RECT  3.33 0.05 3.45 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.565 0.44 5.3 0.56 ;
      RECT  4.15 0.56 4.255 1.11 ;
      RECT  3.55 1.11 4.255 1.29 ;
    END
    ANTENNADIFFAREA 0.616 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.485 0.24 3.215 0.355 ;
      RECT  0.05 0.445 1.915 0.56 ;
      RECT  2.265 0.445 3.035 0.56 ;
      RECT  2.945 0.56 3.035 0.79 ;
      RECT  2.945 0.79 4.055 0.89 ;
      RECT  2.945 0.89 3.035 1.24 ;
      RECT  0.05 1.24 3.035 1.36 ;
      RECT  4.37 1.24 5.555 1.36 ;
      RECT  4.37 1.36 4.49 1.44 ;
      RECT  3.305 1.44 4.49 1.56 ;
  END
END SEN_AN4B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN4B_8
#      Description : "4-Input AND (A inverted input)"
#      Equation    : X=!A&B1&B2&B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN4B_8
  CLASS CORE ;
  FOREIGN SEN_AN4B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.51 7.85 0.71 ;
      RECT  6.35 0.71 7.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.65 0.91 ;
      RECT  2.55 0.91 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.05 0.91 ;
      RECT  1.55 0.91 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.71 0.85 0.91 ;
      RECT  0.42 0.91 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 8.0 1.85 ;
      RECT  0.61 1.43 0.73 1.75 ;
      RECT  1.13 1.43 1.25 1.75 ;
      RECT  1.65 1.43 1.77 1.75 ;
      RECT  2.26 1.43 2.38 1.75 ;
      RECT  2.875 1.43 2.995 1.75 ;
      RECT  3.395 1.19 3.51 1.75 ;
      RECT  5.965 1.245 6.085 1.75 ;
      RECT  6.485 1.245 6.605 1.75 ;
      RECT  7.005 1.245 7.125 1.75 ;
      RECT  7.525 1.245 7.645 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      RECT  4.145 0.05 4.265 0.375 ;
      RECT  4.665 0.05 4.785 0.375 ;
      RECT  5.185 0.05 5.305 0.375 ;
      RECT  5.705 0.05 5.825 0.375 ;
      RECT  6.225 0.05 6.345 0.375 ;
      RECT  6.745 0.05 6.865 0.375 ;
      RECT  7.265 0.05 7.385 0.375 ;
      RECT  7.79 0.05 7.93 0.39 ;
      RECT  0.35 0.05 0.47 0.405 ;
      RECT  0.87 0.05 0.99 0.405 ;
      RECT  3.63 0.05 3.745 0.605 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.525 0.31 7.65 0.465 ;
      RECT  3.835 0.465 7.65 0.595 ;
      RECT  5.35 0.595 6.25 0.69 ;
      RECT  5.35 0.69 5.52 1.11 ;
      RECT  3.75 1.11 5.52 1.115 ;
      RECT  3.75 1.115 5.565 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.35 0.24 3.54 0.36 ;
      RECT  0.09 0.4 0.21 0.5 ;
      RECT  0.09 0.5 2.29 0.62 ;
      RECT  2.17 0.62 2.29 0.715 ;
      RECT  2.565 0.485 3.305 0.605 ;
      RECT  3.2 0.605 3.305 0.785 ;
      RECT  3.2 0.785 5.17 0.895 ;
      RECT  3.2 0.895 3.305 1.22 ;
      RECT  0.3 1.22 3.305 1.34 ;
      RECT  5.68 1.005 6.385 1.035 ;
      RECT  5.68 1.035 7.905 1.155 ;
      RECT  7.785 1.155 7.905 1.255 ;
      RECT  5.68 1.155 5.85 1.41 ;
      RECT  5.145 1.41 5.85 1.44 ;
      RECT  3.6 1.44 5.85 1.56 ;
  END
END SEN_AN4B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AN5_1
#      Description : "5-Input AND"
#      Equation    : X=A1&A2&A3&A4&A5
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN5_1
  CLASS CORE ;
  FOREIGN SEN_AN5_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.95 ;
      RECT  0.52 0.95 0.65 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.485 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.05 1.145 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0465 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.91 ;
      RECT  1.55 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0465 ;
  END A5
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.415 0.185 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  0.585 1.435 0.705 1.75 ;
      RECT  1.49 1.455 1.61 1.75 ;
      RECT  2.0 1.415 2.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  1.55 0.05 1.67 0.41 ;
      RECT  0.94 0.05 1.06 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.475 1.46 0.595 ;
      RECT  1.15 0.595 1.25 1.465 ;
      RECT  0.98 1.465 1.25 1.585 ;
    END
    ANTENNADIFFAREA 0.16 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.19 0.185 0.32 ;
      RECT  0.065 0.32 0.43 0.41 ;
      RECT  0.34 0.41 0.43 1.21 ;
      RECT  0.34 1.21 1.06 1.33 ;
      RECT  0.97 0.755 1.06 1.21 ;
      RECT  0.34 1.33 0.445 1.425 ;
      RECT  2.01 0.37 2.13 0.5 ;
      RECT  1.57 0.5 2.13 0.59 ;
      RECT  1.57 0.59 1.66 0.73 ;
      RECT  1.34 0.73 1.66 0.82 ;
      RECT  1.34 0.82 1.43 1.245 ;
      RECT  1.34 1.245 1.92 1.365 ;
  END
END SEN_AN5_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN5_2
#      Description : "5-Input AND"
#      Equation    : X=A1&A2&A3&A4&A5
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN5_2
  CLASS CORE ;
  FOREIGN SEN_AN5_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.102 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.102 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  1.35 0.91 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.102 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.54 0.71 3.65 0.91 ;
      RECT  3.35 0.91 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.093 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.25 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.093 ;
  END A5
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  1.105 1.415 1.225 1.75 ;
      RECT  1.625 1.415 1.745 1.75 ;
      RECT  2.655 1.43 2.775 1.75 ;
      RECT  3.14 1.465 3.31 1.75 ;
      RECT  3.685 1.455 3.805 1.75 ;
      RECT  4.215 1.21 4.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  1.355 0.05 1.475 0.36 ;
      RECT  3.945 0.05 4.065 0.36 ;
      RECT  2.395 0.05 2.515 0.385 ;
      RECT  1.875 0.05 1.995 0.6 ;
      RECT  2.915 0.05 3.035 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.085 0.475 2.8 0.595 ;
      RECT  2.35 0.595 2.45 1.04 ;
      RECT  2.15 1.04 2.45 1.13 ;
      RECT  2.15 1.13 2.255 1.29 ;
    END
    ANTENNADIFFAREA 0.288 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.215 1.265 0.335 ;
      RECT  0.065 0.335 0.185 0.435 ;
      RECT  3.125 0.24 3.805 0.36 ;
      RECT  3.685 0.36 3.805 0.45 ;
      RECT  3.685 0.45 4.325 0.54 ;
      RECT  4.205 0.32 4.325 0.45 ;
      RECT  0.795 0.475 1.785 0.595 ;
      RECT  3.155 0.475 3.595 0.595 ;
      RECT  3.155 0.595 3.245 0.755 ;
      RECT  2.635 0.755 3.245 0.865 ;
      RECT  3.155 0.865 3.245 1.245 ;
      RECT  3.155 1.245 4.115 1.365 ;
      RECT  1.755 0.755 2.235 0.865 ;
      RECT  1.755 0.865 1.845 1.215 ;
      RECT  0.275 0.475 0.645 0.595 ;
      RECT  0.555 0.595 0.645 1.215 ;
      RECT  0.275 1.215 1.845 1.32 ;
      RECT  2.395 1.22 3.065 1.34 ;
      RECT  2.395 1.34 2.515 1.405 ;
      RECT  1.875 1.405 2.515 1.495 ;
      RECT  1.875 1.495 1.995 1.615 ;
  END
END SEN_AN5_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN5_4
#      Description : "5-Input AND"
#      Equation    : X=A1&A2&A3&A4&A5
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN5_4
  CLASS CORE ;
  FOREIGN SEN_AN5_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.895 ;
      RECT  0.35 0.895 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2034 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.05 0.91 ;
      RECT  1.55 0.91 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2034 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.74 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2034 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.71 7.05 0.91 ;
      RECT  6.95 0.91 7.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1872 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.25 0.91 ;
      RECT  5.83 0.91 6.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1872 ;
  END A5
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  1.105 1.43 1.225 1.75 ;
      RECT  1.66 1.44 1.78 1.75 ;
      RECT  2.245 1.43 2.365 1.75 ;
      RECT  2.795 1.43 2.915 1.75 ;
      RECT  4.62 1.415 4.74 1.75 ;
      RECT  5.14 1.415 5.26 1.75 ;
      RECT  5.66 1.44 5.78 1.75 ;
      RECT  6.18 1.44 6.3 1.75 ;
      RECT  6.7 1.44 6.82 1.75 ;
      RECT  7.22 1.41 7.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  2.255 0.05 2.375 0.36 ;
      RECT  2.795 0.05 2.915 0.36 ;
      RECT  3.84 0.05 3.96 0.385 ;
      RECT  4.36 0.05 4.48 0.385 ;
      RECT  4.88 0.05 5.0 0.385 ;
      RECT  5.92 0.05 6.04 0.405 ;
      RECT  3.32 0.05 3.44 0.63 ;
      RECT  5.4 0.05 5.52 0.63 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.14 0.31 5.26 0.475 ;
      RECT  3.53 0.475 5.26 0.595 ;
      RECT  4.15 0.595 4.25 1.11 ;
      RECT  3.55 1.11 4.25 1.29 ;
    END
    ANTENNADIFFAREA 0.576 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.215 1.795 0.335 ;
      RECT  0.065 0.335 0.185 0.435 ;
      RECT  6.13 0.215 7.34 0.335 ;
      RECT  7.22 0.335 7.34 0.41 ;
      RECT  6.13 0.335 6.245 0.495 ;
      RECT  5.61 0.495 6.245 0.615 ;
      RECT  1.315 0.475 3.205 0.595 ;
      RECT  6.355 0.475 7.13 0.595 ;
      RECT  6.355 0.595 6.445 1.225 ;
      RECT  6.355 1.225 7.13 1.23 ;
      RECT  4.73 0.77 5.7 0.88 ;
      RECT  5.61 0.88 5.7 1.23 ;
      RECT  5.61 1.23 7.13 1.35 ;
      RECT  3.355 0.755 3.98 0.865 ;
      RECT  3.355 0.865 3.445 1.22 ;
      RECT  0.275 0.475 1.14 0.595 ;
      RECT  1.05 0.595 1.14 1.22 ;
      RECT  0.275 1.22 3.445 1.34 ;
      RECT  4.36 1.145 5.52 1.265 ;
      RECT  5.4 1.265 5.52 1.425 ;
      RECT  4.36 1.265 4.48 1.465 ;
      RECT  3.26 1.465 4.48 1.585 ;
  END
END SEN_AN5_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN5_6
#      Description : "5-Input AND"
#      Equation    : X=A1&A2&A3&A4&A5
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN5_6
  CLASS CORE ;
  FOREIGN SEN_AN5_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3054 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.91 ;
      RECT  1.75 0.91 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3054 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.05 0.91 ;
      RECT  2.95 0.91 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3054 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.08 0.71 9.85 0.89 ;
      RECT  9.75 0.89 9.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2724 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.71 7.85 0.91 ;
      RECT  7.75 0.91 8.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2724 ;
  END A5
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 10.0 1.85 ;
      RECT  0.585 1.42 0.705 1.75 ;
      RECT  1.105 1.42 1.225 1.75 ;
      RECT  1.625 1.42 1.745 1.75 ;
      RECT  2.145 1.42 2.265 1.75 ;
      RECT  2.665 1.42 2.785 1.75 ;
      RECT  3.185 1.42 3.305 1.75 ;
      RECT  3.705 1.42 3.825 1.75 ;
      RECT  5.985 1.245 6.105 1.75 ;
      RECT  6.51 1.245 6.63 1.75 ;
      RECT  7.03 1.245 7.15 1.75 ;
      RECT  7.475 1.44 7.595 1.75 ;
      RECT  7.995 1.44 8.115 1.75 ;
      RECT  8.515 1.44 8.635 1.75 ;
      RECT  9.035 1.44 9.155 1.75 ;
      RECT  9.555 1.44 9.675 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.0 0.05 ;
      RECT  2.925 0.05 3.045 0.385 ;
      RECT  3.445 0.05 3.565 0.385 ;
      RECT  4.615 0.05 4.735 0.385 ;
      RECT  5.135 0.05 5.255 0.385 ;
      RECT  5.655 0.05 5.775 0.385 ;
      RECT  6.175 0.05 6.295 0.385 ;
      RECT  6.695 0.05 6.815 0.385 ;
      RECT  7.735 0.05 7.855 0.385 ;
      RECT  8.255 0.05 8.375 0.385 ;
      RECT  4.03 0.05 4.15 0.585 ;
      RECT  7.215 0.05 7.335 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.305 0.475 7.125 0.595 ;
      RECT  5.32 0.595 5.45 1.11 ;
      RECT  4.35 1.11 5.595 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 0.24 2.575 0.36 ;
      RECT  8.515 0.24 9.725 0.36 ;
      RECT  8.515 0.36 8.635 0.475 ;
      RECT  7.425 0.475 8.635 0.595 ;
      RECT  9.815 0.4 9.935 0.5 ;
      RECT  8.775 0.5 9.935 0.62 ;
      RECT  8.775 0.62 8.895 1.23 ;
      RECT  6.2 0.755 7.625 0.865 ;
      RECT  7.535 0.865 7.625 1.23 ;
      RECT  7.535 1.23 9.935 1.35 ;
      RECT  9.815 1.35 9.935 1.45 ;
      RECT  1.57 0.475 3.88 0.595 ;
      RECT  4.165 0.755 5.215 0.865 ;
      RECT  4.165 0.865 4.255 1.205 ;
      RECT  0.065 0.4 0.185 0.5 ;
      RECT  0.065 0.5 1.455 0.62 ;
      RECT  1.365 0.62 1.455 1.205 ;
      RECT  0.275 1.205 4.255 1.325 ;
      RECT  5.72 1.035 7.445 1.155 ;
      RECT  5.72 1.155 5.84 1.465 ;
      RECT  4.11 1.465 5.84 1.585 ;
  END
END SEN_AN5_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AN6_1
#      Description : "6-Input AND"
#      Equation    : X=A1&A2&A3&A4&A5&A6
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN6_1
  CLASS CORE ;
  FOREIGN SEN_AN6_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.865 ;
      RECT  0.52 0.865 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.45 0.685 ;
      RECT  1.35 0.685 1.65 0.775 ;
      RECT  1.525 0.775 1.65 0.99 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.9 ;
      RECT  1.15 0.9 1.395 0.99 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A5
  PIN A6
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.965 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A6
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.845 1.415 0.965 1.75 ;
      RECT  1.365 1.44 1.485 1.75 ;
      RECT  2.405 1.415 2.54 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.885 0.05 2.025 0.36 ;
      RECT  0.845 0.05 0.965 0.385 ;
      RECT  2.405 0.05 2.54 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.3 2.275 0.51 ;
      RECT  2.15 0.51 2.515 0.69 ;
      RECT  2.425 0.69 2.515 1.11 ;
      RECT  2.15 1.11 2.515 1.29 ;
      RECT  2.15 1.29 2.25 1.44 ;
      RECT  1.845 1.44 2.25 1.56 ;
    END
    ANTENNADIFFAREA 0.18 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.57 0.45 2.06 0.57 ;
      RECT  1.97 0.57 2.06 0.86 ;
      RECT  1.97 0.86 2.335 0.95 ;
      RECT  2.235 0.78 2.335 0.86 ;
      RECT  1.97 0.95 2.06 1.26 ;
      RECT  1.12 1.26 2.06 1.35 ;
      RECT  1.12 1.35 1.225 1.55 ;
      RECT  1.625 1.35 1.745 1.55 ;
      RECT  1.79 0.725 1.88 1.08 ;
      RECT  0.94 1.08 1.88 1.17 ;
      RECT  0.94 1.17 1.03 1.235 ;
      RECT  0.065 0.165 0.185 0.295 ;
      RECT  0.065 0.295 0.43 0.385 ;
      RECT  0.34 0.385 0.43 1.235 ;
      RECT  0.065 1.235 1.03 1.325 ;
      RECT  0.065 1.325 0.185 1.55 ;
      RECT  0.585 1.325 0.705 1.55 ;
  END
END SEN_AN6_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AN6_2
#      Description : "6-Input AND"
#      Equation    : X=A1&A2&A3&A4&A5&A6
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN6_2
  CLASS CORE ;
  FOREIGN SEN_AN6_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.205 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.205 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.79 2.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.05 1.05 ;
      RECT  1.95 1.05 2.08 1.22 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A5
  PIN A6
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.105 ;
      RECT  1.55 1.105 1.74 1.205 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A6
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.475 0.47 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.82 1.475 1.0 1.75 ;
      RECT  1.35 1.475 1.52 1.75 ;
      RECT  1.87 1.49 2.04 1.75 ;
      RECT  2.425 1.42 2.545 1.75 ;
      RECT  3.21 1.415 3.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  2.95 0.05 3.07 0.385 ;
      RECT  3.47 0.05 3.59 0.385 ;
      RECT  4.01 0.05 4.13 0.385 ;
      RECT  1.295 0.05 1.43 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.21 0.375 3.33 0.475 ;
      RECT  3.21 0.475 4.05 0.595 ;
      RECT  3.95 0.595 4.05 1.11 ;
      RECT  3.705 1.11 4.05 1.29 ;
    END
    ANTENNADIFFAREA 0.288 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.07 0.17 2.86 0.29 ;
      RECT  0.065 0.22 0.815 0.33 ;
      RECT  0.065 0.33 0.185 0.405 ;
      RECT  1.67 0.38 2.86 0.47 ;
      RECT  1.67 0.47 1.76 0.485 ;
      RECT  2.77 0.47 2.86 0.51 ;
      RECT  1.355 0.485 1.76 0.575 ;
      RECT  2.77 0.51 3.12 0.6 ;
      RECT  1.355 0.575 1.445 1.295 ;
      RECT  3.03 0.6 3.12 0.755 ;
      RECT  3.03 0.755 3.86 0.865 ;
      RECT  0.27 0.44 0.65 0.56 ;
      RECT  0.56 0.56 0.65 1.295 ;
      RECT  0.065 1.295 1.445 1.385 ;
      RECT  0.065 1.385 0.185 1.52 ;
      RECT  0.585 1.385 0.705 1.52 ;
      RECT  1.115 1.385 1.235 1.52 ;
      RECT  2.17 0.56 2.68 0.68 ;
      RECT  2.59 0.68 2.68 0.755 ;
      RECT  2.17 0.68 2.26 1.31 ;
      RECT  2.59 0.755 2.94 0.865 ;
      RECT  2.59 0.865 2.805 0.875 ;
      RECT  2.685 0.875 2.805 1.27 ;
      RECT  1.635 1.31 2.26 1.4 ;
      RECT  2.16 1.4 2.26 1.525 ;
      RECT  1.635 1.4 1.755 1.535 ;
      RECT  2.9 1.155 3.59 1.275 ;
      RECT  3.47 1.275 3.59 1.51 ;
      RECT  3.47 1.51 4.11 1.6 ;
      RECT  3.99 1.38 4.11 1.51 ;
  END
END SEN_AN6_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AN6_4
#      Description : "6-Input AND"
#      Equation    : X=A1&A2&A3&A4&A5&A6
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN6_4
  CLASS CORE ;
  FOREIGN SEN_AN6_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 0.9 ;
      RECT  0.15 0.9 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.9 ;
      RECT  0.95 0.9 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 0.9 ;
      RECT  1.75 0.9 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 0.91 ;
      RECT  4.32 0.91 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.05 0.9 ;
      RECT  3.35 0.9 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A5
  PIN A6
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.9 3.05 1.09 ;
      RECT  2.55 1.09 2.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A6
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.44 0.435 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  0.835 1.44 0.955 1.75 ;
      RECT  1.355 1.44 1.475 1.75 ;
      RECT  1.875 1.44 1.995 1.75 ;
      RECT  2.395 1.44 2.515 1.75 ;
      RECT  2.92 1.44 3.035 1.75 ;
      RECT  3.435 1.44 3.555 1.75 ;
      RECT  3.955 1.44 4.075 1.75 ;
      RECT  4.485 1.44 4.605 1.75 ;
      RECT  5.205 1.415 5.325 1.75 ;
      RECT  5.725 1.415 5.845 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  4.91 0.05 5.08 0.23 ;
      RECT  2.37 0.05 2.54 0.34 ;
      RECT  2.89 0.05 3.06 0.34 ;
      RECT  5.44 0.05 5.61 0.345 ;
      RECT  5.96 0.05 6.13 0.345 ;
      RECT  6.48 0.05 6.65 0.345 ;
      RECT  1.875 0.05 1.995 0.38 ;
      RECT  7.015 0.05 7.145 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.205 0.32 5.325 0.435 ;
      RECT  5.205 0.435 6.885 0.535 ;
      RECT  6.75 0.31 6.885 0.435 ;
      RECT  6.75 0.535 6.85 1.11 ;
      RECT  6.24 1.11 7.05 1.29 ;
    END
    ANTENNADIFFAREA 0.576 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.195 0.14 4.81 0.23 ;
      RECT  4.72 0.23 4.81 0.32 ;
      RECT  3.195 0.23 3.285 0.43 ;
      RECT  4.72 0.32 5.07 0.41 ;
      RECT  4.98 0.41 5.07 0.625 ;
      RECT  2.37 0.43 3.285 0.52 ;
      RECT  2.37 0.52 2.46 1.23 ;
      RECT  4.98 0.625 6.225 0.715 ;
      RECT  6.135 0.715 6.225 0.755 ;
      RECT  6.135 0.755 6.6 0.865 ;
      RECT  0.055 0.175 0.175 0.475 ;
      RECT  0.055 0.475 0.845 0.595 ;
      RECT  0.755 0.595 0.845 1.23 ;
      RECT  0.055 1.23 2.46 1.35 ;
      RECT  0.055 1.35 0.175 1.635 ;
      RECT  0.265 0.22 1.525 0.34 ;
      RECT  3.385 0.345 4.63 0.465 ;
      RECT  1.045 0.495 2.28 0.615 ;
      RECT  2.605 0.61 3.86 0.73 ;
      RECT  4.745 0.5 4.865 0.805 ;
      RECT  4.745 0.805 5.8 0.915 ;
      RECT  4.745 0.915 4.855 1.23 ;
      RECT  4.14 0.595 4.39 0.715 ;
      RECT  4.14 0.715 4.23 1.23 ;
      RECT  2.74 1.23 4.855 1.35 ;
      RECT  2.74 1.35 2.83 1.44 ;
      RECT  4.745 1.35 4.855 1.635 ;
      RECT  2.605 1.44 2.83 1.56 ;
      RECT  4.945 1.005 5.065 1.205 ;
      RECT  4.945 1.205 6.105 1.325 ;
      RECT  5.985 1.325 6.105 1.47 ;
      RECT  5.985 1.47 7.145 1.59 ;
      RECT  7.025 1.41 7.145 1.47 ;
  END
END SEN_AN6_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AN6_8
#      Description : "6-Input AND"
#      Equation    : X=A1&A2&A3&A4&A5&A6
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AN6_8
  CLASS CORE ;
  FOREIGN SEN_AN6_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3234 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.55 0.91 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3234 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.25 0.91 ;
      RECT  3.35 0.91 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3234 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 7.45 0.91 ;
      RECT  7.15 0.91 7.985 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3234 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.71 6.85 0.91 ;
      RECT  5.75 0.91 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3234 ;
  END A5
  PIN A6
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.91 5.25 1.09 ;
      RECT  4.35 1.09 4.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3234 ;
  END A6
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.455 1.44 0.575 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  1.055 1.435 1.175 1.75 ;
      RECT  1.615 1.435 1.735 1.75 ;
      RECT  2.135 1.435 2.255 1.75 ;
      RECT  2.655 1.435 2.775 1.75 ;
      RECT  3.175 1.435 3.295 1.75 ;
      RECT  3.695 1.435 3.815 1.75 ;
      RECT  4.215 1.405 4.335 1.75 ;
      RECT  4.735 1.44 4.855 1.75 ;
      RECT  5.255 1.44 5.375 1.75 ;
      RECT  5.775 1.44 5.895 1.75 ;
      RECT  6.295 1.44 6.415 1.75 ;
      RECT  6.815 1.44 6.935 1.75 ;
      RECT  7.335 1.44 7.455 1.75 ;
      RECT  7.855 1.44 7.98 1.75 ;
      RECT  8.72 1.415 8.845 1.75 ;
      RECT  9.24 1.415 9.365 1.75 ;
      RECT  9.76 1.415 9.885 1.75 ;
      RECT  10.28 1.415 10.4 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  8.955 0.05 9.125 0.305 ;
      RECT  9.475 0.05 9.665 0.305 ;
      RECT  9.995 0.05 10.165 0.305 ;
      RECT  10.515 0.05 10.685 0.305 ;
      RECT  11.035 0.05 11.205 0.305 ;
      RECT  11.555 0.05 11.725 0.305 ;
      RECT  12.075 0.05 12.245 0.305 ;
      RECT  5.23 0.05 5.4 0.31 ;
      RECT  8.415 0.05 8.585 0.31 ;
      RECT  3.15 0.05 3.32 0.32 ;
      RECT  3.67 0.05 3.84 0.32 ;
      RECT  4.19 0.05 4.36 0.32 ;
      RECT  4.71 0.05 4.88 0.32 ;
      RECT  12.62 0.05 12.74 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.67 0.395 9.84 0.415 ;
      RECT  8.67 0.415 12.465 0.485 ;
      RECT  9.72 0.485 12.465 0.545 ;
      RECT  10.245 0.545 12.465 0.565 ;
      RECT  12.315 0.565 12.465 1.11 ;
      RECT  10.785 1.11 12.465 1.29 ;
    END
    ANTENNADIFFAREA 1.152 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.26 0.19 7.515 0.21 ;
      RECT  5.725 0.21 8.025 0.32 ;
      RECT  0.055 0.18 2.825 0.31 ;
      RECT  0.055 0.31 0.175 0.41 ;
      RECT  0.265 0.4 1.5 0.41 ;
      RECT  0.265 0.41 8.545 0.515 ;
      RECT  1.35 0.515 8.545 0.56 ;
      RECT  8.395 0.56 8.545 0.575 ;
      RECT  1.35 0.56 1.45 1.225 ;
      RECT  8.395 0.575 9.63 0.72 ;
      RECT  8.395 0.72 12.225 0.725 ;
      RECT  9.48 0.725 12.225 0.87 ;
      RECT  0.105 1.225 4.075 1.345 ;
      RECT  3.955 1.345 4.075 1.445 ;
      RECT  3.96 0.65 4.06 0.685 ;
      RECT  1.825 0.685 4.06 0.82 ;
      RECT  6.565 0.65 6.66 0.685 ;
      RECT  4.425 0.685 6.66 0.82 ;
      RECT  7.545 0.66 8.27 0.78 ;
      RECT  8.12 0.78 8.27 0.815 ;
      RECT  8.12 0.815 9.39 0.965 ;
      RECT  8.12 0.965 8.24 1.23 ;
      RECT  6.955 0.675 7.22 0.795 ;
      RECT  6.955 0.795 7.045 1.23 ;
      RECT  4.54 1.23 8.24 1.35 ;
      RECT  4.54 1.35 4.63 1.44 ;
      RECT  4.425 1.44 4.63 1.56 ;
      RECT  8.41 1.175 10.68 1.305 ;
      RECT  10.515 1.305 10.68 1.43 ;
      RECT  10.515 1.43 11.225 1.48 ;
      RECT  10.515 1.48 12.74 1.6 ;
      RECT  12.62 1.395 12.74 1.48 ;
  END
END SEN_AN6_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21_1
#      Description : "One 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21_1
  CLASS CORE ;
  FOREIGN SEN_AO21_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0582 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.35 1.42 0.47 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.145 1.22 1.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.96 0.05 1.08 0.35 ;
      RECT  0.065 0.05 0.185 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.45 1.1 ;
      RECT  1.35 1.1 1.525 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.545 0.44 1.25 0.56 ;
      RECT  1.15 0.56 1.25 1.03 ;
      RECT  0.94 1.03 1.25 1.125 ;
      RECT  0.94 1.125 1.04 1.44 ;
      RECT  0.855 1.44 1.04 1.56 ;
      RECT  0.065 1.21 0.795 1.33 ;
      RECT  0.065 1.33 0.185 1.43 ;
  END
END SEN_AO21_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21_2
#      Description : "One 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21_2
  CLASS CORE ;
  FOREIGN SEN_AO21_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1164 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.845 1.415 0.965 1.75 ;
      RECT  1.88 1.21 2.0 1.75 ;
      RECT  2.41 1.21 2.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  2.41 0.05 2.53 0.59 ;
      RECT  1.885 0.05 2.0 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.31 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.24 1.255 0.36 ;
      RECT  0.585 0.36 0.705 0.5 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.59 ;
      RECT  0.815 0.45 1.765 0.57 ;
      RECT  1.675 0.57 1.765 0.825 ;
      RECT  1.675 0.825 2.06 0.925 ;
      RECT  1.96 0.755 2.06 0.825 ;
      RECT  1.675 0.925 1.765 1.23 ;
      RECT  1.34 1.23 1.765 1.35 ;
      RECT  0.065 1.205 1.225 1.325 ;
      RECT  0.065 1.325 0.185 1.42 ;
      RECT  1.105 1.325 1.225 1.44 ;
      RECT  1.105 1.44 1.77 1.56 ;
  END
END SEN_AO21_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21_4
#      Description : "One 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21_4
  CLASS CORE ;
  FOREIGN SEN_AO21_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2328 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.845 1.415 0.965 1.75 ;
      RECT  1.365 1.415 1.485 1.75 ;
      RECT  1.885 1.415 2.005 1.75 ;
      RECT  3.46 1.2 3.58 1.75 ;
      RECT  4.025 1.415 4.145 1.75 ;
      RECT  4.6 1.2 4.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  4.025 0.05 4.145 0.35 ;
      RECT  2.395 0.05 2.515 0.36 ;
      RECT  2.915 0.05 3.035 0.36 ;
      RECT  0.325 0.05 0.445 0.375 ;
      RECT  0.845 0.05 0.965 0.375 ;
      RECT  3.46 0.05 3.58 0.6 ;
      RECT  4.6 0.05 4.72 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.705 0.44 4.45 0.56 ;
      RECT  4.35 0.56 4.45 1.11 ;
      RECT  3.75 1.11 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.46 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.24 2.29 0.36 ;
      RECT  1.105 0.36 1.225 0.465 ;
      RECT  0.065 0.36 0.185 0.465 ;
      RECT  0.065 0.465 1.225 0.585 ;
      RECT  1.34 0.45 3.32 0.57 ;
      RECT  3.23 0.57 3.32 0.79 ;
      RECT  3.23 0.79 4.26 0.89 ;
      RECT  3.23 0.89 3.32 1.23 ;
      RECT  2.38 1.23 3.32 1.35 ;
      RECT  0.065 1.205 2.265 1.325 ;
      RECT  0.065 1.325 0.185 1.43 ;
      RECT  2.145 1.325 2.265 1.44 ;
      RECT  2.145 1.44 3.33 1.56 ;
  END
END SEN_AO21_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21_DG_1
#      Description : "One 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21_DG_1
  CLASS CORE ;
  FOREIGN SEN_AO21_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.08 1.39 1.2 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  0.845 0.05 0.965 0.41 ;
      RECT  1.08 0.05 1.2 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.45 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.19 0.705 0.505 ;
      RECT  0.585 0.505 1.25 0.595 ;
      RECT  1.15 0.595 1.25 1.19 ;
      RECT  0.845 1.19 1.25 1.28 ;
      RECT  0.845 1.28 0.965 1.58 ;
      RECT  0.065 1.235 0.705 1.325 ;
      RECT  0.585 1.325 0.705 1.555 ;
      RECT  0.065 1.325 0.185 1.58 ;
  END
END SEN_AO21_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21_DG_2
#      Description : "One 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21_DG_2
  CLASS CORE ;
  FOREIGN SEN_AO21_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.41 0.445 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.095 1.39 1.215 1.75 ;
      RECT  1.605 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  1.605 0.05 1.74 0.39 ;
      RECT  0.845 0.05 0.965 0.41 ;
      RECT  1.095 0.05 1.215 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.475 0.51 ;
      RECT  1.35 0.51 1.65 0.6 ;
      RECT  1.55 0.6 1.65 1.11 ;
      RECT  1.35 1.11 1.65 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.215 0.705 0.5 ;
      RECT  0.585 0.5 1.24 0.59 ;
      RECT  1.15 0.59 1.24 0.775 ;
      RECT  1.15 0.775 1.45 0.895 ;
      RECT  1.15 0.895 1.24 1.205 ;
      RECT  0.845 1.205 1.24 1.295 ;
      RECT  0.845 1.295 0.965 1.525 ;
      RECT  0.065 1.23 0.705 1.32 ;
      RECT  0.065 1.32 0.185 1.525 ;
      RECT  0.585 1.32 0.705 1.525 ;
  END
END SEN_AO21_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21_DG_4
#      Description : "One 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21_DG_4
  CLASS CORE ;
  FOREIGN SEN_AO21_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.125 1.39 1.245 1.75 ;
      RECT  1.675 1.41 1.795 1.75 ;
      RECT  2.2 1.21 2.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  1.675 0.05 1.795 0.395 ;
      RECT  0.865 0.05 0.985 0.41 ;
      RECT  1.13 0.05 1.25 0.41 ;
      RECT  2.2 0.05 2.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.41 0.355 1.53 0.485 ;
      RECT  1.41 0.485 2.05 0.575 ;
      RECT  1.95 0.575 2.05 1.11 ;
      RECT  1.35 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.365 0.705 0.52 ;
      RECT  0.585 0.52 1.245 0.61 ;
      RECT  1.155 0.61 1.245 0.785 ;
      RECT  1.155 0.785 1.855 0.895 ;
      RECT  1.155 0.895 1.245 1.19 ;
      RECT  0.845 1.19 1.245 1.28 ;
      RECT  0.845 1.28 0.965 1.41 ;
      RECT  0.065 1.205 0.755 1.325 ;
      RECT  0.065 1.325 0.185 1.43 ;
  END
END SEN_AO21_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21_8
#      Description : "One 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21_8
  CLASS CORE ;
  FOREIGN SEN_AO21_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 3.45 0.9 ;
      RECT  3.35 0.9 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4536 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.65 0.9 ;
      RECT  1.55 0.9 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4536 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 5.25 0.9 ;
      RECT  5.15 0.9 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4248 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.43 0.445 1.75 ;
      RECT  0.0 1.75 8.0 1.85 ;
      RECT  0.845 1.43 0.965 1.75 ;
      RECT  1.365 1.43 1.485 1.75 ;
      RECT  1.885 1.455 2.005 1.75 ;
      RECT  2.405 1.455 2.525 1.75 ;
      RECT  2.925 1.455 3.045 1.75 ;
      RECT  3.445 1.455 3.565 1.75 ;
      RECT  5.735 1.395 5.855 1.75 ;
      RECT  6.255 1.405 6.375 1.75 ;
      RECT  6.775 1.405 6.895 1.75 ;
      RECT  7.295 1.405 7.415 1.75 ;
      RECT  7.815 1.21 7.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      RECT  4.0 0.05 4.12 0.36 ;
      RECT  4.6 0.05 4.72 0.36 ;
      RECT  5.215 0.05 5.335 0.36 ;
      RECT  0.585 0.05 0.705 0.38 ;
      RECT  1.105 0.05 1.225 0.38 ;
      RECT  1.625 0.05 1.745 0.38 ;
      RECT  6.255 0.05 6.375 0.395 ;
      RECT  6.775 0.05 6.895 0.395 ;
      RECT  7.295 0.05 7.415 0.395 ;
      RECT  5.735 0.05 5.855 0.4 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  7.815 0.05 7.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.94 0.49 7.675 0.62 ;
      RECT  7.505 0.62 7.675 1.11 ;
      RECT  5.95 1.11 7.675 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.87 0.23 3.59 0.36 ;
      RECT  1.87 0.36 2.02 0.47 ;
      RECT  0.275 0.47 2.02 0.6 ;
      RECT  2.12 0.45 5.66 0.6 ;
      RECT  5.51 0.6 5.66 0.775 ;
      RECT  5.51 0.775 7.39 0.9 ;
      RECT  5.51 0.9 6.705 0.925 ;
      RECT  5.51 0.925 5.66 1.215 ;
      RECT  3.93 1.215 5.66 1.345 ;
      RECT  0.065 1.215 3.84 1.335 ;
      RECT  1.585 1.335 3.84 1.365 ;
      RECT  0.065 1.335 0.185 1.44 ;
      RECT  3.69 1.365 3.84 1.435 ;
      RECT  3.69 1.435 5.435 1.565 ;
  END
END SEN_AO21_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21B_1
#      Description : "One 2-input NAND into 2-input NAND"
#      Equation    : X=(A1&A2)|!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21B_1
  CLASS CORE ;
  FOREIGN SEN_AO21B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.71 ;
      RECT  0.35 0.71 0.495 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.42 0.175 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.63 1.4 0.75 1.75 ;
      RECT  1.225 1.415 1.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.225 0.05 1.345 0.375 ;
      RECT  0.055 0.05 0.175 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.775 0.51 1.05 0.69 ;
      RECT  0.95 0.69 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.199 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.19 0.685 0.785 ;
      RECT  0.585 0.785 0.86 0.895 ;
      RECT  0.585 0.895 0.685 1.21 ;
      RECT  0.315 1.21 0.685 1.3 ;
      RECT  0.315 1.3 0.435 1.49 ;
  END
END SEN_AO21B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21B_2
#      Description : "One 2-input NAND into 2-input NAND"
#      Equation    : X=(A1&A2)|!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21B_2
  CLASS CORE ;
  FOREIGN SEN_AO21B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 0.91 ;
      RECT  0.75 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0852 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0852 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.415 0.185 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.56 1.47 0.73 1.75 ;
      RECT  1.21 1.47 1.38 1.75 ;
      RECT  1.875 1.41 1.995 1.75 ;
      RECT  2.395 1.21 2.515 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.325 0.05 0.445 0.35 ;
      RECT  2.135 0.05 2.255 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.72 0.69 ;
      RECT  1.55 0.69 1.65 1.11 ;
      RECT  1.55 1.11 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.23 1.25 0.35 ;
      RECT  0.585 0.35 0.705 0.44 ;
      RECT  0.065 0.31 0.185 0.44 ;
      RECT  0.065 0.44 0.705 0.56 ;
      RECT  1.355 0.24 1.995 0.36 ;
      RECT  1.875 0.36 1.995 0.44 ;
      RECT  1.355 0.36 1.475 0.455 ;
      RECT  1.875 0.44 2.555 0.56 ;
      RECT  0.805 0.44 1.24 0.56 ;
      RECT  1.15 0.56 1.24 0.78 ;
      RECT  1.15 0.78 1.46 0.89 ;
      RECT  1.15 0.89 1.24 1.26 ;
      RECT  0.29 1.26 1.24 1.38 ;
  END
END SEN_AO21B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21B_4
#      Description : "One 2-input NAND into 2-input NAND"
#      Equation    : X=(A1&A2)|!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21B_4
  CLASS CORE ;
  FOREIGN SEN_AO21B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  0.95 0.91 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1707 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.215 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.585 1.42 0.705 1.75 ;
      RECT  1.105 1.42 1.225 1.75 ;
      RECT  1.72 1.42 1.84 1.75 ;
      RECT  2.33 1.41 2.45 1.75 ;
      RECT  2.85 1.41 2.97 1.75 ;
      RECT  3.385 1.41 3.505 1.75 ;
      RECT  3.94 1.21 4.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  3.11 0.05 3.23 0.35 ;
      RECT  3.645 0.05 3.765 0.35 ;
      RECT  0.065 0.05 0.185 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.71 0.69 ;
      RECT  2.55 0.69 2.65 1.11 ;
      RECT  1.95 1.11 3.77 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.76 0.215 2.97 0.335 ;
      RECT  2.85 0.335 2.97 0.44 ;
      RECT  2.85 0.44 4.08 0.56 ;
      RECT  0.845 0.24 1.54 0.36 ;
      RECT  0.845 0.36 0.965 0.44 ;
      RECT  0.3 0.44 0.965 0.56 ;
      RECT  1.055 0.5 1.81 0.62 ;
      RECT  1.72 0.62 1.81 0.785 ;
      RECT  1.72 0.785 2.46 0.895 ;
      RECT  1.72 0.895 1.81 1.21 ;
      RECT  0.285 1.21 1.81 1.33 ;
  END
END SEN_AO21B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21B_16
#      Description : "One 2-input NAND into 2-input NAND"
#      Equation    : X=(A1&A2)|!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21B_16
  CLASS CORE ;
  FOREIGN SEN_AO21B_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 4.85 0.91 ;
      RECT  3.55 0.91 5.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6939 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 0.91 ;
      RECT  0.55 0.91 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6939 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.15 0.71 14.45 0.815 ;
      RECT  11.15 0.815 14.45 0.91 ;
      RECT  14.35 0.91 14.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9873 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 14.6 1.85 ;
      RECT  0.585 1.455 0.705 1.75 ;
      RECT  1.105 1.455 1.225 1.75 ;
      RECT  1.625 1.455 1.745 1.75 ;
      RECT  2.145 1.455 2.265 1.75 ;
      RECT  2.665 1.455 2.785 1.75 ;
      RECT  3.185 1.455 3.305 1.75 ;
      RECT  3.705 1.455 3.825 1.75 ;
      RECT  4.225 1.455 4.345 1.75 ;
      RECT  4.745 1.455 4.865 1.75 ;
      RECT  5.265 1.455 5.385 1.75 ;
      RECT  5.76 1.455 5.935 1.75 ;
      RECT  6.035 1.215 6.155 1.75 ;
      RECT  6.555 1.415 6.675 1.75 ;
      RECT  7.075 1.415 7.195 1.75 ;
      RECT  7.595 1.415 7.715 1.75 ;
      RECT  8.115 1.415 8.235 1.75 ;
      RECT  8.635 1.415 8.755 1.75 ;
      RECT  9.155 1.415 9.275 1.75 ;
      RECT  9.65 1.47 9.82 1.75 ;
      RECT  10.205 1.47 10.375 1.75 ;
      RECT  10.75 1.455 10.92 1.75 ;
      RECT  11.295 1.43 11.415 1.75 ;
      RECT  11.815 1.415 11.935 1.75 ;
      RECT  12.335 1.415 12.455 1.75 ;
      RECT  12.855 1.415 12.975 1.75 ;
      RECT  13.375 1.415 13.495 1.75 ;
      RECT  13.895 1.415 14.015 1.75 ;
      RECT  14.415 1.21 14.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 14.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 14.6 0.05 ;
      RECT  11.01 0.05 11.18 0.32 ;
      RECT  11.53 0.05 11.7 0.32 ;
      RECT  12.05 0.05 12.22 0.34 ;
      RECT  0.585 0.05 0.705 0.345 ;
      RECT  1.105 0.05 1.225 0.345 ;
      RECT  1.625 0.05 1.745 0.345 ;
      RECT  2.145 0.05 2.265 0.345 ;
      RECT  2.665 0.05 2.785 0.345 ;
      RECT  10.53 0.05 10.635 0.345 ;
      RECT  12.595 0.05 12.715 0.36 ;
      RECT  13.115 0.05 13.235 0.385 ;
      RECT  13.635 0.05 13.755 0.385 ;
      RECT  14.155 0.05 14.275 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 14.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.245 0.51 9.055 0.54 ;
      RECT  6.245 0.54 9.61 0.57 ;
      RECT  6.245 0.57 10.05 0.63 ;
      RECT  7.325 0.63 10.05 0.69 ;
      RECT  8.855 0.69 10.05 0.745 ;
      RECT  8.855 0.745 9.65 0.77 ;
      RECT  9.35 0.77 9.65 1.07 ;
      RECT  9.35 1.07 10.67 1.11 ;
      RECT  6.28 1.11 14.26 1.29 ;
      RECT  8.35 1.29 12.21 1.3 ;
      RECT  8.35 1.3 11.69 1.325 ;
      RECT  9.35 1.325 11.185 1.365 ;
    END
    ANTENNADIFFAREA 2.537 ;
  END X
  OBS
      LAYER M1 ;
      RECT  8.1 0.16 10.44 0.195 ;
      RECT  6.035 0.195 10.44 0.345 ;
      RECT  8.615 0.345 10.44 0.375 ;
      RECT  6.035 0.345 6.155 0.415 ;
      RECT  9.13 0.375 10.44 0.425 ;
      RECT  9.655 0.425 10.44 0.435 ;
      RECT  9.655 0.435 12.48 0.46 ;
      RECT  10.14 0.46 12.48 0.47 ;
      RECT  10.14 0.47 12.99 0.5 ;
      RECT  10.14 0.5 14.535 0.62 ;
      RECT  14.415 0.4 14.535 0.5 ;
      RECT  10.14 0.62 11.95 0.65 ;
      RECT  10.14 0.65 11.415 0.695 ;
      RECT  10.14 0.695 10.905 0.735 ;
      RECT  2.875 0.16 4.625 0.2 ;
      RECT  2.875 0.2 5.7 0.315 ;
      RECT  2.875 0.315 4.1 0.355 ;
      RECT  2.875 0.355 3.57 0.385 ;
      RECT  2.875 0.385 3.1 0.435 ;
      RECT  0.275 0.435 3.1 0.59 ;
      RECT  1.875 0.59 3.1 0.66 ;
      RECT  4.22 0.425 5.92 0.445 ;
      RECT  3.64 0.445 5.92 0.5 ;
      RECT  3.19 0.5 5.92 0.62 ;
      RECT  5.24 0.62 5.92 0.645 ;
      RECT  3.19 0.62 3.77 0.665 ;
      RECT  5.695 0.645 5.92 0.74 ;
      RECT  3.19 0.665 3.34 1.175 ;
      RECT  5.695 0.74 7.23 0.805 ;
      RECT  5.695 0.805 8.495 0.86 ;
      RECT  5.695 0.86 9.205 0.965 ;
      RECT  5.695 0.965 5.92 1.235 ;
      RECT  2.89 1.175 3.34 1.225 ;
      RECT  2.385 1.225 3.34 1.235 ;
      RECT  2.385 1.235 5.92 1.245 ;
      RECT  0.325 1.245 5.92 1.365 ;
      RECT  0.325 1.365 0.445 1.465 ;
  END
END SEN_AO21B_16
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21B_6
#      Description : "One 2-input NAND into 2-input NAND"
#      Equation    : X=(A1&A2)|!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21B_6
  CLASS CORE ;
  FOREIGN SEN_AO21B_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.55 0.91 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2625 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.25 0.91 ;
      RECT  0.35 0.91 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2625 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.85 0.915 ;
      RECT  5.75 0.915 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3708 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  1.625 1.44 1.745 1.75 ;
      RECT  2.145 1.44 2.265 1.75 ;
      RECT  2.67 1.415 2.79 1.75 ;
      RECT  3.19 1.39 3.31 1.75 ;
      RECT  3.71 1.39 3.83 1.75 ;
      RECT  4.23 1.39 4.35 1.75 ;
      RECT  4.75 1.39 4.87 1.75 ;
      RECT  5.27 1.39 5.39 1.75 ;
      RECT  5.795 1.21 5.915 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  0.585 0.05 0.705 0.36 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  4.49 0.05 4.61 0.38 ;
      RECT  5.01 0.05 5.13 0.38 ;
      RECT  5.535 0.05 5.655 0.38 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 4.08 0.69 ;
      RECT  3.95 0.69 4.08 1.11 ;
      RECT  2.75 1.11 5.65 1.29 ;
    END
    ANTENNADIFFAREA 0.95 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.365 0.24 2.55 0.36 ;
      RECT  1.365 0.36 1.485 0.475 ;
      RECT  0.275 0.475 1.485 0.595 ;
      RECT  2.64 0.24 4.35 0.36 ;
      RECT  4.23 0.36 4.35 0.47 ;
      RECT  4.23 0.47 5.915 0.59 ;
      RECT  5.795 0.365 5.915 0.47 ;
      RECT  1.575 0.47 2.605 0.59 ;
      RECT  2.49 0.59 2.605 0.805 ;
      RECT  2.49 0.805 3.84 0.915 ;
      RECT  2.49 0.915 2.605 1.225 ;
      RECT  0.275 1.225 2.605 1.345 ;
  END
END SEN_AO21B_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AO21B_8
#      Description : "One 2-input NAND into 2-input NAND"
#      Equation    : X=(A1&A2)|!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO21B_8
  CLASS CORE ;
  FOREIGN SEN_AO21B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.895 ;
      RECT  1.75 0.895 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.348 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.9 ;
      RECT  0.35 0.9 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.348 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.71 7.65 0.905 ;
      RECT  7.55 0.905 7.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.585 1.415 0.7 1.75 ;
      RECT  1.105 1.415 1.22 1.75 ;
      RECT  1.625 1.415 1.74 1.75 ;
      RECT  2.145 1.415 2.26 1.75 ;
      RECT  2.665 1.415 2.78 1.75 ;
      RECT  3.185 1.19 3.305 1.75 ;
      RECT  3.435 1.19 3.555 1.75 ;
      RECT  3.955 1.39 4.075 1.75 ;
      RECT  4.475 1.39 4.595 1.75 ;
      RECT  4.995 1.39 5.115 1.75 ;
      RECT  5.515 1.39 5.635 1.75 ;
      RECT  6.035 1.39 6.155 1.75 ;
      RECT  6.555 1.39 6.675 1.75 ;
      RECT  7.075 1.39 7.195 1.75 ;
      RECT  7.61 1.21 7.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  5.775 0.05 5.895 0.36 ;
      RECT  6.295 0.05 6.415 0.36 ;
      RECT  0.325 0.05 0.445 0.385 ;
      RECT  0.845 0.05 0.965 0.385 ;
      RECT  1.365 0.05 1.485 0.385 ;
      RECT  6.815 0.05 6.935 0.385 ;
      RECT  7.335 0.05 7.455 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.635 0.51 5.4 0.69 ;
      RECT  5.08 0.69 5.4 0.7 ;
      RECT  5.08 0.7 5.25 1.11 ;
      RECT  3.675 1.11 7.45 1.29 ;
    END
    ANTENNADIFFAREA 1.264 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.62 0.21 3.345 0.34 ;
      RECT  1.62 0.34 1.75 0.475 ;
      RECT  0.065 0.375 0.185 0.475 ;
      RECT  0.065 0.475 1.75 0.595 ;
      RECT  3.435 0.225 5.65 0.375 ;
      RECT  3.435 0.375 3.555 0.445 ;
      RECT  5.5 0.375 5.65 0.45 ;
      RECT  5.5 0.45 6.7 0.5 ;
      RECT  5.5 0.5 7.715 0.62 ;
      RECT  7.595 0.4 7.715 0.5 ;
      RECT  1.84 0.465 3.095 0.595 ;
      RECT  2.965 0.595 3.095 0.8 ;
      RECT  2.965 0.8 4.91 0.93 ;
      RECT  2.965 0.93 3.095 1.195 ;
      RECT  0.275 1.195 3.095 1.325 ;
  END
END SEN_AO21B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AO221_0P5
#      Description : "Two 2-input ANDs into 3 input OR"
#      Equation    : X=(A1&A2)|(B1&B2)|C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO221_0P5
  CLASS CORE ;
  FOREIGN SEN_AO221_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0261 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.68 0.65 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0261 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.26 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.15 0.89 1.26 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0261 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.54 0.665 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0261 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.68 0.25 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0261 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.16 1.43 1.28 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.67 1.41 1.81 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.35 0.05 0.47 0.385 ;
      RECT  1.68 0.05 1.8 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.21 2.05 1.53 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.56 0.24 1.45 0.36 ;
      RECT  0.56 0.36 0.66 0.475 ;
      RECT  1.35 0.36 1.45 0.475 ;
      RECT  0.08 0.19 0.2 0.475 ;
      RECT  0.08 0.475 0.66 0.575 ;
      RECT  1.35 0.475 1.86 0.575 ;
      RECT  0.355 0.575 0.445 1.235 ;
      RECT  1.76 0.575 1.86 0.79 ;
      RECT  0.08 1.235 0.445 1.325 ;
      RECT  0.08 1.325 0.2 1.57 ;
      RECT  0.595 1.25 1.54 1.34 ;
      RECT  0.595 1.34 0.765 1.46 ;
      RECT  1.42 1.34 1.54 1.57 ;
      RECT  0.34 1.43 0.46 1.57 ;
      RECT  0.34 1.57 1.0 1.66 ;
      RECT  0.88 1.43 1.0 1.57 ;
  END
END SEN_AO221_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AO221_1
#      Description : "Two 2-input ANDs into 3 input OR"
#      Equation    : X=(A1&A2)|(B1&B2)|C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO221_1
  CLASS CORE ;
  FOREIGN SEN_AO221_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.86 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.7 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.5 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.91 ;
      RECT  1.35 0.91 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.24 0.71 0.45 0.9 ;
      RECT  0.35 0.9 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0582 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.11 1.42 1.23 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.655 1.215 1.775 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.325 0.05 0.445 0.385 ;
      RECT  1.605 0.05 1.725 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.57 0.27 1.45 0.39 ;
      RECT  0.57 0.39 0.66 0.5 ;
      RECT  1.35 0.39 1.45 0.5 ;
      RECT  0.06 0.35 0.19 0.5 ;
      RECT  0.06 0.5 0.66 0.59 ;
      RECT  1.35 0.5 1.86 0.59 ;
      RECT  0.06 0.59 0.15 1.2 ;
      RECT  1.77 0.59 1.86 0.925 ;
      RECT  0.06 1.2 0.185 1.4 ;
      RECT  0.56 1.21 1.54 1.33 ;
      RECT  0.3 1.45 1.005 1.57 ;
  END
END SEN_AO221_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO221_2
#      Description : "Two 2-input ANDs into 3 input OR"
#      Equation    : X=(A1&A2)|(B1&B2)|C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO221_2
  CLASS CORE ;
  FOREIGN SEN_AO221_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 0.71 ;
      RECT  1.75 0.71 2.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 0.71 ;
      RECT  1.35 0.71 1.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.02 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1164 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.42 0.445 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.845 1.42 0.965 1.75 ;
      RECT  3.12 1.0 3.225 1.75 ;
      RECT  3.625 1.41 3.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  1.535 0.05 1.705 0.19 ;
      RECT  3.625 0.05 3.745 0.36 ;
      RECT  0.325 0.05 0.445 0.365 ;
      RECT  3.12 0.05 3.225 0.575 ;
      RECT  2.575 0.05 2.695 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.34 0.45 3.65 0.57 ;
      RECT  3.55 0.57 3.65 1.11 ;
      RECT  3.35 1.11 3.65 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.19 1.21 0.28 ;
      RECT  1.105 0.28 1.21 0.365 ;
      RECT  0.585 0.28 0.705 0.455 ;
      RECT  0.065 0.33 0.185 0.455 ;
      RECT  0.065 0.455 0.705 0.545 ;
      RECT  2.35 0.2 2.47 0.285 ;
      RECT  1.3 0.285 2.47 0.41 ;
      RECT  1.3 0.41 1.41 0.62 ;
      RECT  2.8 0.44 3.03 0.56 ;
      RECT  2.94 0.56 3.03 0.785 ;
      RECT  2.94 0.785 3.46 0.895 ;
      RECT  2.94 0.895 3.03 1.21 ;
      RECT  2.05 0.5 2.445 0.62 ;
      RECT  2.355 0.62 2.445 1.03 ;
      RECT  0.82 0.465 1.21 0.585 ;
      RECT  1.12 0.585 1.21 1.03 ;
      RECT  1.12 1.03 2.445 1.12 ;
      RECT  2.355 1.12 2.445 1.21 ;
      RECT  2.355 1.21 3.03 1.33 ;
      RECT  0.065 1.21 2.235 1.33 ;
      RECT  0.065 1.33 0.185 1.43 ;
      RECT  1.24 1.465 3.015 1.585 ;
  END
END SEN_AO221_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO221_4
#      Description : "Two 2-input ANDs into 3 input OR"
#      Equation    : X=(A1&A2)|(B1&B2)|C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO221_4
  CLASS CORE ;
  FOREIGN SEN_AO221_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.45 0.71 ;
      RECT  3.35 0.71 4.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.51 3.05 0.71 ;
      RECT  2.55 0.71 3.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.45 0.89 ;
      RECT  4.95 0.89 5.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2328 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.42 0.445 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.845 1.42 0.965 1.75 ;
      RECT  1.365 1.42 1.485 1.75 ;
      RECT  1.885 1.42 2.005 1.75 ;
      RECT  5.755 1.21 5.875 1.75 ;
      RECT  6.275 1.405 6.395 1.75 ;
      RECT  6.795 1.21 6.915 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  2.575 0.05 2.745 0.195 ;
      RECT  3.115 0.05 3.285 0.195 ;
      RECT  5.23 0.05 5.35 0.35 ;
      RECT  6.275 0.05 6.395 0.36 ;
      RECT  0.325 0.05 0.445 0.365 ;
      RECT  0.845 0.05 0.965 0.365 ;
      RECT  4.71 0.05 4.83 0.585 ;
      RECT  5.755 0.05 5.86 0.59 ;
      RECT  6.795 0.05 6.915 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.51 6.65 0.69 ;
      RECT  6.55 0.69 6.65 1.11 ;
      RECT  6.0 1.11 6.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.145 0.16 2.25 0.24 ;
      RECT  1.105 0.24 2.25 0.36 ;
      RECT  1.105 0.36 1.225 0.455 ;
      RECT  0.065 0.35 0.185 0.455 ;
      RECT  0.065 0.455 1.225 0.575 ;
      RECT  2.34 0.285 4.6 0.41 ;
      RECT  2.34 0.41 2.45 0.65 ;
      RECT  4.935 0.44 5.645 0.56 ;
      RECT  5.555 0.56 5.645 0.785 ;
      RECT  5.555 0.785 6.46 0.895 ;
      RECT  5.555 0.895 5.645 1.21 ;
      RECT  3.63 0.5 4.545 0.62 ;
      RECT  4.455 0.62 4.545 1.03 ;
      RECT  1.34 0.5 2.23 0.62 ;
      RECT  2.14 0.62 2.23 1.03 ;
      RECT  2.14 1.03 4.545 1.12 ;
      RECT  4.455 1.12 4.545 1.21 ;
      RECT  4.455 1.21 5.645 1.33 ;
      RECT  0.065 1.21 4.335 1.33 ;
      RECT  0.065 1.33 0.185 1.43 ;
      RECT  2.28 1.465 5.635 1.585 ;
  END
END SEN_AO221_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2222_1
#      Description : "4 NAND2s into a NAND4"
#      Equation    : X=(A1&A2)|(B1&B2)|(C1&C2)|(D1&D2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2222_1
  CLASS CORE ;
  FOREIGN SEN_AO2222_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.525 0.51 0.65 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.945 0.31 1.05 0.71 ;
      RECT  0.945 0.71 1.075 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.95 ;
      RECT  0.75 0.95 0.865 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.94 0.71 3.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.91 ;
      RECT  2.75 0.91 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END C2
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0435 ;
  END D2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.595 1.395 0.715 1.75 ;
      RECT  1.23 1.605 1.4 1.75 ;
      RECT  1.9 1.6 2.07 1.75 ;
      RECT  2.445 1.6 2.615 1.75 ;
      RECT  3.045 1.395 3.165 1.75 ;
      RECT  3.605 1.41 3.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  2.43 0.05 2.63 0.225 ;
      RECT  3.605 0.05 3.74 0.39 ;
      RECT  0.595 0.05 0.715 0.405 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.345 0.235 2.05 0.355 ;
      RECT  1.95 0.355 2.05 1.31 ;
      RECT  1.62 1.31 2.305 1.49 ;
    END
    ANTENNADIFFAREA 0.273 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.185 0.185 0.315 ;
      RECT  0.065 0.315 0.43 0.405 ;
      RECT  0.34 0.405 0.43 1.21 ;
      RECT  0.34 1.21 1.345 1.3 ;
      RECT  1.23 0.785 1.345 1.21 ;
      RECT  0.34 1.3 0.445 1.52 ;
      RECT  2.97 0.18 3.09 0.315 ;
      RECT  2.14 0.315 3.09 0.405 ;
      RECT  2.14 0.405 2.25 1.13 ;
      RECT  2.14 1.13 2.525 1.22 ;
      RECT  2.415 1.22 2.525 1.39 ;
      RECT  2.415 1.39 2.9 1.51 ;
      RECT  1.14 0.34 1.255 0.47 ;
      RECT  1.14 0.47 1.525 0.56 ;
      RECT  1.435 0.56 1.525 0.81 ;
      RECT  1.435 0.81 1.825 0.98 ;
      RECT  1.435 0.98 1.525 1.405 ;
      RECT  0.815 1.405 1.525 1.515 ;
      RECT  2.36 0.5 3.46 0.62 ;
      RECT  2.36 0.62 2.46 1.03 ;
      RECT  3.345 0.62 3.46 1.45 ;
  END
END SEN_AO2222_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2222_2
#      Description : "4 NAND2s into a NAND4"
#      Equation    : X=(A1&A2)|(B1&B2)|(C1&C2)|(D1&D2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2222_2
  CLASS CORE ;
  FOREIGN SEN_AO2222_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.89 1.45 1.1 ;
      RECT  1.15 1.1 1.45 1.205 ;
      RECT  1.15 1.205 1.25 1.35 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.05 1.19 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.21 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.71 6.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.71 5.85 1.21 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END C2
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.9 5.25 1.1 ;
      RECT  5.15 1.1 5.45 1.215 ;
      RECT  5.35 1.215 5.45 1.35 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 1.2 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END D2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.56 1.495 0.73 1.75 ;
      RECT  1.08 1.47 1.25 1.75 ;
      RECT  1.6 1.495 1.77 1.75 ;
      RECT  2.12 1.495 2.29 1.75 ;
      RECT  2.665 1.38 2.785 1.75 ;
      RECT  3.24 1.38 3.36 1.75 ;
      RECT  3.815 1.38 3.935 1.75 ;
      RECT  4.31 1.495 4.48 1.75 ;
      RECT  4.83 1.495 5.0 1.75 ;
      RECT  5.35 1.48 5.52 1.75 ;
      RECT  5.87 1.495 6.04 1.75 ;
      RECT  6.405 1.41 6.54 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.535 0.05 1.705 0.185 ;
      RECT  4.09 0.05 4.26 0.2 ;
      RECT  4.88 0.05 5.05 0.2 ;
      RECT  0.845 0.05 0.965 0.39 ;
      RECT  5.62 0.05 5.74 0.42 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.325 0.595 2.525 0.7 ;
      RECT  2.42 0.7 2.525 1.11 ;
      RECT  2.42 1.11 4.25 1.29 ;
      RECT  3.15 0.71 3.25 1.11 ;
      RECT  2.95 1.29 3.05 1.49 ;
    END
    ANTENNADIFFAREA 0.502 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.83 0.195 1.95 0.275 ;
      RECT  1.24 0.275 1.95 0.395 ;
      RECT  2.04 0.215 3.31 0.32 ;
      RECT  4.385 0.23 4.505 0.32 ;
      RECT  3.845 0.32 4.505 0.43 ;
      RECT  3.845 0.43 3.965 0.68 ;
      RECT  3.34 0.59 3.445 0.68 ;
      RECT  3.34 0.68 3.965 0.78 ;
      RECT  0.065 0.23 0.755 0.35 ;
      RECT  0.065 0.35 0.185 0.45 ;
      RECT  5.83 0.23 6.535 0.35 ;
      RECT  6.415 0.35 6.535 0.45 ;
      RECT  4.595 0.29 5.32 0.41 ;
      RECT  2.045 0.415 2.735 0.485 ;
      RECT  0.27 0.485 2.735 0.505 ;
      RECT  0.27 0.505 2.135 0.585 ;
      RECT  2.635 0.505 2.735 0.825 ;
      RECT  0.27 0.585 0.45 0.605 ;
      RECT  0.35 0.605 0.45 1.3 ;
      RECT  2.635 0.825 2.965 0.945 ;
      RECT  0.35 1.3 1.015 1.38 ;
      RECT  0.325 1.38 1.015 1.405 ;
      RECT  0.325 1.405 0.445 1.575 ;
      RECT  2.83 0.41 3.755 0.5 ;
      RECT  6.05 0.475 6.325 0.52 ;
      RECT  4.065 0.52 6.325 0.61 ;
      RECT  4.065 0.61 4.155 0.88 ;
      RECT  5.95 0.61 6.05 1.3 ;
      RECT  3.515 0.88 4.155 0.99 ;
      RECT  5.585 1.3 6.26 1.405 ;
      RECT  6.155 1.405 6.26 1.525 ;
      RECT  1.08 0.675 1.645 0.765 ;
      RECT  1.08 0.765 1.17 0.795 ;
      RECT  1.555 0.765 1.645 1.3 ;
      RECT  1.03 0.795 1.17 0.975 ;
      RECT  1.375 1.3 2.33 1.405 ;
      RECT  2.24 0.815 2.33 1.3 ;
      RECT  1.375 1.405 1.475 1.53 ;
      RECT  4.955 0.7 5.52 0.79 ;
      RECT  5.43 0.79 5.52 0.805 ;
      RECT  4.955 0.79 5.045 1.3 ;
      RECT  5.43 0.805 5.555 0.98 ;
      RECT  4.245 0.85 4.445 1.02 ;
      RECT  4.355 1.02 4.445 1.3 ;
      RECT  4.355 1.3 5.045 1.305 ;
      RECT  4.355 1.305 5.225 1.405 ;
      RECT  5.125 1.405 5.225 1.54 ;
  END
END SEN_AO2222_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2222_4
#      Description : "4 NAND2s into a NAND4"
#      Equation    : X=(A1&A2)|(B1&B2)|(C1&C2)|(D1&D2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2222_4
  CLASS CORE ;
  FOREIGN SEN_AO2222_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1575 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.91 ;
      RECT  2.15 0.91 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.65 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1575 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.15 0.3 9.25 0.71 ;
      RECT  8.95 0.71 9.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 0.71 8.85 0.92 ;
      RECT  8.55 0.92 8.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1575 ;
  END C2
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.55 0.71 7.65 0.91 ;
      RECT  7.35 0.91 7.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.51 8.25 0.71 ;
      RECT  7.75 0.71 8.25 0.89 ;
      RECT  8.15 0.89 8.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1575 ;
  END D2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.43 0.455 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.855 1.43 0.975 1.75 ;
      RECT  1.375 1.41 1.495 1.75 ;
      RECT  1.955 1.45 2.075 1.75 ;
      RECT  2.52 1.45 2.64 1.75 ;
      RECT  3.045 1.415 3.165 1.75 ;
      RECT  3.565 1.415 3.685 1.75 ;
      RECT  4.085 1.415 4.205 1.75 ;
      RECT  4.605 1.415 4.725 1.75 ;
      RECT  5.135 1.415 5.255 1.75 ;
      RECT  5.73 1.415 5.85 1.75 ;
      RECT  6.315 1.42 6.435 1.75 ;
      RECT  6.835 1.445 6.955 1.75 ;
      RECT  7.355 1.45 7.475 1.75 ;
      RECT  7.875 1.45 7.995 1.75 ;
      RECT  8.63 1.43 8.75 1.75 ;
      RECT  9.15 1.43 9.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  8.67 0.05 8.79 0.36 ;
      RECT  6.135 0.05 6.255 0.365 ;
      RECT  6.655 0.05 6.775 0.365 ;
      RECT  1.115 0.05 1.235 0.385 ;
      RECT  7.62 0.05 7.74 0.385 ;
      RECT  8.145 0.05 8.265 0.385 ;
      RECT  2.34 0.05 2.46 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.76 0.51 3.45 0.69 ;
      RECT  3.35 0.69 3.45 1.11 ;
      RECT  2.75 1.11 6.695 1.29 ;
      RECT  2.75 1.29 2.905 1.39 ;
      RECT  6.55 1.29 6.695 1.49 ;
    END
    ANTENNADIFFAREA 0.984 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.285 0.19 1.02 0.32 ;
      RECT  1.51 0.2 2.245 0.32 ;
      RECT  2.55 0.215 4.72 0.335 ;
      RECT  4.605 0.335 4.72 0.385 ;
      RECT  2.55 0.335 2.65 0.51 ;
      RECT  2.54 0.51 2.65 0.705 ;
      RECT  6.865 0.215 7.085 0.335 ;
      RECT  6.865 0.335 6.985 0.455 ;
      RECT  4.81 0.2 5.995 0.32 ;
      RECT  5.875 0.32 5.995 0.455 ;
      RECT  5.875 0.455 6.985 0.575 ;
      RECT  8.93 0.35 9.05 0.45 ;
      RECT  8.36 0.45 9.05 0.57 ;
      RECT  0.075 0.4 0.195 0.5 ;
      RECT  0.075 0.5 0.84 0.62 ;
      RECT  0.74 0.62 0.84 1.22 ;
      RECT  0.075 1.22 1.235 1.34 ;
      RECT  0.075 1.34 0.195 1.44 ;
      RECT  1.115 1.34 1.235 1.44 ;
      RECT  3.77 0.475 5.785 0.595 ;
      RECT  7.31 0.475 8.05 0.595 ;
      RECT  7.1 0.495 7.21 0.74 ;
      RECT  6.225 0.74 7.21 0.84 ;
      RECT  7.095 0.84 7.21 1.24 ;
      RECT  7.095 1.24 8.255 1.36 ;
      RECT  8.135 1.36 8.255 1.63 ;
      RECT  3.55 0.505 3.65 0.835 ;
      RECT  3.55 0.835 4.37 0.95 ;
      RECT  5.06 0.83 6.005 0.93 ;
      RECT  5.06 0.93 6.96 0.95 ;
      RECT  5.87 0.95 6.96 1.02 ;
      RECT  6.86 1.02 6.96 1.32 ;
      RECT  2.56 0.83 3.225 0.95 ;
      RECT  2.56 0.95 2.65 1.24 ;
      RECT  1.25 0.5 2.05 0.62 ;
      RECT  1.94 0.62 2.05 1.24 ;
      RECT  1.585 1.24 2.65 1.36 ;
      RECT  8.345 1.11 8.445 1.22 ;
      RECT  8.345 1.22 9.535 1.34 ;
      RECT  9.415 0.46 9.535 1.22 ;
      LAYER M2 ;
      RECT  0.7 0.55 3.785 0.65 ;
      RECT  6.815 1.15 8.485 1.25 ;
      LAYER V1 ;
      RECT  0.74 0.55 0.84 0.65 ;
      RECT  3.55 0.55 3.65 0.65 ;
      RECT  6.86 1.15 6.96 1.25 ;
      RECT  8.345 1.15 8.445 1.25 ;
  END
END SEN_AO2222_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO222_1
#      Description : "Three 2-input ANDs into 3-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)|(C1&C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO222_1
  CLASS CORE ;
  FOREIGN SEN_AO222_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.82 ;
      RECT  0.265 0.82 0.45 0.99 ;
      RECT  0.35 0.99 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 0.935 ;
      RECT  0.545 0.935 0.65 1.105 ;
      RECT  0.55 1.105 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.86 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 0.71 ;
      RECT  2.55 0.71 2.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.46 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.38 0.185 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.595 1.395 0.715 1.75 ;
      RECT  1.11 1.605 1.28 1.75 ;
      RECT  1.63 1.6 1.8 1.75 ;
      RECT  2.175 1.6 2.345 1.75 ;
      RECT  2.73 1.41 2.87 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  0.595 0.05 0.715 0.225 ;
      RECT  2.185 0.05 2.305 0.355 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.32 0.22 2.05 0.34 ;
      RECT  1.94 0.34 2.05 1.315 ;
      RECT  1.35 1.315 2.05 1.49 ;
    END
    ANTENNADIFFAREA 0.271 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.425 0.245 2.9 0.355 ;
      RECT  2.425 0.355 2.515 0.445 ;
      RECT  2.14 0.445 2.515 0.565 ;
      RECT  2.14 0.565 2.23 1.39 ;
      RECT  2.14 1.39 2.64 1.51 ;
      RECT  0.065 0.315 1.03 0.405 ;
      RECT  0.94 0.405 1.03 0.645 ;
      RECT  0.065 0.405 0.175 1.18 ;
      RECT  0.94 0.645 1.6 0.735 ;
      RECT  1.5 0.735 1.6 1.0 ;
      RECT  0.065 1.18 0.445 1.285 ;
      RECT  0.325 1.285 0.445 1.485 ;
      RECT  1.12 0.3 1.225 0.465 ;
      RECT  1.12 0.465 1.825 0.555 ;
      RECT  1.735 0.555 1.825 1.135 ;
      RECT  1.17 1.135 1.825 1.225 ;
      RECT  1.17 1.225 1.26 1.38 ;
      RECT  0.805 1.38 1.26 1.49 ;
  END
END SEN_AO222_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO222_2
#      Description : "Three 2-input ANDs into 3-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)|(C1&C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO222_2
  CLASS CORE ;
  FOREIGN SEN_AO222_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0786 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.75 0.91 1.05 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0786 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0786 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 0.91 ;
      RECT  4.285 0.91 4.65 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0786 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.91 4.05 1.145 ;
      RECT  3.95 1.145 4.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0786 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0786 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.345 0.185 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.56 1.47 0.73 1.75 ;
      RECT  1.08 1.47 1.25 1.75 ;
      RECT  1.715 1.38 1.835 1.75 ;
      RECT  2.325 1.38 2.445 1.75 ;
      RECT  2.92 1.445 3.09 1.75 ;
      RECT  3.44 1.445 3.61 1.75 ;
      RECT  3.985 1.38 4.105 1.75 ;
      RECT  4.48 1.445 4.65 1.75 ;
      RECT  5.025 1.39 5.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  3.42 0.05 3.59 0.2 ;
      RECT  2.39 0.05 2.56 0.205 ;
      RECT  2.945 0.05 3.06 0.385 ;
      RECT  4.225 0.05 4.355 0.395 ;
      RECT  0.845 0.05 0.96 0.58 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.46 0.68 ;
      RECT  1.35 0.68 1.45 1.11 ;
      RECT  1.35 1.11 2.85 1.29 ;
    END
    ANTENNADIFFAREA 0.396 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.945 0.205 2.065 0.295 ;
      RECT  1.945 0.295 2.855 0.415 ;
      RECT  0.065 0.195 0.755 0.31 ;
      RECT  0.065 0.31 0.185 0.4 ;
      RECT  4.455 0.2 5.145 0.32 ;
      RECT  5.025 0.32 5.145 0.415 ;
      RECT  1.05 0.235 1.78 0.355 ;
      RECT  1.66 0.355 1.78 0.525 ;
      RECT  1.66 0.525 2.375 0.645 ;
      RECT  3.15 0.29 3.885 0.415 ;
      RECT  4.76 0.41 4.885 0.505 ;
      RECT  2.5 0.505 4.885 0.58 ;
      RECT  2.5 0.58 4.86 0.595 ;
      RECT  2.5 0.595 2.6 0.82 ;
      RECT  4.76 0.595 4.86 1.25 ;
      RECT  1.965 0.82 2.6 0.94 ;
      RECT  4.195 1.25 4.86 1.355 ;
      RECT  4.74 1.355 4.86 1.37 ;
      RECT  4.74 1.37 4.885 1.54 ;
      RECT  3.55 0.715 4.13 0.82 ;
      RECT  3.55 0.82 3.64 1.225 ;
      RECT  2.72 0.775 3.04 0.975 ;
      RECT  2.95 0.975 3.04 1.225 ;
      RECT  2.95 1.225 3.64 1.24 ;
      RECT  2.95 1.24 3.845 1.355 ;
      RECT  3.725 1.355 3.845 1.475 ;
      RECT  0.34 0.4 0.43 1.265 ;
      RECT  0.34 1.265 1.245 1.38 ;
      RECT  1.155 0.75 1.245 1.265 ;
      RECT  0.34 1.38 0.445 1.505 ;
  END
END SEN_AO222_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO222_4
#      Description : "Three 2-input ANDs into 3-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)|(C1&C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO222_4
  CLASS CORE ;
  FOREIGN SEN_AO222_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.925 ;
      RECT  0.15 0.925 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1548 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 0.91 ;
      RECT  0.95 0.91 1.45 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1536 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.25 0.91 ;
      RECT  6.95 0.91 7.25 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1536 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.55 0.705 7.65 0.9 ;
      RECT  7.55 0.9 7.905 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1548 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.71 5.85 0.91 ;
      RECT  5.35 0.91 5.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1536 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.03 0.89 6.65 1.09 ;
      RECT  6.55 1.09 6.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1548 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.56 1.465 0.73 1.75 ;
      RECT  1.08 1.465 1.25 1.75 ;
      RECT  1.625 1.45 1.745 1.75 ;
      RECT  2.145 1.425 2.265 1.75 ;
      RECT  2.665 1.425 2.785 1.75 ;
      RECT  3.185 1.425 3.305 1.75 ;
      RECT  3.765 1.425 3.885 1.75 ;
      RECT  4.335 1.415 4.455 1.75 ;
      RECT  4.895 1.2 5.015 1.75 ;
      RECT  5.415 1.415 5.535 1.75 ;
      RECT  5.935 1.415 6.055 1.75 ;
      RECT  6.455 1.45 6.575 1.75 ;
      RECT  6.95 1.475 7.12 1.75 ;
      RECT  7.47 1.475 7.64 1.75 ;
      RECT  8.015 1.21 8.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  4.06 0.05 4.23 0.2 ;
      RECT  4.6 0.05 4.77 0.2 ;
      RECT  5.89 0.05 6.06 0.2 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  7.495 0.05 7.615 0.36 ;
      RECT  6.455 0.05 6.575 0.38 ;
      RECT  8.015 0.05 8.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 2.65 0.69 ;
      RECT  2.55 0.69 2.65 1.11 ;
      RECT  1.885 1.11 4.715 1.29 ;
      RECT  1.885 1.29 2.05 1.49 ;
      RECT  4.55 1.29 4.715 1.49 ;
    END
    ANTENNADIFFAREA 0.812 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.895 0.185 5.015 0.29 ;
      RECT  3.875 0.29 5.015 0.41 ;
      RECT  3.875 0.41 3.995 0.565 ;
      RECT  2.795 0.565 3.995 0.685 ;
      RECT  5.125 0.19 5.765 0.29 ;
      RECT  5.125 0.29 6.34 0.36 ;
      RECT  5.645 0.36 6.34 0.41 ;
      RECT  0.275 0.2 1.01 0.32 ;
      RECT  0.92 0.32 1.01 0.475 ;
      RECT  0.92 0.475 1.485 0.595 ;
      RECT  1.365 0.595 1.485 0.81 ;
      RECT  6.69 0.215 7.355 0.335 ;
      RECT  7.235 0.335 7.355 0.475 ;
      RECT  7.235 0.475 7.925 0.595 ;
      RECT  1.5 0.235 3.785 0.355 ;
      RECT  4.15 0.5 7.12 0.62 ;
      RECT  4.15 0.62 4.25 0.82 ;
      RECT  6.74 0.62 6.84 1.265 ;
      RECT  2.985 0.82 4.25 0.94 ;
      RECT  6.74 1.265 7.925 1.385 ;
      RECT  6.715 1.385 6.84 1.57 ;
      RECT  5.13 0.71 5.555 0.82 ;
      RECT  4.415 0.82 5.23 0.94 ;
      RECT  5.13 0.94 5.23 1.2 ;
      RECT  5.13 1.2 6.365 1.32 ;
      RECT  1.66 0.82 2.305 0.94 ;
      RECT  1.66 0.94 1.76 1.23 ;
      RECT  0.065 0.31 0.185 0.41 ;
      RECT  0.065 0.41 0.83 0.53 ;
      RECT  0.74 0.53 0.83 1.23 ;
      RECT  0.275 1.23 1.76 1.35 ;
  END
END SEN_AO222_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO222_6
#      Description : "Three 2-input ANDs into 3-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)|(C1&C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO222_6
  CLASS CORE ;
  FOREIGN SEN_AO222_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.715 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.15 0.91 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.75 0.71 10.85 0.87 ;
      RECT  10.455 0.87 10.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.35 0.71 9.45 0.91 ;
      RECT  9.35 0.91 9.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 7.85 0.925 ;
      RECT  7.75 0.925 7.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.71 8.65 0.92 ;
      RECT  8.55 0.92 8.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 11.2 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  1.105 1.415 1.225 1.75 ;
      RECT  1.625 1.415 1.745 1.75 ;
      RECT  2.145 1.2 2.26 1.75 ;
      RECT  2.665 1.38 2.785 1.75 ;
      RECT  3.185 1.39 3.305 1.75 ;
      RECT  3.705 1.39 3.825 1.75 ;
      RECT  4.225 1.39 4.345 1.75 ;
      RECT  4.745 1.39 4.865 1.75 ;
      RECT  5.265 1.395 5.385 1.75 ;
      RECT  5.785 1.395 5.905 1.75 ;
      RECT  6.305 1.395 6.425 1.75 ;
      RECT  6.825 1.2 6.945 1.75 ;
      RECT  7.345 1.405 7.465 1.75 ;
      RECT  7.865 1.405 7.985 1.75 ;
      RECT  8.385 1.405 8.505 1.75 ;
      RECT  8.905 1.2 9.025 1.75 ;
      RECT  9.425 1.415 9.545 1.75 ;
      RECT  9.945 1.415 10.065 1.75 ;
      RECT  10.465 1.415 10.585 1.75 ;
      RECT  11.0 1.21 11.12 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.2 0.05 ;
      RECT  5.535 0.05 5.655 0.36 ;
      RECT  6.055 0.05 6.175 0.36 ;
      RECT  8.125 0.05 8.245 0.36 ;
      RECT  8.645 0.05 8.765 0.36 ;
      RECT  9.685 0.05 9.805 0.36 ;
      RECT  1.375 0.05 1.495 0.385 ;
      RECT  1.895 0.05 2.015 0.575 ;
      RECT  9.165 0.05 9.285 0.575 ;
      RECT  6.575 0.05 6.695 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 3.85 0.69 ;
      RECT  3.72 0.69 3.85 1.1 ;
      RECT  3.72 1.1 6.685 1.105 ;
      RECT  2.35 1.105 6.685 1.29 ;
    END
    ANTENNADIFFAREA 1.186 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.105 0.215 4.9 0.335 ;
      RECT  6.8 0.215 7.985 0.335 ;
      RECT  7.865 0.335 7.985 0.45 ;
      RECT  7.865 0.45 9.075 0.57 ;
      RECT  9.945 0.215 11.105 0.335 ;
      RECT  10.985 0.335 11.105 0.44 ;
      RECT  9.945 0.335 10.065 0.475 ;
      RECT  9.4 0.475 10.065 0.595 ;
      RECT  0.065 0.23 1.225 0.35 ;
      RECT  0.065 0.35 0.185 0.46 ;
      RECT  1.105 0.35 1.225 0.475 ;
      RECT  1.105 0.475 1.805 0.595 ;
      RECT  3.95 0.475 6.46 0.595 ;
      RECT  7.06 0.475 7.75 0.595 ;
      RECT  7.06 0.595 7.165 0.88 ;
      RECT  5.835 0.88 7.165 1.005 ;
      RECT  7.06 1.005 7.165 1.19 ;
      RECT  7.06 1.19 8.815 1.31 ;
      RECT  10.16 0.475 10.895 0.595 ;
      RECT  10.16 0.595 10.26 1.205 ;
      RECT  9.14 1.205 10.895 1.325 ;
      RECT  6.845 0.49 6.945 0.685 ;
      RECT  5.555 0.685 6.945 0.775 ;
      RECT  5.555 0.775 5.655 0.875 ;
      RECT  4.235 0.875 5.655 1.005 ;
      RECT  1.965 0.79 3.31 0.91 ;
      RECT  1.965 0.91 2.055 1.18 ;
      RECT  0.275 0.45 0.99 0.57 ;
      RECT  0.9 0.57 0.99 1.18 ;
      RECT  0.275 1.18 2.055 1.3 ;
      LAYER M2 ;
      RECT  6.795 0.55 10.3 0.65 ;
      LAYER V1 ;
      RECT  6.845 0.55 6.945 0.65 ;
      RECT  10.16 0.55 10.26 0.65 ;
  END
END SEN_AO222_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_1
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_1
  CLASS CORE ;
  FOREIGN SEN_AO22_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.47 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.355 1.44 1.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.23 0.05 1.35 0.35 ;
      RECT  0.065 0.05 0.185 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.735 0.49 ;
      RECT  1.55 0.49 1.65 1.31 ;
      RECT  1.55 1.31 1.73 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.56 0.24 1.14 0.36 ;
      RECT  1.05 0.36 1.14 0.44 ;
      RECT  1.05 0.44 1.46 0.56 ;
      RECT  1.37 0.56 1.46 1.24 ;
      RECT  0.82 1.24 1.46 1.35 ;
      RECT  0.065 1.21 0.71 1.305 ;
      RECT  0.065 1.305 0.185 1.43 ;
      RECT  0.58 1.305 0.71 1.445 ;
      RECT  0.58 1.445 1.25 1.56 ;
  END
END SEN_AO22_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_2
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_2
  CLASS CORE ;
  FOREIGN SEN_AO22_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.345 1.45 0.465 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.905 1.45 1.025 1.75 ;
      RECT  2.66 1.44 2.78 1.75 ;
      RECT  3.21 1.21 3.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  2.11 0.05 2.28 0.21 ;
      RECT  0.345 0.05 0.465 0.35 ;
      RECT  2.68 0.05 2.8 0.59 ;
      RECT  3.21 0.05 3.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.31 3.05 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.615 0.17 1.735 0.3 ;
      RECT  1.615 0.3 2.54 0.39 ;
      RECT  2.42 0.17 2.54 0.3 ;
      RECT  0.81 0.24 1.48 0.355 ;
      RECT  1.36 0.355 1.48 0.485 ;
      RECT  1.36 0.485 2.02 0.605 ;
      RECT  1.93 0.605 2.02 1.24 ;
      RECT  1.48 1.24 2.86 1.35 ;
      RECT  2.77 0.71 2.86 1.24 ;
      RECT  0.085 0.34 0.205 0.445 ;
      RECT  0.085 0.445 1.27 0.56 ;
      RECT  0.085 1.24 1.34 1.36 ;
      RECT  1.22 1.36 1.34 1.44 ;
      RECT  0.085 1.36 0.205 1.46 ;
      RECT  1.22 1.44 2.49 1.56 ;
  END
END SEN_AO22_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_4
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_4
  CLASS CORE ;
  FOREIGN SEN_AO22_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.45 0.45 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.85 1.45 0.97 1.75 ;
      RECT  1.37 1.45 1.49 1.75 ;
      RECT  1.89 1.45 2.01 1.75 ;
      RECT  4.76 1.2 4.88 1.75 ;
      RECT  5.28 1.425 5.4 1.75 ;
      RECT  5.815 1.21 5.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  3.67 0.05 3.84 0.21 ;
      RECT  0.33 0.05 0.45 0.36 ;
      RECT  0.85 0.05 0.97 0.36 ;
      RECT  4.24 0.05 4.36 0.38 ;
      RECT  5.28 0.05 5.4 0.385 ;
      RECT  5.815 0.05 5.935 0.59 ;
      RECT  4.76 0.05 4.88 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.02 0.51 5.65 0.69 ;
      RECT  5.55 0.69 5.65 1.11 ;
      RECT  5.03 1.11 5.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.635 0.3 4.1 0.42 ;
      RECT  3.98 0.42 4.1 0.47 ;
      RECT  3.98 0.47 4.645 0.59 ;
      RECT  0.07 0.34 0.19 0.45 ;
      RECT  0.07 0.45 2.295 0.56 ;
      RECT  4.56 0.79 5.415 0.89 ;
      RECT  4.56 0.89 4.65 1.24 ;
      RECT  1.345 0.24 2.525 0.36 ;
      RECT  2.4 0.36 2.525 0.51 ;
      RECT  2.4 0.51 3.65 0.62 ;
      RECT  3.56 0.62 3.65 1.24 ;
      RECT  2.6 1.24 4.65 1.355 ;
      RECT  0.07 1.24 2.395 1.36 ;
      RECT  2.27 1.36 2.395 1.445 ;
      RECT  0.07 1.36 0.19 1.46 ;
      RECT  2.27 1.445 4.655 1.56 ;
  END
END SEN_AO22_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_DG_1
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_DG_1
  CLASS CORE ;
  FOREIGN SEN_AO22_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.14 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.4 0.45 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.355 1.41 1.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  1.2 0.05 1.33 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.65 1.235 ;
      RECT  1.55 1.235 1.735 1.49 ;
    END
    ANTENNADIFFAREA 0.182 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.54 0.25 1.05 0.37 ;
      RECT  0.95 0.37 1.05 0.495 ;
      RECT  0.95 0.495 1.46 0.585 ;
      RECT  1.35 0.585 1.46 0.955 ;
      RECT  0.95 0.585 1.05 1.23 ;
      RECT  0.845 1.23 1.05 1.32 ;
      RECT  0.845 1.32 0.965 1.48 ;
      RECT  0.065 1.21 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.55 ;
      RECT  0.585 1.305 0.705 1.57 ;
      RECT  0.585 1.57 1.225 1.66 ;
      RECT  1.105 1.395 1.225 1.57 ;
  END
END SEN_AO22_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_DG_10
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_DG_10
  CLASS CORE ;
  FOREIGN SEN_AO22_DG_10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.45 0.9 ;
      RECT  2.35 0.9 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.05 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  3.39 1.01 3.56 1.29 ;
      RECT  3.44 1.29 3.56 1.75 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  3.905 1.41 4.035 1.75 ;
      RECT  4.425 1.41 4.555 1.75 ;
      RECT  4.945 1.41 5.075 1.75 ;
      RECT  5.465 1.41 5.595 1.75 ;
      RECT  6.015 1.21 6.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  2.68 0.05 2.85 0.19 ;
      RECT  0.56 0.05 0.73 0.365 ;
      RECT  3.905 0.05 4.035 0.39 ;
      RECT  4.425 0.05 4.555 0.39 ;
      RECT  4.945 0.05 5.075 0.39 ;
      RECT  5.465 0.05 5.595 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.015 0.05 6.135 0.59 ;
      RECT  3.37 0.05 3.49 0.665 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.6 0.505 5.855 0.69 ;
      RECT  5.43 0.69 5.65 1.11 ;
      RECT  3.65 1.11 5.85 1.29 ;
    END
    ANTENNADIFFAREA 1.108 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.245 1.54 0.365 ;
      RECT  0.845 0.365 0.965 0.465 ;
      RECT  0.3 0.465 0.965 0.585 ;
      RECT  1.83 0.28 3.18 0.4 ;
      RECT  1.08 0.49 3.27 0.61 ;
      RECT  3.15 0.61 3.27 0.785 ;
      RECT  3.15 0.785 5.32 0.9 ;
      RECT  3.15 0.9 3.27 1.23 ;
      RECT  1.835 1.23 3.27 1.35 ;
      RECT  0.065 1.23 1.745 1.35 ;
      RECT  0.065 1.35 0.185 1.45 ;
      RECT  1.625 1.35 1.745 1.465 ;
      RECT  1.625 1.465 3.35 1.585 ;
  END
END SEN_AO22_DG_10
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_DG_2
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_DG_2
  CLASS CORE ;
  FOREIGN SEN_AO22_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.14 0.71 1.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.4 0.45 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.305 1.19 1.41 1.75 ;
      RECT  1.81 1.21 1.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  1.22 0.05 1.35 0.39 ;
      RECT  1.81 0.05 1.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.67 0.585 ;
      RECT  1.55 0.585 1.65 1.235 ;
      RECT  1.55 1.235 1.67 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.54 0.26 1.05 0.38 ;
      RECT  0.95 0.38 1.05 0.51 ;
      RECT  0.95 0.51 1.46 0.6 ;
      RECT  1.35 0.6 1.46 0.955 ;
      RECT  0.95 0.6 1.05 1.23 ;
      RECT  0.845 1.23 1.05 1.32 ;
      RECT  0.845 1.32 0.965 1.48 ;
      RECT  0.065 1.21 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.53 ;
      RECT  0.585 1.305 0.705 1.57 ;
      RECT  0.585 1.57 1.215 1.66 ;
      RECT  1.105 1.41 1.215 1.57 ;
  END
END SEN_AO22_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_DG_3
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_DG_3
  CLASS CORE ;
  FOREIGN SEN_AO22_DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.4 0.45 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.355 1.21 1.475 1.75 ;
      RECT  1.87 1.41 2.0 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  1.265 0.05 1.395 0.39 ;
      RECT  1.87 0.05 2.0 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.615 0.51 2.25 0.69 ;
      RECT  2.135 0.69 2.25 1.11 ;
      RECT  1.615 1.11 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.54 0.27 1.05 0.39 ;
      RECT  0.95 0.39 1.05 0.51 ;
      RECT  0.95 0.51 1.51 0.6 ;
      RECT  1.4 0.6 1.51 0.785 ;
      RECT  0.95 0.6 1.05 1.23 ;
      RECT  1.4 0.785 2.02 0.895 ;
      RECT  0.845 1.23 1.05 1.32 ;
      RECT  0.845 1.32 0.965 1.45 ;
      RECT  0.065 1.21 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.43 ;
      RECT  0.585 1.305 0.705 1.57 ;
      RECT  0.585 1.57 1.225 1.66 ;
      RECT  1.105 1.395 1.225 1.57 ;
  END
END SEN_AO22_DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_DG_4
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_DG_4
  CLASS CORE ;
  FOREIGN SEN_AO22_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.4 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.355 1.21 1.475 1.75 ;
      RECT  1.87 1.41 2.0 1.75 ;
      RECT  2.405 1.215 2.525 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  1.87 0.05 2.0 0.39 ;
      RECT  1.265 0.05 1.395 0.405 ;
      RECT  2.405 0.05 2.525 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.615 0.51 2.25 0.69 ;
      RECT  2.135 0.69 2.25 1.11 ;
      RECT  1.615 1.11 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.56 0.28 1.05 0.4 ;
      RECT  0.95 0.4 1.05 0.51 ;
      RECT  0.95 0.51 1.51 0.6 ;
      RECT  1.4 0.6 1.51 0.785 ;
      RECT  0.95 0.6 1.05 1.23 ;
      RECT  1.4 0.785 2.02 0.895 ;
      RECT  0.845 1.23 1.05 1.32 ;
      RECT  0.845 1.32 0.965 1.45 ;
      RECT  0.065 1.21 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.43 ;
      RECT  0.585 1.305 0.705 1.57 ;
      RECT  0.585 1.57 1.225 1.66 ;
      RECT  1.105 1.41 1.225 1.57 ;
  END
END SEN_AO22_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_DG_8
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_DG_8
  CLASS CORE ;
  FOREIGN SEN_AO22_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  1.15 0.91 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.45 0.91 ;
      RECT  2.1 0.91 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  2.695 1.435 2.865 1.75 ;
      RECT  3.235 1.39 3.365 1.75 ;
      RECT  3.755 1.39 3.885 1.75 ;
      RECT  4.275 1.39 4.405 1.75 ;
      RECT  4.81 1.21 4.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  2.16 0.05 2.33 0.305 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  3.235 0.05 3.365 0.41 ;
      RECT  3.755 0.05 3.885 0.41 ;
      RECT  4.275 0.05 4.405 0.41 ;
      RECT  2.72 0.05 2.84 0.57 ;
      RECT  4.81 0.05 4.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.51 4.665 0.69 ;
      RECT  4.495 0.69 4.665 1.11 ;
      RECT  2.95 1.11 4.665 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.215 1.27 0.335 ;
      RECT  0.585 0.335 0.705 0.5 ;
      RECT  0.065 0.4 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.62 ;
      RECT  1.36 0.24 2.045 0.36 ;
      RECT  1.925 0.36 2.045 0.4 ;
      RECT  1.925 0.4 2.59 0.52 ;
      RECT  2.615 0.785 4.285 0.905 ;
      RECT  2.615 0.905 2.735 1.215 ;
      RECT  0.82 0.45 1.8 0.57 ;
      RECT  1.68 0.57 1.8 1.215 ;
      RECT  1.34 1.215 2.735 1.335 ;
      RECT  0.065 1.205 1.225 1.325 ;
      RECT  0.065 1.325 0.185 1.43 ;
      RECT  1.105 1.325 1.225 1.445 ;
      RECT  1.105 1.445 2.35 1.565 ;
  END
END SEN_AO22_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AO22_8
#      Description : "Two 2-input ANDs into 2-input OR"
#      Equation    : X=(A1&A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO22_8
  CLASS CORE ;
  FOREIGN SEN_AO22_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.95 0.71 10.65 0.925 ;
      RECT  9.95 0.925 10.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3378 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.35 0.71 9.05 0.91 ;
      RECT  8.95 0.91 9.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3378 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.25 0.925 ;
      RECT  0.55 0.925 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3378 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.85 0.925 ;
      RECT  2.15 0.925 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3378 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.18 1.75 ;
      RECT  0.0 1.75 11.0 1.85 ;
      RECT  0.57 1.415 0.7 1.75 ;
      RECT  1.09 1.415 1.22 1.75 ;
      RECT  1.61 1.415 1.74 1.75 ;
      RECT  2.13 1.415 2.26 1.75 ;
      RECT  2.65 1.415 2.78 1.75 ;
      RECT  3.28 1.415 3.41 1.75 ;
      RECT  3.875 1.41 4.005 1.75 ;
      RECT  4.395 1.41 4.525 1.75 ;
      RECT  4.915 1.41 5.045 1.75 ;
      RECT  5.435 1.41 5.565 1.75 ;
      RECT  5.955 1.41 6.085 1.75 ;
      RECT  6.475 1.41 6.605 1.75 ;
      RECT  6.995 1.41 7.125 1.75 ;
      RECT  7.61 1.21 7.73 1.75 ;
      RECT  8.22 1.41 8.35 1.75 ;
      RECT  8.74 1.41 8.87 1.75 ;
      RECT  9.26 1.41 9.39 1.75 ;
      RECT  9.78 1.41 9.91 1.75 ;
      RECT  10.3 1.41 10.43 1.75 ;
      RECT  10.82 1.41 10.945 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      RECT  3.615 0.05 3.745 0.36 ;
      RECT  4.135 0.05 4.265 0.36 ;
      RECT  4.655 0.05 4.785 0.36 ;
      RECT  5.175 0.05 5.305 0.36 ;
      RECT  1.87 0.05 2.0 0.385 ;
      RECT  2.39 0.05 2.52 0.385 ;
      RECT  2.91 0.05 3.04 0.385 ;
      RECT  7.96 0.05 8.09 0.39 ;
      RECT  8.48 0.05 8.61 0.39 ;
      RECT  9.0 0.05 9.13 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.7 0.51 7.45 0.69 ;
      RECT  5.905 0.69 6.075 1.11 ;
      RECT  3.635 1.11 7.45 1.29 ;
    END
    ANTENNADIFFAREA 1.264 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.2 1.735 0.32 ;
      RECT  0.055 0.32 0.175 0.42 ;
      RECT  1.615 0.32 1.735 0.475 ;
      RECT  1.615 0.475 3.28 0.595 ;
      RECT  3.175 0.595 3.28 0.69 ;
      RECT  9.265 0.215 10.945 0.335 ;
      RECT  10.825 0.335 10.945 0.42 ;
      RECT  9.265 0.335 9.385 0.5 ;
      RECT  7.65 0.5 9.385 0.62 ;
      RECT  5.415 0.23 7.69 0.38 ;
      RECT  5.415 0.38 5.585 0.45 ;
      RECT  3.37 0.18 3.48 0.45 ;
      RECT  3.37 0.45 5.585 0.62 ;
      RECT  9.5 0.475 10.74 0.595 ;
      RECT  9.5 0.595 9.59 1.18 ;
      RECT  6.165 0.805 8.03 0.93 ;
      RECT  7.91 0.93 8.03 1.18 ;
      RECT  7.91 1.18 10.74 1.3 ;
      RECT  3.395 0.8 5.05 0.93 ;
      RECT  3.395 0.93 3.515 1.205 ;
      RECT  0.29 0.475 1.505 0.595 ;
      RECT  1.415 0.595 1.505 1.205 ;
      RECT  0.26 1.205 3.515 1.325 ;
  END
END SEN_AO22_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_0P5
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_0P5
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.675 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.49 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.525 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.585 1.41 0.715 1.75 ;
      RECT  1.435 1.41 1.565 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.095 0.05 1.265 0.185 ;
      RECT  0.585 0.05 0.71 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.21 1.735 0.38 ;
      RECT  1.55 0.38 1.65 1.22 ;
      RECT  1.15 1.22 1.65 1.31 ;
      RECT  1.15 1.31 1.25 1.53 ;
    END
    ANTENNADIFFAREA 0.112 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.18 0.19 0.27 ;
      RECT  0.07 0.27 0.435 0.39 ;
      RECT  0.345 0.39 0.435 0.485 ;
      RECT  0.345 0.485 1.445 0.575 ;
      RECT  1.355 0.575 1.445 0.985 ;
      RECT  0.345 0.575 0.435 1.63 ;
      RECT  1.355 0.2 1.46 0.275 ;
      RECT  0.8 0.275 1.46 0.395 ;
  END
END SEN_AO2BB2_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_1
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_1
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.14 0.67 1.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0408 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.525 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0408 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.62 1.4 0.74 1.75 ;
      RECT  1.565 1.6 1.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.105 0.05 1.225 0.37 ;
      RECT  0.58 0.05 0.71 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.735 0.49 ;
      RECT  1.55 0.49 1.65 1.38 ;
      RECT  1.18 1.38 1.65 1.5 ;
    END
    ANTENNADIFFAREA 0.207 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 1.2 ;
      RECT  0.34 1.2 1.46 1.29 ;
      RECT  1.35 0.72 1.46 1.2 ;
      RECT  0.34 1.29 0.445 1.49 ;
      RECT  1.355 0.36 1.46 0.46 ;
      RECT  0.795 0.46 1.46 0.58 ;
  END
END SEN_AO2BB2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_2
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_2
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.65 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.05 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0816 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0816 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.56 1.48 0.73 1.75 ;
      RECT  1.1 1.48 1.27 1.75 ;
      RECT  1.665 1.24 1.785 1.75 ;
      RECT  2.725 1.4 2.845 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  2.185 0.05 2.305 0.38 ;
      RECT  2.725 0.05 2.845 0.38 ;
      RECT  0.325 0.05 0.445 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.585 0.44 1.85 0.56 ;
      RECT  1.75 0.56 1.85 1.025 ;
      RECT  1.35 1.025 2.29 1.145 ;
      RECT  1.35 1.145 1.51 1.29 ;
      RECT  2.15 1.145 2.29 1.29 ;
    END
    ANTENNADIFFAREA 0.334 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.215 1.25 0.335 ;
      RECT  0.585 0.335 0.705 0.5 ;
      RECT  0.065 0.33 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.59 ;
      RECT  1.355 0.26 2.045 0.35 ;
      RECT  1.94 0.35 2.045 0.47 ;
      RECT  1.355 0.35 1.475 0.48 ;
      RECT  1.94 0.47 3.13 0.59 ;
      RECT  3.01 0.37 3.13 0.47 ;
      RECT  0.815 0.43 1.25 0.55 ;
      RECT  1.14 0.55 1.25 0.79 ;
      RECT  1.14 0.79 1.66 0.89 ;
      RECT  1.14 0.89 1.25 1.27 ;
      RECT  0.285 1.27 1.25 1.39 ;
      RECT  2.445 1.18 3.13 1.3 ;
      RECT  3.01 1.3 3.13 1.42 ;
      RECT  2.445 1.3 2.565 1.445 ;
      RECT  1.925 1.35 2.045 1.445 ;
      RECT  1.925 1.445 2.565 1.57 ;
  END
END SEN_AO2BB2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_4
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_4
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.85 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 4.85 0.89 ;
      RECT  4.75 0.89 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1629 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1629 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.59 1.415 0.71 1.75 ;
      RECT  1.11 1.415 1.23 1.75 ;
      RECT  1.63 1.415 1.75 1.75 ;
      RECT  2.15 1.415 2.27 1.75 ;
      RECT  2.67 1.415 2.79 1.75 ;
      RECT  4.23 1.415 4.35 1.75 ;
      RECT  4.75 1.42 4.87 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  0.59 0.05 0.71 0.375 ;
      RECT  3.19 0.05 3.31 0.38 ;
      RECT  3.71 0.05 3.83 0.38 ;
      RECT  4.23 0.05 4.35 0.38 ;
      RECT  4.75 0.05 4.87 0.38 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.85 0.69 ;
      RECT  2.75 0.69 2.85 1.11 ;
      RECT  1.89 1.11 3.65 1.18 ;
      RECT  1.89 1.18 3.855 1.29 ;
    END
    ANTENNADIFFAREA 0.668 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.23 1.515 0.35 ;
      RECT  0.845 0.35 0.975 0.465 ;
      RECT  0.29 0.465 0.975 0.59 ;
      RECT  1.855 0.24 3.05 0.36 ;
      RECT  2.94 0.36 3.05 0.47 ;
      RECT  2.94 0.47 5.13 0.59 ;
      RECT  5.01 0.37 5.13 0.47 ;
      RECT  1.085 0.44 1.78 0.56 ;
      RECT  1.67 0.56 1.78 0.79 ;
      RECT  1.67 0.79 2.4 0.89 ;
      RECT  1.67 0.89 1.78 1.205 ;
      RECT  0.3 1.205 1.78 1.325 ;
      RECT  3.97 1.18 5.13 1.3 ;
      RECT  5.01 1.3 5.13 1.42 ;
      RECT  3.97 1.3 4.09 1.45 ;
      RECT  2.905 1.45 4.09 1.57 ;
  END
END SEN_AO2BB2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_8
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_8
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 6.05 0.89 ;
      RECT  5.95 0.89 6.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.71 8.05 0.89 ;
      RECT  7.95 0.89 8.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2232 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.985 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2232 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.24 1.21 0.36 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.845 1.45 0.975 1.75 ;
      RECT  1.365 1.45 1.495 1.75 ;
      RECT  1.99 1.45 2.12 1.75 ;
      RECT  2.62 1.41 2.75 1.75 ;
      RECT  3.14 1.41 3.27 1.75 ;
      RECT  3.66 1.41 3.79 1.75 ;
      RECT  4.18 1.44 4.31 1.75 ;
      RECT  6.775 1.255 6.895 1.75 ;
      RECT  7.295 1.255 7.415 1.75 ;
      RECT  7.815 1.425 7.945 1.75 ;
      RECT  8.34 1.425 8.47 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  4.69 0.05 4.82 0.345 ;
      RECT  5.21 0.05 5.34 0.345 ;
      RECT  5.73 0.05 5.86 0.345 ;
      RECT  6.25 0.05 6.38 0.345 ;
      RECT  6.77 0.05 6.9 0.345 ;
      RECT  7.29 0.05 7.42 0.345 ;
      RECT  7.815 0.05 7.945 0.345 ;
      RECT  8.34 0.05 8.47 0.345 ;
      RECT  0.325 0.05 0.455 0.35 ;
      RECT  0.845 0.05 0.975 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.59 0.435 4.32 0.56 ;
      RECT  4.08 0.56 4.25 1.11 ;
      RECT  2.35 1.11 5.85 1.225 ;
      RECT  2.35 1.225 6.4 1.29 ;
      RECT  5.765 1.29 6.4 1.345 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.88 0.185 4.58 0.205 ;
      RECT  2.355 0.205 4.58 0.335 ;
      RECT  4.41 0.335 4.58 0.435 ;
      RECT  2.355 0.335 2.475 0.67 ;
      RECT  4.41 0.435 8.725 0.57 ;
      RECT  8.605 0.35 8.725 0.435 ;
      RECT  4.41 0.57 6.67 0.605 ;
      RECT  1.11 0.22 2.265 0.335 ;
      RECT  1.11 0.335 1.23 0.44 ;
      RECT  2.15 0.335 2.265 0.44 ;
      RECT  0.07 0.345 0.19 0.44 ;
      RECT  0.07 0.44 1.23 0.56 ;
      RECT  1.345 0.445 2.05 0.56 ;
      RECT  1.96 0.56 2.05 0.77 ;
      RECT  1.96 0.77 3.91 0.895 ;
      RECT  1.96 0.895 2.05 1.24 ;
      RECT  0.54 1.24 2.05 1.36 ;
      RECT  6.495 1.015 7.835 1.165 ;
      RECT  7.7 1.165 7.835 1.18 ;
      RECT  6.495 1.165 6.66 1.435 ;
      RECT  7.7 1.18 8.725 1.315 ;
      RECT  8.605 1.315 8.725 1.4 ;
      RECT  4.41 1.435 6.66 1.57 ;
      RECT  5.95 1.57 6.66 1.585 ;
  END
END SEN_AO2BB2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_DG_1
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_DG_1
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.63 0.85 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.645 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.51 0.65 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.41 0.21 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.61 1.44 0.74 1.75 ;
      RECT  1.43 1.54 1.62 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.55 0.05 0.68 0.36 ;
      RECT  1.095 0.05 1.225 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.215 1.73 0.385 ;
      RECT  1.55 0.385 1.65 1.36 ;
      RECT  1.105 1.36 1.65 1.45 ;
      RECT  1.105 1.45 1.225 1.58 ;
    END
    ANTENNADIFFAREA 0.197 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.84 0.32 0.96 0.45 ;
      RECT  0.84 0.45 1.46 0.54 ;
      RECT  1.35 0.32 1.46 0.45 ;
      RECT  1.355 0.725 1.445 1.18 ;
      RECT  0.925 1.18 1.445 1.26 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 1.26 ;
      RECT  0.34 1.26 1.445 1.27 ;
      RECT  0.34 1.27 1.015 1.35 ;
      RECT  0.34 1.35 0.465 1.59 ;
  END
END SEN_AO2BB2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_DG_2
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_DG_2
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.75 ;
      RECT  0.35 0.75 0.545 0.93 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.4 1.23 1.75 ;
      RECT  2.13 1.44 2.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.61 0.05 1.74 0.36 ;
      RECT  2.13 0.05 2.26 0.36 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.07 0.495 1.25 0.615 ;
      RECT  1.15 0.615 1.25 1.11 ;
      RECT  0.845 1.11 1.735 1.29 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.81 0.215 1.475 0.335 ;
      RECT  1.355 0.335 1.475 0.45 ;
      RECT  1.355 0.45 2.515 0.57 ;
      RECT  2.395 0.35 2.515 0.45 ;
      RECT  0.585 0.21 0.705 0.45 ;
      RECT  0.585 0.45 0.755 0.54 ;
      RECT  0.665 0.54 0.755 0.785 ;
      RECT  0.665 0.785 1.055 0.895 ;
      RECT  0.665 0.895 0.755 1.26 ;
      RECT  0.375 1.26 0.755 1.35 ;
      RECT  0.375 1.35 0.47 1.425 ;
      RECT  0.3 1.425 0.47 1.545 ;
      RECT  1.875 1.26 2.515 1.35 ;
      RECT  1.875 1.35 1.995 1.405 ;
      RECT  2.395 1.35 2.515 1.48 ;
      RECT  1.33 1.405 1.995 1.525 ;
  END
END SEN_AO2BB2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_DG_4
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_DG_4
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.85 0.895 ;
      RECT  3.75 0.895 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.755 ;
      RECT  0.35 0.755 0.535 0.925 ;
      RECT  0.35 0.925 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  3.17 1.44 3.3 1.75 ;
      RECT  3.69 1.44 3.82 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  2.13 0.05 2.26 0.36 ;
      RECT  2.65 0.05 2.78 0.36 ;
      RECT  3.17 0.05 3.3 0.36 ;
      RECT  3.69 0.05 3.82 0.36 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.045 0.475 1.85 0.595 ;
      RECT  1.75 0.595 1.85 1.11 ;
      RECT  0.845 1.11 2.795 1.29 ;
      RECT  0.845 1.29 0.965 1.56 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.785 0.265 2.03 0.385 ;
      RECT  1.94 0.385 2.03 0.45 ;
      RECT  1.94 0.45 4.12 0.57 ;
      RECT  0.54 0.475 0.755 0.595 ;
      RECT  0.665 0.595 0.755 0.785 ;
      RECT  0.665 0.785 1.44 0.895 ;
      RECT  0.665 0.895 0.755 1.23 ;
      RECT  0.3 1.23 0.755 1.35 ;
      RECT  2.915 1.23 4.12 1.35 ;
      RECT  2.915 1.35 3.035 1.435 ;
      RECT  1.85 1.435 3.035 1.555 ;
  END
END SEN_AO2BB2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO2BB2_DG_8
#      Description : "One 2-input NOR, and one 2-input AND, into a 2-input OR"
#      Equation    : X=(!A1&!A2)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO2BB2_DG_8
  CLASS CORE ;
  FOREIGN SEN_AO2BB2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.71 7.45 0.89 ;
      RECT  7.35 0.89 7.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  1.62 1.44 1.75 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  2.66 1.44 2.79 1.75 ;
      RECT  3.16 1.44 3.33 1.75 ;
      RECT  5.77 1.44 5.9 1.75 ;
      RECT  6.29 1.44 6.42 1.75 ;
      RECT  6.81 1.44 6.94 1.75 ;
      RECT  7.33 1.44 7.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  3.69 0.05 3.82 0.36 ;
      RECT  4.21 0.05 4.34 0.36 ;
      RECT  4.73 0.05 4.86 0.36 ;
      RECT  5.25 0.05 5.38 0.36 ;
      RECT  5.77 0.05 5.9 0.36 ;
      RECT  6.29 0.05 6.42 0.36 ;
      RECT  6.81 0.05 6.94 0.36 ;
      RECT  7.33 0.05 7.46 0.36 ;
      RECT  0.32 0.05 0.45 0.405 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.565 0.47 3.32 0.59 ;
      RECT  2.68 0.59 2.85 1.11 ;
      RECT  1.35 1.11 5.38 1.29 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.24 1.25 0.36 ;
      RECT  0.585 0.36 0.705 0.5 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.59 ;
      RECT  1.355 0.21 3.585 0.38 ;
      RECT  3.41 0.38 3.585 0.45 ;
      RECT  3.41 0.45 7.715 0.62 ;
      RECT  0.795 0.475 1.23 0.595 ;
      RECT  1.14 0.595 1.23 0.765 ;
      RECT  1.14 0.765 2.505 0.895 ;
      RECT  1.14 0.895 1.23 1.23 ;
      RECT  0.28 1.23 1.23 1.35 ;
      RECT  5.47 1.18 7.715 1.35 ;
      RECT  5.47 1.35 5.64 1.44 ;
      RECT  3.435 1.44 5.64 1.61 ;
  END
END SEN_AO2BB2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AO31_0P5
#      Description : "One 3-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO31_0P5
  CLASS CORE ;
  FOREIGN SEN_AO31_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.08 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0264 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.71 0.85 1.295 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0264 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0264 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0255 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.34 1.36 0.465 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.86 1.615 1.03 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.32 0.05 0.49 0.185 ;
      RECT  1.415 0.05 1.535 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.055 0.29 0.25 0.49 ;
      RECT  0.055 0.49 0.155 0.91 ;
      RECT  0.055 0.91 0.25 1.06 ;
      RECT  0.09 1.06 0.25 1.49 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.355 0.275 1.3 0.365 ;
      RECT  0.355 0.365 0.445 0.65 ;
      RECT  1.17 0.365 1.26 1.225 ;
      RECT  0.245 0.65 0.445 0.82 ;
      RECT  1.17 1.225 1.535 1.315 ;
      RECT  1.415 1.315 1.535 1.57 ;
      RECT  0.565 1.405 1.325 1.525 ;
  END
END SEN_AO31_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AO31_1
#      Description : "One 3-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO31_1
  CLASS CORE ;
  FOREIGN SEN_AO31_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.51 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.08 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.057 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.555 1.24 1.225 1.36 ;
      RECT  1.105 1.36 1.225 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  1.07 0.05 1.28 0.21 ;
      RECT  0.065 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.45 0.51 ;
      RECT  1.35 0.51 1.535 0.69 ;
      RECT  1.435 0.69 1.535 1.11 ;
      RECT  1.35 1.11 1.535 1.2 ;
      RECT  1.35 1.2 1.48 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.17 0.47 0.3 ;
      RECT  0.34 0.3 1.26 0.39 ;
      RECT  1.17 0.39 1.26 0.79 ;
      RECT  0.34 0.39 0.43 1.23 ;
      RECT  1.17 0.79 1.345 0.89 ;
      RECT  0.065 1.23 0.43 1.32 ;
      RECT  0.065 1.32 0.185 1.45 ;
      RECT  0.28 1.45 0.99 1.57 ;
  END
END SEN_AO31_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO31_2
#      Description : "One 3-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO31_2
  CLASS CORE ;
  FOREIGN SEN_AO31_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.114 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.285 1.445 0.465 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.85 1.565 1.02 1.75 ;
      RECT  1.46 1.565 1.63 1.75 ;
      RECT  2.52 1.015 2.63 1.75 ;
      RECT  3.02 1.41 3.15 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  1.355 0.05 1.475 0.375 ;
      RECT  3.025 0.05 3.145 0.39 ;
      RECT  1.875 0.05 1.995 0.56 ;
      RECT  2.52 0.05 2.625 0.565 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.31 2.875 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.23 1.265 0.34 ;
      RECT  0.055 0.34 0.175 0.43 ;
      RECT  2.1 0.45 2.43 0.555 ;
      RECT  2.34 0.555 2.43 0.755 ;
      RECT  2.34 0.755 2.65 0.925 ;
      RECT  2.34 0.925 2.43 1.18 ;
      RECT  0.26 0.475 0.65 0.59 ;
      RECT  0.56 0.59 0.65 1.02 ;
      RECT  0.56 1.02 0.86 1.115 ;
      RECT  0.77 1.115 0.86 1.18 ;
      RECT  0.77 1.18 2.43 1.28 ;
      RECT  0.81 0.465 1.76 0.585 ;
      RECT  0.055 1.23 0.68 1.35 ;
      RECT  0.575 1.35 0.68 1.37 ;
      RECT  0.055 1.35 0.17 1.59 ;
      RECT  0.575 1.37 1.915 1.47 ;
      RECT  1.795 1.47 1.915 1.5 ;
      RECT  1.795 1.5 2.43 1.59 ;
      RECT  2.315 1.415 2.43 1.5 ;
  END
END SEN_AO31_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO31_4
#      Description : "One 3-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO31_4
  CLASS CORE ;
  FOREIGN SEN_AO31_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.55 0.89 2.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  3.75 0.89 3.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.228 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.38 1.41 1.51 1.75 ;
      RECT  1.975 1.41 2.105 1.75 ;
      RECT  2.57 1.41 2.7 1.75 ;
      RECT  3.09 1.41 3.22 1.75 ;
      RECT  4.655 1.21 4.77 1.75 ;
      RECT  5.25 1.41 5.38 1.75 ;
      RECT  5.81 1.2 5.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  3.695 0.05 3.82 0.39 ;
      RECT  4.19 0.05 4.34 0.39 ;
      RECT  0.57 0.05 0.72 0.4 ;
      RECT  1.09 0.05 1.215 0.4 ;
      RECT  5.27 0.05 5.41 0.405 ;
      RECT  0.05 0.05 0.19 0.59 ;
      RECT  4.72 0.05 4.85 0.59 ;
      RECT  5.81 0.05 5.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.51 5.65 0.69 ;
      RECT  5.55 0.69 5.65 1.11 ;
      RECT  4.91 1.11 5.65 1.29 ;
    END
    ANTENNADIFFAREA 0.47 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.325 0.25 3.585 0.35 ;
      RECT  0.325 0.37 0.445 0.49 ;
      RECT  0.325 0.49 2.31 0.59 ;
      RECT  3.945 0.33 4.065 0.49 ;
      RECT  2.6 0.49 4.585 0.59 ;
      RECT  4.465 0.33 4.585 0.49 ;
      RECT  4.355 0.59 4.445 0.8 ;
      RECT  4.355 0.8 5.44 0.89 ;
      RECT  4.355 0.89 4.445 1.21 ;
      RECT  3.57 1.21 4.445 1.31 ;
      RECT  0.065 1.21 3.475 1.31 ;
      RECT  0.065 1.31 0.185 1.43 ;
      RECT  3.355 1.31 3.475 1.45 ;
      RECT  3.355 1.45 4.545 1.55 ;
  END
END SEN_AO31_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO31_8
#      Description : "One 3-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO31_8
  CLASS CORE ;
  FOREIGN SEN_AO31_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 6.05 0.915 ;
      RECT  5.95 0.915 6.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5064 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.65 0.92 ;
      RECT  2.75 0.92 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5064 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.915 ;
      RECT  0.75 0.915 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5064 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.71 8.05 0.89 ;
      RECT  7.95 0.89 8.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4566 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.445 0.45 1.75 ;
      RECT  0.0 1.75 11.0 1.85 ;
      RECT  0.84 1.445 0.97 1.75 ;
      RECT  1.36 1.445 1.49 1.75 ;
      RECT  1.88 1.445 2.01 1.75 ;
      RECT  2.4 1.445 2.53 1.75 ;
      RECT  2.92 1.445 3.05 1.75 ;
      RECT  3.44 1.445 3.57 1.75 ;
      RECT  3.96 1.445 4.09 1.75 ;
      RECT  4.48 1.445 4.61 1.75 ;
      RECT  5.0 1.445 5.13 1.75 ;
      RECT  5.52 1.445 5.65 1.75 ;
      RECT  6.04 1.445 6.17 1.75 ;
      RECT  8.635 1.21 8.755 1.75 ;
      RECT  9.15 1.41 9.28 1.75 ;
      RECT  9.67 1.41 9.8 1.75 ;
      RECT  10.19 1.41 10.32 1.75 ;
      RECT  10.73 1.21 10.85 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      RECT  6.905 0.05 7.075 0.34 ;
      RECT  7.485 0.05 7.655 0.34 ;
      RECT  8.005 0.05 8.175 0.34 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  0.84 0.05 0.97 0.36 ;
      RECT  1.36 0.05 1.49 0.36 ;
      RECT  1.88 0.05 2.01 0.36 ;
      RECT  9.065 0.05 9.195 0.36 ;
      RECT  9.585 0.05 9.715 0.36 ;
      RECT  10.105 0.05 10.235 0.36 ;
      RECT  8.55 0.05 8.67 0.59 ;
      RECT  10.66 0.05 10.78 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.785 0.455 10.515 0.585 ;
      RECT  10.08 0.585 10.25 1.11 ;
      RECT  8.91 1.11 10.585 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.35 0.17 6.45 0.34 ;
      RECT  6.565 0.33 6.685 0.43 ;
      RECT  4.485 0.43 8.425 0.6 ;
      RECT  8.255 0.6 8.425 0.755 ;
      RECT  8.255 0.755 9.94 0.925 ;
      RECT  8.255 0.925 8.425 1.18 ;
      RECT  6.56 1.18 8.425 1.35 ;
      RECT  0.065 0.37 0.185 0.45 ;
      RECT  0.065 0.45 4.37 0.59 ;
      RECT  0.065 1.185 6.425 1.355 ;
      RECT  6.27 1.355 6.425 1.445 ;
      RECT  6.27 1.445 8.53 1.615 ;
  END
END SEN_AO31_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AO32_0P5
#      Description : "One 3-input AND one 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO32_0P5
  CLASS CORE ;
  FOREIGN SEN_AO32_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.95 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.69 1.45 1.175 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0243 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.465 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.89 1.42 1.02 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.44 1.41 1.57 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.08 0.05 0.21 0.39 ;
      RECT  1.44 0.05 1.57 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.21 1.85 1.54 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.37 0.23 1.275 0.35 ;
      RECT  1.185 0.35 1.275 0.495 ;
      RECT  0.37 0.35 0.46 1.415 ;
      RECT  1.185 0.495 1.63 0.585 ;
      RECT  1.54 0.585 1.63 0.88 ;
      RECT  0.625 1.24 1.275 1.33 ;
      RECT  0.625 1.33 0.745 1.525 ;
      RECT  1.155 1.33 1.275 1.61 ;
      RECT  0.085 1.41 0.205 1.525 ;
      RECT  0.085 1.525 0.745 1.62 ;
  END
END SEN_AO32_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AO32_1
#      Description : "One 3-input AND one 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO32_1
  CLASS CORE ;
  FOREIGN SEN_AO32_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.5 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.5 1.05 0.71 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.24 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.88 1.57 1.05 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.5 1.39 1.63 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.45 0.05 1.63 0.21 ;
      RECT  0.07 0.05 0.21 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.3 1.91 0.69 ;
      RECT  1.82 0.69 1.91 1.1 ;
      RECT  1.75 1.1 1.91 1.5 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.56 0.3 1.64 0.39 ;
      RECT  1.55 0.39 1.64 0.78 ;
      RECT  1.55 0.78 1.725 0.9 ;
      RECT  1.55 0.9 1.64 1.21 ;
      RECT  0.34 1.21 1.64 1.3 ;
      RECT  0.34 1.3 0.445 1.43 ;
      RECT  0.585 1.39 1.345 1.48 ;
      RECT  0.585 1.48 0.705 1.54 ;
      RECT  1.225 1.48 1.345 1.61 ;
      RECT  0.065 1.41 0.185 1.54 ;
      RECT  0.065 1.54 0.705 1.64 ;
  END
END SEN_AO32_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO32_2
#      Description : "One 3-input AND one 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO32_2
  CLASS CORE ;
  FOREIGN SEN_AO32_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.7 2.45 0.9 ;
      RECT  2.15 0.9 2.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.84 0.71 3.05 0.9 ;
      RECT  2.95 0.9 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.7 3.65 0.9 ;
      RECT  3.55 0.9 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.685 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  2.135 1.405 2.255 1.75 ;
      RECT  2.585 1.41 2.705 1.75 ;
      RECT  3.105 1.41 3.225 1.75 ;
      RECT  3.625 1.41 3.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.065 0.05 0.185 0.39 ;
      RECT  1.105 0.05 1.225 0.39 ;
      RECT  3.365 0.05 3.485 0.39 ;
      RECT  0.585 0.05 0.705 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.335 0.31 0.45 0.51 ;
      RECT  0.15 0.51 0.45 0.69 ;
      RECT  0.15 0.69 0.25 1.0 ;
      RECT  0.15 1.0 0.45 1.09 ;
      RECT  0.335 1.09 0.45 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.135 0.14 2.965 0.23 ;
      RECT  2.135 0.23 2.255 0.38 ;
      RECT  2.845 0.23 2.965 0.385 ;
      RECT  2.37 0.32 2.54 0.415 ;
      RECT  2.37 0.415 2.46 0.505 ;
      RECT  1.355 0.17 1.995 0.28 ;
      RECT  1.355 0.28 1.475 0.39 ;
      RECT  1.875 0.28 1.995 0.505 ;
      RECT  1.875 0.505 2.46 0.595 ;
      RECT  1.875 0.595 1.995 1.0 ;
      RECT  1.615 1.0 1.995 1.105 ;
      RECT  1.615 1.105 1.735 1.21 ;
      RECT  0.34 0.79 0.65 0.89 ;
      RECT  0.56 0.89 0.65 1.21 ;
      RECT  0.56 1.21 1.735 1.32 ;
      RECT  3.62 0.19 3.75 0.495 ;
      RECT  2.585 0.495 3.75 0.6 ;
      RECT  2.585 0.6 2.705 0.71 ;
      RECT  0.845 0.37 0.965 0.5 ;
      RECT  0.845 0.5 1.735 0.59 ;
      RECT  1.615 0.37 1.735 0.5 ;
      RECT  1.875 1.195 3.54 1.315 ;
      RECT  1.875 1.315 1.995 1.44 ;
      RECT  0.81 1.44 1.995 1.56 ;
  END
END SEN_AO32_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO32_4
#      Description : "One 3-input AND one 2-input AND into 2-input OR"
#      Equation    : X=(A1&A2&A3)|(B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO32_4
  CLASS CORE ;
  FOREIGN SEN_AO32_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.45 0.9 ;
      RECT  3.95 0.9 4.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.45 0.9 ;
      RECT  4.95 0.9 5.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.71 6.85 0.9 ;
      RECT  6.35 0.9 6.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.9 ;
      RECT  2.55 0.9 2.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.9 ;
      RECT  1.55 0.9 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  0.59 1.41 0.72 1.75 ;
      RECT  1.115 1.21 1.225 1.75 ;
      RECT  3.7 1.41 3.83 1.75 ;
      RECT  4.225 1.41 4.355 1.75 ;
      RECT  4.745 1.41 4.875 1.75 ;
      RECT  5.265 1.41 5.395 1.75 ;
      RECT  5.815 1.41 5.945 1.75 ;
      RECT  6.39 1.41 6.52 1.75 ;
      RECT  6.96 1.21 7.08 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  5.97 0.05 6.1 0.38 ;
      RECT  0.59 0.05 0.72 0.39 ;
      RECT  1.1 0.05 1.255 0.39 ;
      RECT  1.6 0.05 1.73 0.39 ;
      RECT  2.12 0.05 2.25 0.39 ;
      RECT  6.49 0.05 6.62 0.39 ;
      RECT  0.075 0.05 0.195 0.59 ;
      RECT  7.015 0.05 7.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.51 1.05 0.69 ;
      RECT  0.34 0.69 0.46 1.11 ;
      RECT  0.34 1.11 0.99 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.425 0.19 3.545 0.3 ;
      RECT  2.385 0.3 3.545 0.4 ;
      RECT  2.385 0.4 2.49 0.49 ;
      RECT  1.29 0.49 2.49 0.59 ;
      RECT  3.655 0.19 3.775 0.3 ;
      RECT  3.655 0.3 5.865 0.4 ;
      RECT  5.745 0.19 5.865 0.3 ;
      RECT  6.755 0.37 6.875 0.49 ;
      RECT  4.9 0.49 6.875 0.59 ;
      RECT  2.6 0.49 4.61 0.59 ;
      RECT  3.175 0.59 3.31 1.21 ;
      RECT  0.57 0.795 1.445 0.885 ;
      RECT  1.355 0.885 1.445 1.21 ;
      RECT  1.355 1.21 3.31 1.31 ;
      RECT  3.445 1.21 6.85 1.31 ;
      RECT  3.445 1.31 3.565 1.42 ;
      RECT  1.335 1.42 3.565 1.52 ;
  END
END SEN_AO32_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AO33_1
#      Description : "Two 3-input ANDs into a 2-input OR"
#      Equation    : X=(A1&A2&A3)|(B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO33_1
  CLASS CORE ;
  FOREIGN SEN_AO33_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.705 0.665 0.85 0.835 ;
      RECT  0.75 0.835 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0396 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0396 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0396 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0396 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.745 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0396 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.005 ;
      RECT  1.55 1.005 1.69 1.215 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0396 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.48 0.5 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.85 1.48 1.02 1.75 ;
      RECT  1.395 1.485 1.565 1.75 ;
      RECT  1.915 1.485 2.085 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.43 0.05 1.605 0.32 ;
      RECT  0.085 0.05 0.225 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.92 0.215 1.27 0.335 ;
      RECT  1.15 0.335 1.27 1.29 ;
    END
    ANTENNADIFFAREA 0.19 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.2 0.2 2.32 0.3 ;
      RECT  1.695 0.3 2.32 0.42 ;
      RECT  1.695 0.42 1.785 0.435 ;
      RECT  1.37 0.435 1.785 0.53 ;
      RECT  1.37 0.53 1.46 1.305 ;
      RECT  1.37 1.305 2.32 1.395 ;
      RECT  1.68 1.395 1.8 1.54 ;
      RECT  2.2 1.395 2.32 1.54 ;
      RECT  0.72 0.455 1.06 0.575 ;
      RECT  0.96 0.575 1.06 1.3 ;
      RECT  0.095 1.3 1.06 1.39 ;
      RECT  0.095 1.39 0.215 1.54 ;
      RECT  0.615 1.39 0.735 1.54 ;
  END
END SEN_AO33_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AO33_2
#      Description : "Two 3-input ANDs into a 2-input OR"
#      Equation    : X=(A1&A2&A3)|(B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO33_2
  CLASS CORE ;
  FOREIGN SEN_AO33_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.25 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0744 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 3.65 0.91 ;
      RECT  3.55 0.91 3.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0744 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0744 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.695 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0744 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.75 0.91 1.05 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0744 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0744 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.05 1.41 0.18 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.81 1.495 0.98 1.75 ;
      RECT  1.555 1.495 1.725 1.75 ;
      RECT  2.235 1.41 2.365 1.75 ;
      RECT  2.855 1.495 3.025 1.75 ;
      RECT  3.62 1.495 3.79 1.75 ;
      RECT  4.42 1.41 4.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.31 0.05 0.48 0.32 ;
      RECT  4.125 0.05 4.255 0.345 ;
      RECT  1.975 0.05 2.105 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.475 0.575 2.65 0.665 ;
      RECT  2.55 0.665 2.65 1.11 ;
      RECT  1.95 1.11 2.65 1.29 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.96 0.19 3.68 0.305 ;
      RECT  2.96 0.305 3.065 0.365 ;
      RECT  0.93 0.225 1.705 0.335 ;
      RECT  0.075 0.31 0.195 0.415 ;
      RECT  0.075 0.415 0.79 0.535 ;
      RECT  4.39 0.31 4.51 0.435 ;
      RECT  3.795 0.435 4.51 0.54 ;
      RECT  2.24 0.395 2.875 0.485 ;
      RECT  2.24 0.485 2.36 0.495 ;
      RECT  2.76 0.485 2.875 0.645 ;
      RECT  1.695 0.495 2.36 0.615 ;
      RECT  3.155 0.42 3.445 0.54 ;
      RECT  3.355 0.54 3.445 1.3 ;
      RECT  2.74 0.755 2.835 1.3 ;
      RECT  2.74 1.3 4.145 1.405 ;
      RECT  3.325 1.405 3.445 1.55 ;
      RECT  4.025 1.405 4.145 1.55 ;
      RECT  1.755 0.785 2.16 0.895 ;
      RECT  1.755 0.895 1.86 1.3 ;
      RECT  1.155 0.425 1.45 0.54 ;
      RECT  1.155 0.54 1.245 1.3 ;
      RECT  0.455 1.3 1.86 1.405 ;
      RECT  0.455 1.405 0.575 1.55 ;
      RECT  1.19 1.405 1.31 1.55 ;
  END
END SEN_AO33_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AO33_4
#      Description : "Two 3-input ANDs into a 2-input OR"
#      Equation    : X=(A1&A2&A3)|(B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AO33_4
  CLASS CORE ;
  FOREIGN SEN_AO33_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1419 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.945 0.71 6.45 0.89 ;
      RECT  6.35 0.89 6.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1419 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.71 7.05 0.89 ;
      RECT  6.95 0.89 7.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1419 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1419 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1419 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1419 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.24 1.21 0.36 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  0.82 1.455 0.99 1.75 ;
      RECT  1.34 1.45 1.51 1.75 ;
      RECT  1.6 1.45 1.77 1.75 ;
      RECT  2.155 1.455 2.325 1.75 ;
      RECT  2.59 1.21 2.71 1.75 ;
      RECT  3.105 1.41 3.235 1.75 ;
      RECT  3.625 1.41 3.755 1.75 ;
      RECT  4.145 1.41 4.275 1.75 ;
      RECT  4.67 1.21 4.79 1.75 ;
      RECT  4.98 1.46 5.155 1.75 ;
      RECT  5.535 1.46 5.705 1.75 ;
      RECT  5.87 1.46 6.04 1.75 ;
      RECT  6.39 1.465 6.56 1.75 ;
      RECT  7.04 1.21 7.16 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  2.845 0.05 2.975 0.35 ;
      RECT  3.365 0.05 3.48 0.35 ;
      RECT  6.67 0.05 6.8 0.35 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  7.215 0.05 7.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.44 4.58 0.565 ;
      RECT  3.75 0.565 3.85 1.11 ;
      RECT  2.85 1.11 4.53 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.57 0.24 4.84 0.35 ;
      RECT  3.57 0.35 3.66 0.44 ;
      RECT  2.6 0.17 2.725 0.44 ;
      RECT  2.6 0.44 3.66 0.56 ;
      RECT  5.06 0.24 6.33 0.35 ;
      RECT  1.055 0.24 2.325 0.36 ;
      RECT  0.275 0.45 1.535 0.56 ;
      RECT  1.83 0.45 2.51 0.56 ;
      RECT  2.395 0.56 2.51 0.78 ;
      RECT  2.395 0.78 3.425 0.895 ;
      RECT  2.395 0.895 2.5 1.24 ;
      RECT  0.535 1.24 2.5 1.36 ;
      RECT  4.855 0.44 5.545 0.56 ;
      RECT  4.855 0.56 4.97 0.785 ;
      RECT  3.99 0.785 4.97 0.895 ;
      RECT  4.88 0.895 4.97 1.25 ;
      RECT  4.88 1.25 6.845 1.37 ;
      RECT  5.84 0.44 7.105 0.57 ;
  END
END SEN_AO33_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOA211_DG_1
#      Description : "One 2-input AND into 2-input OR into 2-input AND"
#      Equation    : X=((A1&A2)|B)&C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOA211_DG_1
  CLASS CORE ;
  FOREIGN SEN_AOA211_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.63 0.85 0.995 ;
      RECT  0.655 0.995 0.85 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.635 1.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.13 1.44 1.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.555 0.05 0.685 0.35 ;
      RECT  1.35 0.05 1.48 0.5 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.615 0.3 1.735 0.6 ;
      RECT  1.55 0.6 1.735 0.69 ;
      RECT  1.55 0.69 1.65 1.3 ;
    END
    ANTENNADIFFAREA 0.185 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.44 0.39 ;
      RECT  0.35 0.39 0.44 0.44 ;
      RECT  0.35 0.44 0.965 0.53 ;
      RECT  0.845 0.25 0.965 0.44 ;
      RECT  1.12 0.25 1.24 0.42 ;
      RECT  1.15 0.42 1.24 0.785 ;
      RECT  1.15 0.785 1.45 0.895 ;
      RECT  1.15 0.895 1.24 1.26 ;
      RECT  0.845 1.26 1.24 1.35 ;
      RECT  0.845 1.35 0.965 1.59 ;
      RECT  0.065 1.26 0.705 1.35 ;
      RECT  0.065 1.35 0.185 1.59 ;
      RECT  0.585 1.35 0.705 1.59 ;
  END
END SEN_AOA211_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOA211_DG_2
#      Description : "One 2-input AND into 2-input OR into 2-input AND"
#      Equation    : X=((A1&A2)|B)&C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOA211_DG_2
  CLASS CORE ;
  FOREIGN SEN_AOA211_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.63 0.85 0.995 ;
      RECT  0.64 0.995 0.85 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.635 1.05 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.44 0.44 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.09 1.44 1.22 1.75 ;
      RECT  1.66 1.41 1.79 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.545 0.05 0.675 0.35 ;
      RECT  1.82 0.05 1.945 0.39 ;
      RECT  1.32 0.05 1.43 0.68 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.67 1.11 ;
      RECT  1.33 1.11 1.67 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.17 0.175 0.3 ;
      RECT  0.055 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 0.44 ;
      RECT  0.34 0.44 0.955 0.53 ;
      RECT  0.835 0.21 0.955 0.44 ;
      RECT  1.11 0.195 1.23 0.365 ;
      RECT  1.14 0.365 1.23 0.785 ;
      RECT  1.14 0.785 1.45 0.895 ;
      RECT  1.14 0.895 1.23 1.26 ;
      RECT  0.835 1.26 1.23 1.35 ;
      RECT  0.835 1.35 0.955 1.53 ;
      RECT  0.055 1.26 0.695 1.35 ;
      RECT  0.575 1.35 0.695 1.53 ;
      RECT  0.055 1.35 0.175 1.61 ;
  END
END SEN_AOA211_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOA211_DG_4
#      Description : "One 2-input AND into 2-input OR into 2-input AND"
#      Equation    : X=((A1&A2)|B)&C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOA211_DG_4
  CLASS CORE ;
  FOREIGN SEN_AOA211_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.6 0.45 0.755 ;
      RECT  0.35 0.755 0.525 0.925 ;
      RECT  0.35 0.925 0.45 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.6 0.85 0.755 ;
      RECT  0.69 0.755 0.85 0.925 ;
      RECT  0.75 0.925 0.85 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.6 1.05 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.44 0.44 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.09 1.44 1.22 1.75 ;
      RECT  1.61 1.41 1.74 1.75 ;
      RECT  2.16 1.21 2.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.525 0.05 0.695 0.31 ;
      RECT  1.8 0.05 1.97 0.345 ;
      RECT  2.36 0.05 2.48 0.59 ;
      RECT  1.32 0.05 1.425 0.67 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.3 1.685 0.475 ;
      RECT  1.55 0.475 2.25 0.565 ;
      RECT  2.085 0.3 2.25 0.475 ;
      RECT  1.95 0.565 2.05 1.11 ;
      RECT  1.35 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.17 0.175 0.3 ;
      RECT  0.055 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 0.4 ;
      RECT  0.34 0.4 0.955 0.49 ;
      RECT  0.835 0.27 0.955 0.4 ;
      RECT  1.11 0.195 1.23 0.365 ;
      RECT  1.14 0.365 1.23 0.785 ;
      RECT  1.14 0.785 1.84 0.895 ;
      RECT  1.14 0.895 1.23 1.26 ;
      RECT  0.835 1.26 1.23 1.35 ;
      RECT  0.835 1.35 0.955 1.5 ;
      RECT  0.055 1.26 0.695 1.35 ;
      RECT  0.575 1.35 0.695 1.5 ;
      RECT  0.055 1.35 0.175 1.61 ;
  END
END SEN_AOA211_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOA211_DG_8
#      Description : "One 2-input AND into 2-input OR into 2-input AND"
#      Equation    : X=((A1&A2)|B)&C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOA211_DG_8
  CLASS CORE ;
  FOREIGN SEN_AOA211_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.47 2.45 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.455 0.445 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.845 1.455 0.965 1.75 ;
      RECT  2.07 1.44 2.19 1.75 ;
      RECT  2.535 1.425 2.655 1.75 ;
      RECT  3.055 1.425 3.175 1.75 ;
      RECT  3.575 1.425 3.695 1.75 ;
      RECT  4.095 1.425 4.215 1.75 ;
      RECT  4.615 1.24 4.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  1.55 0.05 1.67 0.36 ;
      RECT  3.055 0.05 3.175 0.365 ;
      RECT  3.575 0.05 3.695 0.365 ;
      RECT  4.095 0.05 4.215 0.365 ;
      RECT  4.615 0.05 4.735 0.56 ;
      RECT  2.54 0.05 2.655 0.655 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 4.5 0.69 ;
      RECT  4.08 0.69 4.25 1.11 ;
      RECT  2.75 1.11 4.49 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.81 0.18 2.45 0.27 ;
      RECT  2.33 0.27 2.45 0.36 ;
      RECT  1.81 0.27 1.93 0.5 ;
      RECT  0.82 0.5 1.93 0.62 ;
      RECT  0.585 0.21 1.25 0.335 ;
      RECT  0.585 0.335 0.69 0.45 ;
      RECT  0.065 0.32 0.185 0.45 ;
      RECT  0.065 0.45 0.69 0.54 ;
      RECT  2.56 0.78 3.895 0.9 ;
      RECT  2.56 0.9 2.65 1.05 ;
      RECT  2.07 0.36 2.19 1.05 ;
      RECT  2.07 1.05 2.65 1.17 ;
      RECT  2.07 1.17 2.185 1.21 ;
      RECT  1.305 1.01 1.41 1.21 ;
      RECT  1.305 1.21 2.185 1.33 ;
      RECT  0.065 1.245 1.215 1.365 ;
      RECT  1.105 1.365 1.215 1.455 ;
      RECT  0.065 1.365 0.185 1.47 ;
      RECT  1.105 1.455 1.72 1.575 ;
  END
END SEN_AOA211_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_1
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_1
  CLASS CORE ;
  FOREIGN SEN_AOAI211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.345 0.71 0.65 0.89 ;
      RECT  0.345 0.89 0.45 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.805 1.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.305 1.435 0.475 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.2 1.41 1.355 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.595 0.05 0.805 0.24 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.335 0.485 ;
      RECT  1.15 0.485 1.255 0.51 ;
      RECT  0.95 0.51 1.255 0.69 ;
      RECT  0.95 0.69 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.205 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.19 0.185 0.33 ;
      RECT  0.065 0.33 1.05 0.42 ;
      RECT  0.94 0.2 1.05 0.33 ;
      RECT  0.065 1.225 0.81 1.325 ;
      RECT  0.065 1.325 0.185 1.45 ;
  END
END SEN_AOAI211_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_2
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_2
  CLASS CORE ;
  FOREIGN SEN_AOAI211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.085 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.485 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.685 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.8 ;
      RECT  2.185 0.8 2.45 0.91 ;
      RECT  2.35 0.91 2.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.435 0.47 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.82 1.435 0.99 1.75 ;
      RECT  2.11 1.435 2.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.59 0.05 1.76 0.305 ;
      RECT  0.28 0.05 0.49 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.145 0.415 2.25 0.575 ;
      RECT  1.945 0.575 2.25 0.69 ;
      RECT  1.945 0.69 2.055 1.21 ;
      RECT  1.88 1.21 2.535 1.3 ;
      RECT  1.88 1.3 1.99 1.43 ;
      RECT  2.415 1.3 2.535 1.43 ;
      RECT  1.3 1.43 1.99 1.55 ;
    END
    ANTENNADIFFAREA 0.414 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.875 0.17 2.525 0.26 ;
      RECT  2.405 0.26 2.525 0.39 ;
      RECT  1.875 0.26 1.995 0.395 ;
      RECT  1.35 0.395 1.995 0.485 ;
      RECT  1.35 0.485 1.48 0.49 ;
      RECT  0.82 0.49 1.48 0.59 ;
      RECT  0.585 0.24 1.25 0.345 ;
      RECT  0.585 0.345 0.705 0.5 ;
      RECT  0.06 0.37 0.19 0.5 ;
      RECT  0.06 0.5 0.705 0.59 ;
      RECT  0.065 1.185 1.77 1.285 ;
      RECT  0.065 1.285 0.185 1.42 ;
  END
END SEN_AOAI211_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_3
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_3
  CLASS CORE ;
  FOREIGN SEN_AOAI211_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.215 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.225 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.08 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1908 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.485 0.47 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.82 1.475 0.99 1.75 ;
      RECT  1.34 1.485 1.51 1.75 ;
      RECT  2.83 1.465 3.0 1.75 ;
      RECT  3.415 1.42 3.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  2.35 0.05 2.52 0.32 ;
      RECT  1.83 0.05 2.0 0.335 ;
      RECT  0.56 0.05 0.73 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.9 0.42 3.05 0.5 ;
      RECT  2.9 0.5 3.535 0.59 ;
      RECT  3.415 0.41 3.535 0.5 ;
      RECT  2.95 0.59 3.05 1.11 ;
      RECT  2.545 1.11 3.26 1.29 ;
      RECT  2.545 1.29 2.65 1.48 ;
      RECT  1.93 1.48 2.65 1.6 ;
    END
    ANTENNADIFFAREA 0.548 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.63 0.21 3.3 0.32 ;
      RECT  2.63 0.32 2.76 0.445 ;
      RECT  1.08 0.23 1.74 0.34 ;
      RECT  1.63 0.34 1.74 0.445 ;
      RECT  1.63 0.445 2.76 0.55 ;
      RECT  0.3 0.48 1.51 0.59 ;
      RECT  0.065 1.245 2.435 1.36 ;
      RECT  0.065 1.36 0.185 1.48 ;
  END
END SEN_AOAI211_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_4
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_4
  CLASS CORE ;
  FOREIGN SEN_AOAI211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.45 0.435 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.835 1.45 0.955 1.75 ;
      RECT  1.355 1.45 1.475 1.75 ;
      RECT  1.875 1.45 1.995 1.75 ;
      RECT  3.63 1.425 3.755 1.75 ;
      RECT  4.14 1.43 4.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.315 0.05 0.435 0.385 ;
      RECT  0.835 0.05 0.955 0.385 ;
      RECT  2.58 0.05 2.7 0.385 ;
      RECT  3.1 0.05 3.22 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.615 0.47 4.295 0.58 ;
      RECT  3.615 0.58 3.85 0.665 ;
      RECT  3.75 0.665 3.85 1.11 ;
      RECT  3.42 1.11 4.25 1.22 ;
      RECT  3.42 1.22 4.52 1.31 ;
      RECT  4.4 1.31 4.52 1.44 ;
      RECT  3.42 1.31 3.54 1.475 ;
      RECT  2.37 1.475 3.54 1.6 ;
    END
    ANTENNADIFFAREA 0.714 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.34 0.17 4.52 0.32 ;
      RECT  4.395 0.32 4.52 0.39 ;
      RECT  3.34 0.32 3.485 0.475 ;
      RECT  1.33 0.23 2.465 0.35 ;
      RECT  2.35 0.35 2.465 0.475 ;
      RECT  2.35 0.475 3.485 0.59 ;
      RECT  0.05 0.19 0.18 0.475 ;
      RECT  0.05 0.475 2.24 0.59 ;
      RECT  2.15 0.59 2.24 0.68 ;
      RECT  3.175 1.09 3.295 1.2 ;
      RECT  0.05 1.2 3.295 1.315 ;
      RECT  0.05 1.315 0.18 1.61 ;
  END
END SEN_AOAI211_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_6
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_6
  CLASS CORE ;
  FOREIGN SEN_AOAI211_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.935 0.9 ;
      RECT  1.46 0.71 1.85 0.89 ;
      RECT  0.43 0.71 0.85 0.89 ;
      LAYER M2 ;
      RECT  0.435 0.75 2.73 0.85 ;
      LAYER V1 ;
      RECT  2.565 0.75 2.665 0.85 ;
      RECT  1.505 0.75 1.605 0.85 ;
      RECT  1.705 0.75 1.805 0.85 ;
      RECT  0.475 0.75 0.575 0.85 ;
      RECT  0.675 0.75 0.775 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.005 ;
      RECT  0.15 1.005 3.25 1.095 ;
      RECT  1.15 0.71 1.25 1.005 ;
      RECT  2.15 0.71 2.25 1.005 ;
      RECT  3.095 0.71 3.25 1.005 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 4.45 0.89 ;
      RECT  3.55 0.89 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.51 6.65 0.71 ;
      RECT  5.75 0.71 6.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3798 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  1.88 1.44 2.01 1.75 ;
      RECT  2.4 1.44 2.53 1.75 ;
      RECT  2.92 1.44 3.05 1.75 ;
      RECT  4.99 1.41 5.12 1.75 ;
      RECT  5.51 1.41 5.64 1.75 ;
      RECT  6.03 1.41 6.16 1.75 ;
      RECT  6.57 1.21 6.69 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  3.18 0.05 3.31 0.36 ;
      RECT  3.7 0.05 3.83 0.36 ;
      RECT  4.22 0.05 4.35 0.36 ;
      RECT  4.74 0.05 4.87 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.215 0.47 6.46 0.59 ;
      RECT  5.32 0.59 5.45 1.11 ;
      RECT  3.75 1.11 6.45 1.2 ;
      RECT  3.42 1.2 6.45 1.3 ;
    END
    ANTENNADIFFAREA 0.996 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.985 0.23 6.71 0.36 ;
      RECT  4.985 0.36 5.115 0.45 ;
      RECT  0.525 0.45 5.115 0.58 ;
      RECT  0.065 1.22 3.305 1.35 ;
      RECT  0.065 1.35 0.185 1.44 ;
      RECT  3.175 1.35 3.305 1.45 ;
      RECT  3.175 1.45 4.89 1.58 ;
  END
END SEN_AOAI211_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_8
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_8
  CLASS CORE ;
  FOREIGN SEN_AOAI211_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.43 0.71 3.975 0.89 ;
      RECT  2.55 0.71 2.85 0.9 ;
      RECT  1.55 0.71 1.875 0.9 ;
      RECT  0.55 0.71 0.85 0.89 ;
      LAYER M2 ;
      RECT  0.51 0.75 3.89 0.85 ;
      LAYER V1 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.25 1.0 ;
      RECT  3.15 1.0 3.605 1.005 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.45 1.005 ;
      RECT  0.15 1.005 4.25 1.095 ;
      RECT  1.15 0.71 1.25 1.005 ;
      RECT  2.15 0.71 2.25 1.005 ;
      RECT  4.135 0.71 4.25 1.005 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 5.65 0.89 ;
      RECT  4.55 0.89 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.48 0.71 8.65 0.9 ;
      RECT  8.55 0.9 8.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5064 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.455 0.45 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.84 1.455 0.97 1.75 ;
      RECT  1.36 1.455 1.49 1.75 ;
      RECT  1.88 1.455 2.01 1.75 ;
      RECT  2.4 1.455 2.53 1.75 ;
      RECT  2.92 1.455 3.05 1.75 ;
      RECT  3.44 1.455 3.57 1.75 ;
      RECT  3.96 1.455 4.085 1.75 ;
      RECT  6.53 1.41 6.66 1.75 ;
      RECT  7.05 1.41 7.18 1.75 ;
      RECT  7.57 1.41 7.7 1.75 ;
      RECT  8.09 1.41 8.22 1.75 ;
      RECT  8.62 1.41 8.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  3.18 0.05 3.31 0.36 ;
      RECT  4.22 0.05 4.35 0.36 ;
      RECT  4.74 0.05 4.87 0.36 ;
      RECT  5.26 0.05 5.39 0.36 ;
      RECT  5.78 0.05 5.91 0.36 ;
      RECT  6.3 0.05 6.425 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.775 0.45 8.53 0.585 ;
      RECT  6.775 0.585 7.32 0.595 ;
      RECT  7.15 0.595 7.32 1.11 ;
      RECT  4.75 1.11 8.45 1.19 ;
      RECT  4.46 1.19 8.45 1.2 ;
      RECT  4.46 1.2 8.545 1.3 ;
    END
    ANTENNADIFFAREA 1.332 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.515 0.19 8.74 0.36 ;
      RECT  6.515 0.36 6.685 0.45 ;
      RECT  0.585 0.45 6.685 0.62 ;
      RECT  0.065 1.195 4.345 1.365 ;
      RECT  4.175 1.365 4.345 1.44 ;
      RECT  4.175 1.44 6.44 1.61 ;
  END
END SEN_AOAI211_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_0P5
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_0P5
  CLASS CORE ;
  FOREIGN SEN_AOAI211_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.63 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.815 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.125 1.41 1.255 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.555 0.05 0.685 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.105 0.21 1.25 0.625 ;
      RECT  0.95 0.625 1.25 0.725 ;
      RECT  0.95 0.725 1.05 1.225 ;
      RECT  0.845 1.225 1.05 1.315 ;
      RECT  0.845 1.315 0.965 1.55 ;
    END
    ANTENNADIFFAREA 0.097 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.44 0.39 ;
      RECT  0.35 0.39 0.44 0.445 ;
      RECT  0.35 0.445 0.965 0.535 ;
      RECT  0.845 0.21 0.965 0.445 ;
      RECT  0.065 1.26 0.705 1.35 ;
      RECT  0.065 1.35 0.185 1.53 ;
      RECT  0.585 1.35 0.705 1.53 ;
  END
END SEN_AOAI211_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_0P75
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_0P75
  CLASS CORE ;
  FOREIGN SEN_AOAI211_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.63 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.815 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.12 1.42 1.25 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.555 0.05 0.685 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.105 0.31 1.25 0.625 ;
      RECT  0.95 0.625 1.25 0.725 ;
      RECT  0.95 0.725 1.05 1.26 ;
      RECT  0.845 1.26 1.05 1.35 ;
      RECT  0.845 1.35 0.965 1.48 ;
    END
    ANTENNADIFFAREA 0.145 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.44 0.39 ;
      RECT  0.35 0.39 0.44 0.435 ;
      RECT  0.35 0.435 0.965 0.525 ;
      RECT  0.845 0.3 0.965 0.435 ;
      RECT  0.065 1.26 0.705 1.35 ;
      RECT  0.065 1.35 0.185 1.48 ;
      RECT  0.585 1.35 0.705 1.48 ;
  END
END SEN_AOAI211_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_G_0P5
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_G_0P5
  CLASS CORE ;
  FOREIGN SEN_AOAI211_G_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.63 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.815 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.125 1.41 1.255 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.555 0.05 0.685 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.105 0.21 1.25 0.625 ;
      RECT  0.95 0.625 1.25 0.725 ;
      RECT  0.95 0.725 1.05 1.26 ;
      RECT  0.845 1.26 1.05 1.35 ;
      RECT  0.845 1.35 0.965 1.53 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.44 0.39 ;
      RECT  0.35 0.39 0.44 0.445 ;
      RECT  0.35 0.445 0.965 0.535 ;
      RECT  0.845 0.21 0.965 0.445 ;
      RECT  0.065 1.26 0.705 1.35 ;
      RECT  0.065 1.35 0.185 1.53 ;
      RECT  0.585 1.35 0.705 1.53 ;
  END
END SEN_AOAI211_G_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_G_0P75
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_G_0P75
  CLASS CORE ;
  FOREIGN SEN_AOAI211_G_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.63 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.815 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.135 1.41 1.265 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.555 0.05 0.685 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.105 0.31 1.25 0.625 ;
      RECT  0.95 0.625 1.25 0.725 ;
      RECT  0.95 0.725 1.05 1.26 ;
      RECT  0.845 1.26 1.05 1.35 ;
      RECT  0.845 1.35 0.965 1.48 ;
    END
    ANTENNADIFFAREA 0.147 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.44 0.39 ;
      RECT  0.35 0.39 0.44 0.435 ;
      RECT  0.35 0.435 0.965 0.525 ;
      RECT  0.845 0.3 0.965 0.435 ;
      RECT  0.065 1.26 0.705 1.35 ;
      RECT  0.065 1.35 0.185 1.48 ;
      RECT  0.585 1.35 0.705 1.48 ;
  END
END SEN_AOAI211_G_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_G_1
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_G_1
  CLASS CORE ;
  FOREIGN SEN_AOAI211_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.63 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.8 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.39 0.45 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.125 1.41 1.255 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.555 0.05 0.685 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.105 0.31 1.25 0.62 ;
      RECT  0.95 0.62 1.25 0.71 ;
      RECT  0.95 0.71 1.05 1.21 ;
      RECT  0.845 1.21 1.05 1.3 ;
      RECT  0.845 1.3 0.965 1.43 ;
    END
    ANTENNADIFFAREA 0.197 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.17 0.185 0.3 ;
      RECT  0.065 0.3 0.44 0.39 ;
      RECT  0.35 0.39 0.44 0.44 ;
      RECT  0.35 0.44 0.965 0.53 ;
      RECT  0.845 0.31 0.965 0.44 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.585 1.3 0.705 1.43 ;
  END
END SEN_AOAI211_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_G_2
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_G_2
  CLASS CORE ;
  FOREIGN SEN_AOAI211_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.85 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 1.02 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.455 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.84 1.455 0.97 1.75 ;
      RECT  2.13 1.41 2.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  1.61 0.05 1.74 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.36 2.25 1.11 ;
      RECT  1.35 1.11 2.515 1.29 ;
    END
    ANTENNADIFFAREA 0.408 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.875 0.18 2.515 0.27 ;
      RECT  2.395 0.27 2.515 0.41 ;
      RECT  1.875 0.27 1.995 0.475 ;
      RECT  0.82 0.475 1.995 0.595 ;
      RECT  0.585 0.21 1.28 0.335 ;
      RECT  0.585 0.335 0.705 0.45 ;
      RECT  0.065 0.32 0.185 0.45 ;
      RECT  0.065 0.45 0.705 0.54 ;
      RECT  0.065 1.24 1.225 1.36 ;
      RECT  1.105 1.36 1.225 1.425 ;
      RECT  0.065 1.36 0.185 1.46 ;
      RECT  1.105 1.425 1.79 1.545 ;
  END
END SEN_AOAI211_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_G_3
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_G_3
  CLASS CORE ;
  FOREIGN SEN_AOAI211_G_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.9 ;
      RECT  1.35 0.9 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.9 ;
      RECT  0.55 0.9 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.45 0.9 ;
      RECT  1.75 0.9 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.45 0.925 ;
      RECT  3.35 0.925 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.18 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.575 1.44 0.7 1.75 ;
      RECT  1.09 1.44 1.22 1.75 ;
      RECT  1.61 1.44 1.74 1.75 ;
      RECT  2.9 1.41 3.03 1.75 ;
      RECT  3.425 1.41 3.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.57 0.05 0.7 0.36 ;
      RECT  1.86 0.05 1.99 0.36 ;
      RECT  2.38 0.05 2.51 0.36 ;
      RECT  0.055 0.05 0.18 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.425 0.19 3.545 0.45 ;
      RECT  2.905 0.45 3.545 0.54 ;
      RECT  2.905 0.54 3.05 0.62 ;
      RECT  2.95 0.62 3.05 1.11 ;
      RECT  2.125 1.11 3.05 1.205 ;
      RECT  2.125 1.205 3.335 1.3 ;
    END
    ANTENNADIFFAREA 0.52 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.645 0.215 3.335 0.335 ;
      RECT  2.645 0.335 2.765 0.45 ;
      RECT  1.04 0.24 1.735 0.36 ;
      RECT  1.615 0.36 1.735 0.45 ;
      RECT  1.615 0.45 2.765 0.57 ;
      RECT  0.26 0.475 1.525 0.595 ;
      RECT  0.265 1.23 1.985 1.35 ;
      RECT  1.865 1.35 1.985 1.44 ;
      RECT  1.865 1.44 2.56 1.56 ;
  END
END SEN_AOAI211_G_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOAI211_G_4
#      Description : "One 2-input AND into 2-input OR into 2-input NAND"
#      Equation    : X=!(((A1&A2)|B)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOAI211_G_4
  CLASS CORE ;
  FOREIGN SEN_AOAI211_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 3.05 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  1.88 1.44 2.01 1.75 ;
      RECT  3.625 1.395 3.755 1.75 ;
      RECT  4.145 1.395 4.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.59 0.05 2.715 0.36 ;
      RECT  3.105 0.05 3.235 0.36 ;
      RECT  0.32 0.05 0.45 0.375 ;
      RECT  0.84 0.05 0.97 0.375 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.58 0.475 4.32 0.595 ;
      RECT  3.75 0.595 3.85 1.11 ;
      RECT  2.405 1.11 3.85 1.205 ;
      RECT  2.405 1.205 4.53 1.295 ;
      RECT  4.41 1.295 4.53 1.425 ;
    END
    ANTENNADIFFAREA 0.724 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.37 0.2 4.53 0.32 ;
      RECT  4.41 0.32 4.53 0.43 ;
      RECT  3.37 0.32 3.49 0.475 ;
      RECT  1.315 0.215 2.5 0.335 ;
      RECT  2.41 0.335 2.5 0.475 ;
      RECT  2.41 0.475 3.49 0.595 ;
      RECT  0.065 0.375 0.185 0.475 ;
      RECT  0.065 0.475 2.32 0.595 ;
      RECT  0.065 1.23 2.265 1.35 ;
      RECT  0.065 1.35 0.185 1.45 ;
      RECT  2.145 1.35 2.265 1.465 ;
      RECT  2.145 1.465 3.355 1.585 ;
  END
END SEN_AOAI211_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_0P5
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI211_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.05 ;
      RECT  0.35 1.05 0.575 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.64 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.75 ;
      RECT  0.55 0.75 0.68 0.935 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.435 0.435 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.775 0.05 0.945 0.18 ;
      RECT  0.045 0.05 0.215 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.45 0.275 1.135 0.395 ;
      RECT  1.015 0.395 1.135 0.55 ;
      RECT  0.75 0.395 0.86 0.69 ;
      RECT  0.77 0.69 0.86 1.015 ;
      RECT  0.75 1.015 0.86 1.285 ;
      RECT  0.75 1.285 1.145 1.375 ;
      RECT  0.95 1.375 1.145 1.49 ;
    END
    ANTENNADIFFAREA 0.127 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.06 1.245 0.65 1.335 ;
      RECT  0.55 1.335 0.65 1.465 ;
      RECT  0.06 1.335 0.17 1.62 ;
      RECT  0.55 1.465 0.75 1.575 ;
  END
END SEN_AOI211_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_1
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_1
  CLASS CORE ;
  FOREIGN SEN_AOI211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.5 0.45 0.755 ;
      RECT  0.35 0.755 0.535 0.925 ;
      RECT  0.35 0.925 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.055 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.735 0.51 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.495 0.52 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.86 0.05 1.03 0.23 ;
      RECT  0.095 0.05 0.24 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.615 0.2 0.735 0.32 ;
      RECT  0.615 0.32 1.26 0.42 ;
      RECT  1.15 0.21 1.26 0.32 ;
      RECT  1.15 0.42 1.26 1.3 ;
    END
    ANTENNADIFFAREA 0.261 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.09 1.3 0.74 1.39 ;
      RECT  0.09 1.39 0.22 1.52 ;
      RECT  0.61 1.39 0.74 1.52 ;
  END
END SEN_AOI211_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_2
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_2
  CLASS CORE ;
  FOREIGN SEN_AOI211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.21 0.19 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.56 1.48 0.73 1.75 ;
      RECT  1.08 1.48 1.25 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.605 0.05 1.775 0.36 ;
      RECT  2.125 0.05 2.295 0.36 ;
      RECT  0.28 0.05 0.49 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.37 2.53 0.49 ;
      RECT  0.82 0.49 2.53 0.59 ;
      RECT  1.95 0.59 2.05 1.11 ;
      RECT  1.95 1.11 2.26 1.29 ;
    END
    ANTENNADIFFAREA 0.45 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.58 0.235 1.28 0.35 ;
      RECT  0.58 0.35 0.705 0.5 ;
      RECT  0.06 0.37 0.19 0.5 ;
      RECT  0.06 0.5 0.705 0.59 ;
      RECT  0.28 1.25 1.8 1.355 ;
      RECT  2.41 1.34 2.53 1.46 ;
      RECT  1.345 1.46 2.53 1.56 ;
  END
END SEN_AOI211_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_3
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_3
  CLASS CORE ;
  FOREIGN SEN_AOI211_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.189 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.189 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.82 1.48 0.99 1.75 ;
      RECT  1.34 1.48 1.51 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.54 0.05 0.75 0.34 ;
      RECT  1.86 0.05 2.03 0.365 ;
      RECT  2.38 0.05 2.55 0.365 ;
      RECT  2.9 0.05 3.07 0.365 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.185 0.355 3.305 0.47 ;
      RECT  1.08 0.47 3.305 0.575 ;
      RECT  2.55 0.575 2.65 1.11 ;
      RECT  2.55 1.11 3.05 1.265 ;
      RECT  2.55 1.265 3.29 1.29 ;
      RECT  2.95 1.29 3.29 1.355 ;
      RECT  3.19 1.355 3.29 1.49 ;
    END
    ANTENNADIFFAREA 0.659 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.24 1.54 0.34 ;
      RECT  0.845 0.34 0.965 0.44 ;
      RECT  0.28 0.44 0.965 0.545 ;
      RECT  0.065 1.21 2.29 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  1.83 1.46 3.1 1.56 ;
  END
END SEN_AOI211_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_4
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_4
  CLASS CORE ;
  FOREIGN SEN_AOI211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.815 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.21 0.19 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.56 1.415 0.73 1.75 ;
      RECT  1.08 1.415 1.25 1.75 ;
      RECT  1.6 1.415 1.77 1.75 ;
      RECT  2.12 1.415 2.255 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.82 0.05 0.99 0.32 ;
      RECT  0.28 0.05 0.49 0.325 ;
      RECT  2.565 0.05 2.735 0.34 ;
      RECT  3.085 0.05 3.255 0.34 ;
      RECT  3.605 0.05 3.775 0.34 ;
      RECT  4.125 0.05 4.295 0.34 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.41 0.34 4.53 0.445 ;
      RECT  1.34 0.445 4.53 0.56 ;
      RECT  3.55 0.56 3.65 1.11 ;
      RECT  3.55 1.11 4.255 1.29 ;
    END
    ANTENNADIFFAREA 0.832 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.19 2.32 0.325 ;
      RECT  1.105 0.325 1.225 0.44 ;
      RECT  0.065 0.34 0.185 0.44 ;
      RECT  0.065 0.44 1.225 0.56 ;
      RECT  1.975 0.91 2.715 1.03 ;
      RECT  1.975 1.03 2.095 1.2 ;
      RECT  2.585 1.03 2.715 1.245 ;
      RECT  0.325 1.2 2.095 1.325 ;
      RECT  2.585 1.245 3.29 1.36 ;
      RECT  0.325 1.325 0.44 1.42 ;
      RECT  2.325 1.14 2.45 1.32 ;
      RECT  2.345 1.32 2.45 1.45 ;
      RECT  2.345 1.45 4.53 1.565 ;
      RECT  4.405 1.34 4.53 1.45 ;
  END
END SEN_AOI211_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_0P75
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_0P75
  CLASS CORE ;
  FOREIGN SEN_AOI211_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.635 1.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.68 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.355 1.44 0.48 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.95 0.05 1.08 0.365 ;
      RECT  0.075 0.05 0.205 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.615 0.22 0.85 0.34 ;
      RECT  0.75 0.34 0.85 0.455 ;
      RECT  0.75 0.455 1.335 0.545 ;
      RECT  1.215 0.24 1.335 0.455 ;
      RECT  0.95 0.545 1.05 1.31 ;
      RECT  0.95 1.31 1.335 1.49 ;
    END
    ANTENNADIFFAREA 0.188 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.085 1.26 0.66 1.35 ;
      RECT  0.57 1.35 0.66 1.44 ;
      RECT  0.085 1.35 0.205 1.48 ;
      RECT  0.57 1.44 0.835 1.56 ;
  END
END SEN_AOI211_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_12
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_12
  CLASS CORE ;
  FOREIGN SEN_AOI211_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 5.85 0.765 ;
      RECT  2.95 0.765 5.85 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7257 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 2.45 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7257 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.91 0.71 11.85 0.89 ;
      RECT  11.75 0.89 11.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.693 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.71 8.85 0.89 ;
      RECT  8.75 0.89 8.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.693 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 12.6 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  1.88 1.44 2.01 1.75 ;
      RECT  2.38 1.48 2.55 1.75 ;
      RECT  2.9 1.485 3.07 1.75 ;
      RECT  3.44 1.44 3.57 1.75 ;
      RECT  3.96 1.44 4.09 1.75 ;
      RECT  4.48 1.44 4.61 1.75 ;
      RECT  5.0 1.44 5.13 1.75 ;
      RECT  5.52 1.44 5.65 1.75 ;
      RECT  6.04 1.44 6.17 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.6 0.05 ;
      RECT  6.325 0.05 6.51 0.305 ;
      RECT  6.89 0.05 7.07 0.305 ;
      RECT  7.41 0.05 7.58 0.305 ;
      RECT  7.925 0.05 8.1 0.305 ;
      RECT  8.45 0.05 8.665 0.305 ;
      RECT  8.97 0.05 9.14 0.305 ;
      RECT  9.53 0.05 9.7 0.32 ;
      RECT  1.88 0.05 2.01 0.345 ;
      RECT  2.4 0.05 2.53 0.345 ;
      RECT  2.92 0.05 3.045 0.35 ;
      RECT  10.07 0.05 10.2 0.36 ;
      RECT  10.59 0.05 10.72 0.36 ;
      RECT  11.11 0.05 11.24 0.36 ;
      RECT  11.63 0.05 11.76 0.36 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      RECT  0.29 0.05 0.41 0.59 ;
      RECT  12.185 0.05 12.305 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.025 0.395 9.375 0.405 ;
      RECT  5.5 0.405 9.375 0.42 ;
      RECT  5.5 0.42 9.97 0.44 ;
      RECT  3.42 0.44 9.97 0.45 ;
      RECT  3.42 0.45 12.065 0.58 ;
      RECT  3.42 0.58 10.49 0.6 ;
      RECT  8.95 0.6 10.49 0.62 ;
      RECT  5.95 0.6 6.85 0.69 ;
      RECT  8.95 0.62 9.78 0.69 ;
      RECT  9.55 0.69 9.78 1.1 ;
      RECT  9.55 1.1 10.85 1.205 ;
      RECT  9.55 1.205 12.325 1.3 ;
      RECT  10.57 1.3 12.325 1.335 ;
    END
    ANTENNADIFFAREA 2.137 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.135 0.155 3.85 0.19 ;
      RECT  3.135 0.19 5.96 0.315 ;
      RECT  3.135 0.315 4.9 0.35 ;
      RECT  3.135 0.35 3.33 0.45 ;
      RECT  1.59 0.45 3.33 0.48 ;
      RECT  0.53 0.48 3.33 0.61 ;
      RECT  2.635 0.61 3.33 0.645 ;
      RECT  3.15 1.085 7.06 1.125 ;
      RECT  3.15 1.125 7.58 1.155 ;
      RECT  3.15 1.155 8.105 1.18 ;
      RECT  1.61 1.18 9.17 1.21 ;
      RECT  0.065 1.21 9.17 1.315 ;
      RECT  0.065 1.315 3.33 1.33 ;
      RECT  2.12 1.33 3.33 1.365 ;
      RECT  0.065 1.33 0.185 1.43 ;
      RECT  2.64 1.365 3.33 1.395 ;
      RECT  12.415 1.33 12.535 1.425 ;
      RECT  6.605 1.425 12.535 1.545 ;
      RECT  7.67 1.545 11.0 1.61 ;
      RECT  8.71 1.61 9.92 1.64 ;
  END
END SEN_AOI211_12
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_6
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_6
  CLASS CORE ;
  FOREIGN SEN_AOI211_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.85 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3618 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.45 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3618 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.71 6.25 0.89 ;
      RECT  6.15 0.89 6.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3465 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.675 4.65 0.89 ;
      RECT  4.55 0.89 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3456 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.44 0.465 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.855 1.44 0.985 1.75 ;
      RECT  1.375 1.44 1.505 1.75 ;
      RECT  1.895 1.44 2.025 1.75 ;
      RECT  2.415 1.44 2.545 1.75 ;
      RECT  2.98 1.44 3.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  3.805 0.05 3.935 0.345 ;
      RECT  4.325 0.05 4.455 0.345 ;
      RECT  4.845 0.05 4.975 0.345 ;
      RECT  5.365 0.05 5.495 0.345 ;
      RECT  5.885 0.05 6.015 0.345 ;
      RECT  1.375 0.05 1.505 0.37 ;
      RECT  0.335 0.05 0.465 0.385 ;
      RECT  0.855 0.05 0.985 0.385 ;
      RECT  6.405 0.05 6.53 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.85 0.435 6.32 0.565 ;
      RECT  4.95 0.565 6.32 0.58 ;
      RECT  4.95 0.58 5.25 0.69 ;
      RECT  5.12 0.69 5.25 1.215 ;
      RECT  5.12 1.215 6.32 1.335 ;
    END
    ANTENNADIFFAREA 1.077 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.62 0.23 3.43 0.345 ;
      RECT  1.62 0.345 1.76 0.465 ;
      RECT  1.085 0.465 1.76 0.495 ;
      RECT  0.08 0.38 0.2 0.495 ;
      RECT  0.08 0.495 1.76 0.615 ;
      RECT  0.08 1.23 4.685 1.35 ;
      RECT  0.08 1.35 0.2 1.45 ;
      RECT  6.41 1.375 6.53 1.455 ;
      RECT  3.68 1.455 6.53 1.575 ;
  END
END SEN_AOI211_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_8
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_8
  CLASS CORE ;
  FOREIGN SEN_AOI211_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4833 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4833 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.645 0.71 7.85 0.89 ;
      RECT  7.75 0.89 7.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4623 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4623 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  1.88 1.44 2.01 1.75 ;
      RECT  2.4 1.44 2.53 1.75 ;
      RECT  2.92 1.44 3.05 1.75 ;
      RECT  3.44 1.44 3.57 1.75 ;
      RECT  3.96 1.44 4.09 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  4.28 0.05 4.41 0.36 ;
      RECT  4.83 0.05 4.96 0.36 ;
      RECT  5.35 0.05 5.48 0.36 ;
      RECT  5.87 0.05 6.0 0.36 ;
      RECT  6.39 0.05 6.52 0.36 ;
      RECT  6.91 0.05 7.04 0.36 ;
      RECT  7.43 0.05 7.56 0.36 ;
      RECT  7.95 0.05 8.08 0.36 ;
      RECT  1.88 0.05 2.01 0.37 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  0.29 0.05 0.41 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.135 0.31 6.255 0.45 ;
      RECT  2.37 0.45 8.335 0.58 ;
      RECT  8.215 0.34 8.335 0.45 ;
      RECT  3.95 0.58 6.52 0.62 ;
      RECT  3.95 0.62 4.45 0.69 ;
      RECT  5.75 0.62 6.52 0.69 ;
      RECT  6.35 0.69 6.52 1.11 ;
      RECT  6.35 1.11 6.65 1.21 ;
      RECT  6.35 1.21 8.125 1.34 ;
    END
    ANTENNADIFFAREA 1.412 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.13 0.21 2.81 0.24 ;
      RECT  2.13 0.24 3.875 0.36 ;
      RECT  2.13 0.36 2.28 0.465 ;
      RECT  1.59 0.465 2.28 0.495 ;
      RECT  0.535 0.495 2.28 0.615 ;
      RECT  2.1 1.18 4.98 1.22 ;
      RECT  0.065 1.22 4.98 1.23 ;
      RECT  0.065 1.23 6.05 1.35 ;
      RECT  0.065 1.35 0.185 1.44 ;
      RECT  8.215 1.34 8.335 1.44 ;
      RECT  4.52 1.44 8.335 1.56 ;
      RECT  5.59 1.56 6.81 1.59 ;
  END
END SEN_AOI211_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_G_0P5
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_G_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI211_G_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.755 ;
      RECT  0.125 0.755 0.25 0.925 ;
      RECT  0.15 0.925 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.635 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.68 0.68 0.85 ;
      RECT  0.55 0.85 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.42 0.44 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.76 0.05 0.89 0.365 ;
      RECT  0.055 0.05 0.18 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.455 0.22 0.65 0.34 ;
      RECT  0.55 0.34 0.65 0.455 ;
      RECT  0.55 0.455 1.145 0.545 ;
      RECT  1.025 0.275 1.145 0.455 ;
      RECT  0.77 0.545 0.86 0.91 ;
      RECT  0.75 0.91 0.86 1.23 ;
      RECT  0.75 1.23 1.05 1.32 ;
      RECT  0.95 1.32 1.05 1.395 ;
      RECT  0.95 1.395 1.145 1.565 ;
    END
    ANTENNADIFFAREA 0.125 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 1.24 0.64 1.33 ;
      RECT  0.55 1.33 0.64 1.42 ;
      RECT  0.055 1.33 0.175 1.465 ;
      RECT  0.55 1.42 0.75 1.54 ;
  END
END SEN_AOI211_G_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_G_0P75
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_G_0P75
  CLASS CORE ;
  FOREIGN SEN_AOI211_G_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.635 1.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.68 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.35 1.44 0.48 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.95 0.05 1.08 0.365 ;
      RECT  0.07 0.05 0.2 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.615 0.22 0.85 0.34 ;
      RECT  0.75 0.34 0.85 0.455 ;
      RECT  0.75 0.455 1.335 0.545 ;
      RECT  1.215 0.325 1.335 0.455 ;
      RECT  0.95 0.545 1.05 1.31 ;
      RECT  0.95 1.31 1.335 1.49 ;
    END
    ANTENNADIFFAREA 0.218 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.085 1.26 0.66 1.35 ;
      RECT  0.57 1.35 0.66 1.44 ;
      RECT  0.085 1.35 0.205 1.48 ;
      RECT  0.57 1.44 0.83 1.56 ;
  END
END SEN_AOI211_G_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_G_1
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_G_1
  CLASS CORE ;
  FOREIGN SEN_AOI211_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.635 1.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.68 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.35 1.44 0.48 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.95 0.05 1.08 0.365 ;
      RECT  0.07 0.05 0.2 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.615 0.22 0.85 0.34 ;
      RECT  0.75 0.34 0.85 0.455 ;
      RECT  0.75 0.455 1.335 0.545 ;
      RECT  1.215 0.325 1.335 0.455 ;
      RECT  0.95 0.545 1.05 1.31 ;
      RECT  0.95 1.31 1.335 1.49 ;
    END
    ANTENNADIFFAREA 0.295 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.085 1.26 0.66 1.35 ;
      RECT  0.57 1.35 0.66 1.44 ;
      RECT  0.085 1.35 0.205 1.48 ;
      RECT  0.57 1.44 0.84 1.56 ;
  END
END SEN_AOI211_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_G_2
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_G_2
  CLASS CORE ;
  FOREIGN SEN_AOI211_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.35 0.05 1.48 0.36 ;
      RECT  1.88 0.05 2.01 0.36 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  2.415 0.05 2.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.795 0.455 2.325 0.575 ;
      RECT  1.95 0.575 2.05 1.22 ;
      RECT  1.95 1.22 2.31 1.34 ;
    END
    ANTENNADIFFAREA 0.408 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.24 1.26 0.36 ;
      RECT  0.585 0.36 0.705 0.49 ;
      RECT  0.065 0.37 0.185 0.49 ;
      RECT  0.065 0.49 0.705 0.59 ;
      RECT  0.275 1.23 1.785 1.35 ;
      RECT  1.33 1.44 2.535 1.56 ;
      RECT  2.415 1.56 2.535 1.63 ;
  END
END SEN_AOI211_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_G_3
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_G_3
  CLASS CORE ;
  FOREIGN SEN_AOI211_G_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  1.88 0.05 2.01 0.36 ;
      RECT  2.4 0.05 2.53 0.36 ;
      RECT  2.935 0.05 3.065 0.36 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.215 0.355 3.335 0.455 ;
      RECT  1.055 0.455 3.335 0.575 ;
      RECT  2.55 0.575 2.65 1.22 ;
      RECT  2.55 1.22 3.335 1.34 ;
      RECT  3.215 1.34 3.335 1.445 ;
    END
    ANTENNADIFFAREA 0.677 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.24 1.535 0.36 ;
      RECT  0.845 0.36 0.965 0.495 ;
      RECT  0.275 0.495 0.965 0.615 ;
      RECT  0.065 1.23 2.315 1.35 ;
      RECT  0.065 1.35 0.185 1.45 ;
      RECT  1.83 1.44 3.115 1.56 ;
  END
END SEN_AOI211_G_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_G_4
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_G_4
  CLASS CORE ;
  FOREIGN SEN_AOI211_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.44 0.44 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.83 1.44 0.96 1.75 ;
      RECT  1.35 1.44 1.48 1.75 ;
      RECT  1.87 1.44 2.0 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.6 0.05 2.73 0.36 ;
      RECT  3.12 0.05 3.25 0.36 ;
      RECT  3.64 0.05 3.77 0.36 ;
      RECT  4.16 0.05 4.29 0.36 ;
      RECT  0.31 0.05 0.44 0.385 ;
      RECT  0.83 0.05 0.96 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.305 0.455 4.545 0.575 ;
      RECT  2.345 0.575 2.46 0.72 ;
      RECT  4.425 0.575 4.545 0.72 ;
      RECT  3.55 0.575 3.65 1.22 ;
      RECT  3.55 1.22 4.32 1.34 ;
    END
    ANTENNADIFFAREA 0.844 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.135 0.17 2.255 0.24 ;
      RECT  1.095 0.24 2.255 0.36 ;
      RECT  1.095 0.36 1.215 0.495 ;
      RECT  0.055 0.18 0.175 0.495 ;
      RECT  0.055 0.495 1.215 0.615 ;
      RECT  2.135 0.96 2.255 1.23 ;
      RECT  0.055 1.23 3.295 1.35 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  2.295 1.44 4.545 1.56 ;
      RECT  4.425 1.56 4.545 1.63 ;
  END
END SEN_AOI211_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_G_5
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_G_5
  CLASS CORE ;
  FOREIGN SEN_AOI211_G_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.45 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 5.25 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.85 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  1.91 1.44 2.04 1.75 ;
      RECT  2.485 1.44 2.615 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  3.03 0.05 3.16 0.36 ;
      RECT  3.55 0.05 3.68 0.36 ;
      RECT  4.09 0.05 4.22 0.36 ;
      RECT  4.63 0.05 4.76 0.36 ;
      RECT  5.15 0.05 5.28 0.36 ;
      RECT  1.1 0.05 1.23 0.37 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.415 0.35 5.535 0.45 ;
      RECT  1.575 0.45 5.535 0.57 ;
      RECT  4.35 0.57 4.45 1.22 ;
      RECT  4.35 1.22 5.535 1.34 ;
      RECT  5.415 1.34 5.535 1.44 ;
    END
    ANTENNADIFFAREA 1.085 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.365 0.24 2.66 0.36 ;
      RECT  1.365 0.36 1.485 0.495 ;
      RECT  0.275 0.495 1.485 0.615 ;
      RECT  0.065 1.225 3.985 1.345 ;
      RECT  0.065 1.345 0.185 1.445 ;
      RECT  2.98 1.44 5.325 1.56 ;
  END
END SEN_AOI211_G_5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI211_G_8
#      Description : "One 2-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI211_G_8
  CLASS CORE ;
  FOREIGN SEN_AOI211_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.045 0.71 8.25 0.89 ;
      RECT  8.15 0.89 8.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.905 0.71 6.05 0.89 ;
      RECT  5.95 0.89 6.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  1.88 1.44 2.01 1.75 ;
      RECT  2.4 1.44 2.53 1.75 ;
      RECT  2.92 1.44 3.05 1.75 ;
      RECT  3.44 1.44 3.57 1.75 ;
      RECT  3.96 1.44 4.09 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  4.46 0.05 4.58 0.36 ;
      RECT  4.97 0.05 5.1 0.36 ;
      RECT  5.49 0.05 5.62 0.36 ;
      RECT  6.01 0.05 6.14 0.36 ;
      RECT  6.53 0.05 6.66 0.36 ;
      RECT  7.05 0.05 7.18 0.36 ;
      RECT  7.57 0.05 7.7 0.36 ;
      RECT  8.09 0.05 8.22 0.36 ;
      RECT  1.88 0.05 2.01 0.37 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  8.615 0.05 8.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.37 0.45 4.12 0.51 ;
      RECT  2.37 0.51 8.525 0.58 ;
      RECT  4.49 0.45 8.525 0.51 ;
      RECT  3.95 0.58 6.92 0.62 ;
      RECT  3.95 0.62 4.67 0.69 ;
      RECT  6.15 0.62 6.92 0.69 ;
      RECT  6.75 0.69 6.92 1.11 ;
      RECT  6.75 1.11 7.05 1.21 ;
      RECT  6.75 1.21 8.525 1.34 ;
    END
    ANTENNADIFFAREA 1.632 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.13 0.21 2.81 0.24 ;
      RECT  2.13 0.24 4.37 0.36 ;
      RECT  2.13 0.36 2.28 0.465 ;
      RECT  1.59 0.465 2.28 0.495 ;
      RECT  0.065 0.385 0.185 0.495 ;
      RECT  0.065 0.495 2.28 0.615 ;
      RECT  2.1 1.18 5.38 1.22 ;
      RECT  0.065 1.22 5.38 1.23 ;
      RECT  0.065 1.23 6.445 1.35 ;
      RECT  0.065 1.35 0.185 1.44 ;
      RECT  8.615 1.34 8.735 1.44 ;
      RECT  4.405 1.44 8.735 1.56 ;
      RECT  5.99 1.56 7.21 1.59 ;
  END
END SEN_AOI211_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_0P5
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI21_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.69 0.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.385 1.43 0.505 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.67 0.05 0.79 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.085 0.24 0.45 0.36 ;
      RECT  0.35 0.36 0.45 0.455 ;
      RECT  0.35 0.455 1.06 0.545 ;
      RECT  0.94 0.275 1.06 0.455 ;
      RECT  0.94 0.545 1.06 1.5 ;
    END
    ANTENNADIFFAREA 0.124 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.11 1.24 0.79 1.33 ;
      RECT  0.11 1.33 0.23 1.53 ;
      RECT  0.67 1.33 0.79 1.53 ;
  END
END SEN_AOI21_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_1
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_1
  CLASS CORE ;
  FOREIGN SEN_AOI21_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.69 0.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.385 1.45 0.505 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.67 0.05 0.79 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.085 0.24 0.45 0.36 ;
      RECT  0.35 0.36 0.45 0.455 ;
      RECT  0.35 0.455 1.06 0.545 ;
      RECT  0.94 0.3 1.06 0.455 ;
      RECT  0.94 0.545 1.06 1.5 ;
    END
    ANTENNADIFFAREA 0.25 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.085 1.24 0.83 1.36 ;
  END
END SEN_AOI21_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_2
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_2
  CLASS CORE ;
  FOREIGN SEN_AOI21_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.78 1.85 0.885 ;
      RECT  1.75 0.885 1.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.45 0.445 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.845 1.45 0.965 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.325 0.05 0.445 0.35 ;
      RECT  1.565 0.05 1.685 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.82 0.51 1.945 0.62 ;
      RECT  1.15 0.62 1.945 0.69 ;
      RECT  1.35 0.69 1.45 1.385 ;
      RECT  1.35 1.385 1.71 1.48 ;
    END
    ANTENNADIFFAREA 0.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.24 1.25 0.36 ;
      RECT  0.585 0.36 0.705 0.44 ;
      RECT  0.065 0.34 0.185 0.44 ;
      RECT  0.065 0.44 0.705 0.56 ;
      RECT  0.065 1.24 1.26 1.36 ;
      RECT  0.065 1.36 0.19 1.46 ;
      RECT  1.14 1.36 1.26 1.57 ;
      RECT  1.14 1.57 1.945 1.66 ;
      RECT  1.825 1.41 1.945 1.57 ;
  END
END SEN_AOI21_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_3
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_3
  CLASS CORE ;
  FOREIGN SEN_AOI21_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.5 2.45 0.71 ;
      RECT  2.14 0.71 2.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.455 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.85 1.45 0.97 1.75 ;
      RECT  1.37 1.45 1.49 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.59 0.05 0.71 0.35 ;
      RECT  1.89 0.05 2.01 0.35 ;
      RECT  2.41 0.05 2.53 0.39 ;
      RECT  0.07 0.05 0.19 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.31 2.26 0.445 ;
      RECT  1.08 0.445 2.26 0.56 ;
      RECT  1.95 0.56 2.05 1.11 ;
      RECT  1.89 1.11 2.53 1.29 ;
    END
    ANTENNADIFFAREA 0.504 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.85 0.24 1.55 0.355 ;
      RECT  0.85 0.355 0.97 0.44 ;
      RECT  0.305 0.44 0.97 0.56 ;
      RECT  0.07 1.24 1.75 1.36 ;
      RECT  1.63 1.36 1.75 1.44 ;
      RECT  0.07 1.36 0.19 1.46 ;
      RECT  1.63 1.44 2.32 1.56 ;
  END
END SEN_AOI21_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_4
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_4
  CLASS CORE ;
  FOREIGN SEN_AOI21_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.85 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.45 0.435 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.835 1.45 0.955 1.75 ;
      RECT  1.355 1.45 1.475 1.75 ;
      RECT  1.875 1.455 1.995 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.835 0.05 0.955 0.35 ;
      RECT  0.315 0.05 0.435 0.36 ;
      RECT  2.385 0.05 2.505 0.39 ;
      RECT  2.905 0.05 3.025 0.39 ;
      RECT  3.425 0.05 3.545 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.33 0.5 3.34 0.62 ;
      RECT  1.95 0.62 2.85 0.69 ;
      RECT  2.75 0.69 2.85 1.11 ;
      RECT  2.645 1.11 3.25 1.2 ;
      RECT  2.645 1.2 3.31 1.29 ;
    END
    ANTENNADIFFAREA 0.624 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.1 0.24 2.28 0.36 ;
      RECT  1.1 0.36 1.215 0.45 ;
      RECT  0.055 0.45 1.215 0.56 ;
      RECT  0.055 0.56 0.175 0.69 ;
      RECT  0.055 1.24 2.39 1.36 ;
      RECT  2.27 1.36 2.39 1.465 ;
      RECT  0.055 1.36 0.175 1.63 ;
      RECT  2.27 1.465 3.545 1.585 ;
      RECT  3.425 1.41 3.545 1.465 ;
  END
END SEN_AOI21_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_16
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_16
  CLASS CORE ;
  FOREIGN SEN_AOI21_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.76 0.71 8.06 0.9 ;
      RECT  6.605 0.71 6.905 0.9 ;
      RECT  5.825 0.71 6.125 0.9 ;
      RECT  4.735 0.71 5.035 0.9 ;
      RECT  3.75 0.71 4.125 0.9 ;
      RECT  2.635 0.71 2.975 0.9 ;
      RECT  1.615 0.71 1.915 0.9 ;
      RECT  0.62 0.71 0.98 0.9 ;
      LAYER M2 ;
      RECT  0.795 0.75 8.29 0.85 ;
      LAYER V1 ;
      RECT  7.76 0.75 7.86 0.85 ;
      RECT  7.96 0.75 8.06 0.85 ;
      RECT  6.605 0.75 6.705 0.85 ;
      RECT  6.805 0.75 6.905 0.85 ;
      RECT  5.825 0.75 5.925 0.85 ;
      RECT  6.025 0.75 6.125 0.85 ;
      RECT  4.735 0.75 4.835 0.85 ;
      RECT  4.935 0.75 5.035 0.85 ;
      RECT  3.825 0.75 3.925 0.85 ;
      RECT  4.025 0.75 4.125 0.85 ;
      RECT  2.675 0.75 2.775 0.85 ;
      RECT  2.875 0.75 2.975 0.85 ;
      RECT  1.615 0.75 1.715 0.85 ;
      RECT  1.815 0.75 1.915 0.85 ;
      RECT  0.835 0.75 0.935 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.755 8.335 0.91 ;
      RECT  8.15 0.91 8.565 1.09 ;
      RECT  7.315 0.755 7.415 0.91 ;
      RECT  7.11 0.91 7.415 1.09 ;
      RECT  6.39 0.755 6.515 0.91 ;
      RECT  6.215 0.91 6.515 1.09 ;
      RECT  5.35 0.755 5.475 0.91 ;
      RECT  5.175 0.91 5.475 1.09 ;
      RECT  4.315 0.755 4.415 0.91 ;
      RECT  4.315 0.91 4.645 1.09 ;
      RECT  3.275 0.755 3.395 0.91 ;
      RECT  3.275 0.91 3.605 1.09 ;
      RECT  2.15 0.745 2.25 0.91 ;
      RECT  2.15 0.91 2.455 1.09 ;
      RECT  1.145 0.735 1.255 0.91 ;
      RECT  1.145 0.91 1.455 1.09 ;
      RECT  0.15 0.71 0.275 0.91 ;
      RECT  0.15 0.91 0.455 1.09 ;
      LAYER M2 ;
      RECT  0.275 0.95 8.49 1.05 ;
      LAYER V1 ;
      RECT  8.15 0.95 8.25 1.05 ;
      RECT  8.35 0.95 8.45 1.05 ;
      RECT  7.11 0.95 7.21 1.05 ;
      RECT  7.31 0.95 7.41 1.05 ;
      RECT  6.215 0.95 6.315 1.05 ;
      RECT  6.415 0.95 6.515 1.05 ;
      RECT  5.175 0.95 5.275 1.05 ;
      RECT  5.375 0.95 5.475 1.05 ;
      RECT  4.345 0.95 4.445 1.05 ;
      RECT  4.545 0.95 4.645 1.05 ;
      RECT  3.305 0.95 3.405 1.05 ;
      RECT  3.505 0.95 3.605 1.05 ;
      RECT  2.15 0.95 2.25 1.05 ;
      RECT  2.35 0.95 2.45 1.05 ;
      RECT  1.15 0.95 1.25 1.05 ;
      RECT  1.35 0.95 1.45 1.05 ;
      RECT  0.315 0.95 0.415 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.02 0.71 12.65 0.89 ;
      RECT  12.55 0.89 12.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  0.82 1.48 0.99 1.75 ;
      RECT  1.34 1.48 1.51 1.75 ;
      RECT  1.86 1.48 2.03 1.75 ;
      RECT  2.38 1.48 2.55 1.75 ;
      RECT  2.9 1.48 3.07 1.75 ;
      RECT  3.42 1.48 3.59 1.75 ;
      RECT  3.94 1.48 4.11 1.75 ;
      RECT  4.46 1.48 4.63 1.75 ;
      RECT  4.98 1.48 5.15 1.75 ;
      RECT  5.5 1.48 5.67 1.75 ;
      RECT  6.02 1.48 6.19 1.75 ;
      RECT  6.54 1.48 6.71 1.75 ;
      RECT  7.06 1.48 7.23 1.75 ;
      RECT  7.58 1.48 7.75 1.75 ;
      RECT  8.125 1.44 8.25 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  1.08 0.05 1.25 0.305 ;
      RECT  2.12 0.05 2.29 0.305 ;
      RECT  3.16 0.05 3.33 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  5.24 0.05 5.41 0.305 ;
      RECT  6.28 0.05 6.45 0.305 ;
      RECT  7.32 0.05 7.49 0.305 ;
      RECT  8.4 0.05 8.57 0.305 ;
      RECT  8.95 0.05 9.12 0.305 ;
      RECT  9.47 0.05 9.64 0.305 ;
      RECT  9.99 0.05 10.16 0.305 ;
      RECT  10.51 0.05 10.68 0.305 ;
      RECT  11.03 0.05 11.2 0.305 ;
      RECT  11.55 0.05 11.72 0.305 ;
      RECT  12.07 0.05 12.24 0.305 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  12.615 0.05 12.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.6 0.35 0.83 0.415 ;
      RECT  0.6 0.415 12.475 0.59 ;
      RECT  1.6 0.35 1.98 0.415 ;
      RECT  2.64 0.35 3.02 0.415 ;
      RECT  3.68 0.35 4.06 0.415 ;
      RECT  4.72 0.35 5.1 0.415 ;
      RECT  5.76 0.35 6.14 0.415 ;
      RECT  6.8 0.35 7.18 0.415 ;
      RECT  7.84 0.35 8.22 0.415 ;
      RECT  8.68 0.35 8.86 0.415 ;
      RECT  9.2 0.35 9.38 0.415 ;
      RECT  9.73 0.35 9.91 0.415 ;
      RECT  10.25 0.35 10.43 0.415 ;
      RECT  10.77 0.35 10.95 0.415 ;
      RECT  11.285 0.35 11.465 0.415 ;
      RECT  6.84 0.59 6.93 0.6 ;
      RECT  8.55 0.59 12.475 0.6 ;
      RECT  8.55 0.6 9.85 0.69 ;
      RECT  9.55 0.69 9.85 1.07 ;
      RECT  9.55 1.07 12.46 1.11 ;
      RECT  12.365 1.01 12.46 1.07 ;
      RECT  8.73 1.11 12.46 1.19 ;
      RECT  8.73 1.19 11.46 1.29 ;
      LAYER M2 ;
      RECT  0.645 0.35 11.465 0.45 ;
      LAYER V1 ;
      RECT  0.685 0.35 0.785 0.45 ;
      RECT  1.64 0.35 1.74 0.45 ;
      RECT  1.84 0.35 1.94 0.45 ;
      RECT  2.68 0.35 2.78 0.45 ;
      RECT  2.88 0.35 2.98 0.45 ;
      RECT  3.72 0.35 3.82 0.45 ;
      RECT  3.92 0.35 4.02 0.45 ;
      RECT  4.76 0.35 4.86 0.45 ;
      RECT  4.96 0.35 5.06 0.45 ;
      RECT  5.8 0.35 5.9 0.45 ;
      RECT  6.0 0.35 6.1 0.45 ;
      RECT  6.84 0.35 6.94 0.45 ;
      RECT  7.04 0.35 7.14 0.45 ;
      RECT  7.88 0.35 7.98 0.45 ;
      RECT  8.08 0.35 8.18 0.45 ;
      RECT  8.72 0.35 8.82 0.45 ;
      RECT  9.24 0.35 9.34 0.45 ;
      RECT  9.77 0.35 9.87 0.45 ;
      RECT  10.29 0.35 10.39 0.45 ;
      RECT  10.81 0.35 10.91 0.45 ;
      RECT  11.325 0.35 11.425 0.45 ;
    END
    ANTENNADIFFAREA 2.496 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 1.18 8.64 1.35 ;
      RECT  0.08 1.35 7.975 1.37 ;
      RECT  8.34 1.35 8.64 1.43 ;
      RECT  2.66 1.37 2.76 1.49 ;
      RECT  3.195 1.37 3.295 1.49 ;
      RECT  3.715 1.37 3.815 1.49 ;
      RECT  4.235 1.37 4.335 1.49 ;
      RECT  4.75 1.37 4.85 1.49 ;
      RECT  5.27 1.37 5.37 1.49 ;
      RECT  7.355 1.37 7.455 1.49 ;
      RECT  7.875 1.37 7.975 1.49 ;
      RECT  8.34 1.43 12.72 1.64 ;
      RECT  11.685 1.35 12.72 1.43 ;
      LAYER M2 ;
      RECT  2.62 1.35 12.465 1.45 ;
      LAYER V1 ;
      RECT  2.66 1.35 2.76 1.45 ;
      RECT  3.195 1.35 3.295 1.45 ;
      RECT  3.715 1.35 3.815 1.45 ;
      RECT  4.235 1.35 4.335 1.45 ;
      RECT  4.75 1.35 4.85 1.45 ;
      RECT  5.27 1.35 5.37 1.45 ;
      RECT  7.355 1.35 7.455 1.45 ;
      RECT  7.875 1.35 7.975 1.45 ;
      RECT  8.34 1.35 8.44 1.45 ;
      RECT  8.54 1.35 8.64 1.45 ;
      RECT  11.725 1.35 11.825 1.45 ;
      RECT  11.925 1.35 12.025 1.45 ;
      RECT  12.125 1.35 12.225 1.45 ;
      RECT  12.325 1.35 12.425 1.45 ;
  END
END SEN_AOI21_16
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_6
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_6
  CLASS CORE ;
  FOREIGN SEN_AOI21_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.495 0.71 2.795 0.9 ;
      RECT  1.635 0.71 1.935 0.9 ;
      RECT  0.705 0.71 1.05 0.93 ;
      LAYER M2 ;
      RECT  0.71 0.75 3.09 0.85 ;
      LAYER V1 ;
      RECT  2.495 0.75 2.595 0.85 ;
      RECT  2.695 0.75 2.795 0.85 ;
      RECT  1.635 0.75 1.735 0.85 ;
      RECT  1.835 0.75 1.935 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
      RECT  0.95 0.75 1.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.095 0.755 3.185 0.91 ;
      RECT  2.885 0.91 3.185 1.09 ;
      RECT  2.105 0.75 2.195 0.91 ;
      RECT  2.105 0.91 2.405 1.09 ;
      RECT  1.19 0.755 1.29 0.91 ;
      RECT  1.19 0.91 1.49 1.09 ;
      RECT  0.15 0.71 0.275 0.91 ;
      RECT  0.15 0.91 0.615 1.09 ;
      LAYER M2 ;
      RECT  0.275 0.95 3.29 1.05 ;
      LAYER V1 ;
      RECT  2.885 0.95 2.985 1.05 ;
      RECT  3.085 0.95 3.185 1.05 ;
      RECT  2.105 0.95 2.205 1.05 ;
      RECT  2.305 0.95 2.405 1.05 ;
      RECT  1.19 0.95 1.29 1.05 ;
      RECT  1.39 0.95 1.49 1.05 ;
      RECT  0.315 0.95 0.415 1.05 ;
      RECT  0.515 0.95 0.615 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.84 0.71 4.85 0.89 ;
      RECT  4.75 0.89 4.85 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.495 0.47 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.82 1.495 0.99 1.75 ;
      RECT  1.34 1.495 1.51 1.75 ;
      RECT  1.86 1.495 2.03 1.75 ;
      RECT  2.38 1.495 2.55 1.75 ;
      RECT  2.9 1.495 3.07 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  1.08 0.05 1.25 0.305 ;
      RECT  2.12 0.05 2.29 0.305 ;
      RECT  3.16 0.05 3.33 0.305 ;
      RECT  3.68 0.05 3.85 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  4.76 0.05 4.88 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.545 0.43 4.645 0.56 ;
      RECT  0.545 0.56 3.68 0.57 ;
      RECT  3.55 0.57 3.68 1.11 ;
      RECT  3.445 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.936 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.235 3.31 1.365 ;
      RECT  0.065 1.365 0.185 1.455 ;
      RECT  3.16 1.365 3.31 1.48 ;
      RECT  3.16 1.48 4.865 1.61 ;
      RECT  4.75 1.41 4.865 1.48 ;
  END
END SEN_AOI21_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_8
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_8
  CLASS CORE ;
  FOREIGN SEN_AOI21_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.63 0.71 3.93 0.9 ;
      RECT  2.68 0.71 3.085 0.9 ;
      RECT  1.65 0.71 2.045 0.9 ;
      RECT  0.705 0.71 1.135 0.9 ;
      LAYER M2 ;
      RECT  0.795 0.75 4.09 0.85 ;
      LAYER V1 ;
      RECT  3.63 0.75 3.73 0.85 ;
      RECT  3.83 0.75 3.93 0.85 ;
      RECT  2.785 0.75 2.885 0.85 ;
      RECT  2.985 0.75 3.085 0.85 ;
      RECT  1.705 0.75 1.805 0.85 ;
      RECT  1.945 0.75 2.045 0.85 ;
      RECT  0.835 0.75 0.935 0.85 ;
      RECT  1.035 0.75 1.135 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.11 0.755 4.225 0.91 ;
      RECT  4.11 0.91 4.41 1.09 ;
      RECT  3.24 0.755 3.33 0.91 ;
      RECT  3.24 0.91 3.54 1.09 ;
      RECT  2.265 0.755 2.355 0.91 ;
      RECT  2.265 0.91 2.565 1.09 ;
      RECT  1.225 0.725 1.33 0.91 ;
      RECT  1.225 0.91 1.525 1.09 ;
      RECT  0.15 0.71 0.275 0.91 ;
      RECT  0.15 0.91 0.615 1.09 ;
      LAYER M2 ;
      RECT  0.275 0.95 4.49 1.05 ;
      LAYER V1 ;
      RECT  4.11 0.95 4.21 1.05 ;
      RECT  4.31 0.95 4.41 1.05 ;
      RECT  3.24 0.95 3.34 1.05 ;
      RECT  3.44 0.95 3.54 1.05 ;
      RECT  2.265 0.95 2.365 1.05 ;
      RECT  2.465 0.95 2.565 1.05 ;
      RECT  1.225 0.95 1.325 1.05 ;
      RECT  1.425 0.95 1.525 1.05 ;
      RECT  0.315 0.95 0.415 1.05 ;
      RECT  0.515 0.95 0.615 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.035 0.71 6.45 0.9 ;
      RECT  6.35 0.9 6.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.495 0.47 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.82 1.495 0.99 1.75 ;
      RECT  1.34 1.495 1.51 1.75 ;
      RECT  1.86 1.495 2.03 1.75 ;
      RECT  2.38 1.495 2.55 1.75 ;
      RECT  2.9 1.495 3.07 1.75 ;
      RECT  3.42 1.495 3.59 1.75 ;
      RECT  3.94 1.495 4.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.08 0.05 1.25 0.305 ;
      RECT  2.12 0.05 2.29 0.305 ;
      RECT  3.16 0.05 3.33 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.72 0.05 4.89 0.305 ;
      RECT  5.24 0.05 5.41 0.305 ;
      RECT  5.76 0.05 5.93 0.305 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.33 0.05 6.45 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.415 6.17 0.585 ;
      RECT  4.75 0.585 4.93 1.11 ;
      RECT  4.5 1.11 6.17 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.215 4.38 1.385 ;
      RECT  4.2 1.385 4.38 1.415 ;
      RECT  4.2 1.415 6.425 1.585 ;
  END
END SEN_AOI21_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_G_6
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_G_6
  CLASS CORE ;
  FOREIGN SEN_AOI21_G_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.495 0.71 2.795 0.9 ;
      RECT  1.67 0.71 2.015 0.895 ;
      RECT  0.705 0.71 1.135 0.925 ;
      LAYER M2 ;
      RECT  0.795 0.75 3.09 0.85 ;
      LAYER V1 ;
      RECT  2.495 0.75 2.595 0.85 ;
      RECT  2.695 0.75 2.795 0.85 ;
      RECT  1.715 0.75 1.815 0.85 ;
      RECT  1.915 0.75 2.015 0.85 ;
      RECT  0.835 0.75 0.935 0.85 ;
      RECT  1.035 0.75 1.135 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.095 0.755 3.185 0.91 ;
      RECT  2.885 0.91 3.185 1.09 ;
      RECT  2.105 0.755 2.195 0.91 ;
      RECT  2.105 0.91 2.405 1.09 ;
      RECT  1.225 0.755 1.325 0.91 ;
      RECT  1.225 0.91 1.525 1.09 ;
      RECT  0.15 0.71 0.275 0.91 ;
      RECT  0.15 0.91 0.615 1.09 ;
      LAYER M2 ;
      RECT  0.275 0.95 3.29 1.05 ;
      LAYER V1 ;
      RECT  2.885 0.95 2.985 1.05 ;
      RECT  3.085 0.95 3.185 1.05 ;
      RECT  2.105 0.95 2.205 1.05 ;
      RECT  2.305 0.95 2.405 1.05 ;
      RECT  1.225 0.95 1.325 1.05 ;
      RECT  1.425 0.95 1.525 1.05 ;
      RECT  0.315 0.95 0.415 1.05 ;
      RECT  0.515 0.95 0.615 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.82 0.71 4.85 0.89 ;
      RECT  4.75 0.89 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.495 0.47 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.82 1.495 0.99 1.75 ;
      RECT  1.34 1.495 1.51 1.75 ;
      RECT  1.86 1.495 2.03 1.75 ;
      RECT  2.38 1.495 2.55 1.75 ;
      RECT  2.9 1.495 3.07 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  1.08 0.05 1.25 0.305 ;
      RECT  2.12 0.05 2.29 0.305 ;
      RECT  3.16 0.05 3.33 0.305 ;
      RECT  3.68 0.05 3.85 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  4.76 0.05 4.88 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.545 0.43 4.65 0.56 ;
      RECT  0.545 0.56 3.68 0.57 ;
      RECT  3.55 0.57 3.68 1.11 ;
      RECT  3.445 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.936 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.23 3.31 1.37 ;
      RECT  0.065 1.37 0.185 1.45 ;
      RECT  3.16 1.37 3.31 1.48 ;
      RECT  3.16 1.48 4.865 1.61 ;
      RECT  4.75 1.38 4.865 1.48 ;
  END
END SEN_AOI21_G_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_G_8
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_G_8
  CLASS CORE ;
  FOREIGN SEN_AOI21_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.63 0.71 3.93 0.9 ;
      RECT  2.725 0.71 3.085 0.925 ;
      RECT  1.665 0.71 2.045 0.9 ;
      RECT  0.705 0.71 1.135 0.94 ;
      LAYER M2 ;
      RECT  0.795 0.75 4.09 0.85 ;
      LAYER V1 ;
      RECT  3.63 0.75 3.73 0.85 ;
      RECT  3.83 0.75 3.93 0.85 ;
      RECT  2.785 0.75 2.885 0.85 ;
      RECT  2.985 0.75 3.085 0.85 ;
      RECT  1.705 0.75 1.805 0.85 ;
      RECT  1.945 0.75 2.045 0.85 ;
      RECT  0.835 0.75 0.935 0.85 ;
      RECT  1.035 0.75 1.135 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.11 0.755 4.225 0.91 ;
      RECT  4.11 0.91 4.41 1.09 ;
      RECT  3.24 0.755 3.33 0.91 ;
      RECT  3.24 0.91 3.54 1.09 ;
      RECT  2.235 0.755 2.325 0.91 ;
      RECT  2.235 0.91 2.565 1.09 ;
      RECT  1.225 0.755 1.325 0.91 ;
      RECT  1.225 0.91 1.525 1.09 ;
      RECT  0.15 0.71 0.275 0.91 ;
      RECT  0.15 0.91 0.615 1.09 ;
      LAYER M2 ;
      RECT  0.275 0.95 4.49 1.05 ;
      LAYER V1 ;
      RECT  4.11 0.95 4.21 1.05 ;
      RECT  4.31 0.95 4.41 1.05 ;
      RECT  3.24 0.95 3.34 1.05 ;
      RECT  3.44 0.95 3.54 1.05 ;
      RECT  2.265 0.95 2.365 1.05 ;
      RECT  2.465 0.95 2.565 1.05 ;
      RECT  1.225 0.95 1.325 1.05 ;
      RECT  1.425 0.95 1.525 1.05 ;
      RECT  0.315 0.95 0.415 1.05 ;
      RECT  0.515 0.95 0.615 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.095 0.71 6.45 0.9 ;
      RECT  6.35 0.9 6.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.495 0.47 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.82 1.495 0.99 1.75 ;
      RECT  1.34 1.495 1.51 1.75 ;
      RECT  1.86 1.495 2.03 1.75 ;
      RECT  2.38 1.495 2.55 1.75 ;
      RECT  2.9 1.495 3.07 1.75 ;
      RECT  3.42 1.495 3.59 1.75 ;
      RECT  3.94 1.495 4.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.08 0.05 1.25 0.305 ;
      RECT  2.12 0.05 2.29 0.305 ;
      RECT  3.16 0.05 3.33 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.72 0.05 4.89 0.305 ;
      RECT  5.24 0.05 5.41 0.305 ;
      RECT  5.76 0.05 5.93 0.305 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.33 0.05 6.45 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.415 6.17 0.585 ;
      RECT  4.75 0.585 4.92 1.11 ;
      RECT  4.5 1.11 6.17 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.215 4.38 1.385 ;
      RECT  4.2 1.385 4.38 1.415 ;
      RECT  2.68 1.385 2.77 1.42 ;
      RECT  4.2 1.415 6.44 1.585 ;
  END
END SEN_AOI21_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_S_0P5
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_S_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI21_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.41 0.46 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  1.0 0.05 1.13 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.63 0.235 0.85 0.355 ;
      RECT  0.75 0.355 0.85 1.18 ;
      RECT  0.75 1.18 1.1 1.32 ;
      RECT  0.95 1.32 1.1 1.53 ;
    END
    ANTENNADIFFAREA 0.096 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.21 0.64 1.3 ;
      RECT  0.55 1.3 0.64 1.465 ;
      RECT  0.065 1.3 0.185 1.53 ;
      RECT  0.55 1.465 0.85 1.585 ;
  END
END SEN_AOI21_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_S_1
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_S_1
  CLASS CORE ;
  FOREIGN SEN_AOI21_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0474 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.46 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.98 0.05 1.11 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.63 0.235 0.85 0.355 ;
      RECT  0.75 0.355 0.85 1.18 ;
      RECT  0.75 1.18 1.1 1.32 ;
      RECT  0.95 1.32 1.1 1.49 ;
    END
    ANTENNADIFFAREA 0.169 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.2 0.64 1.29 ;
      RECT  0.065 1.29 0.185 1.42 ;
      RECT  0.55 1.29 0.64 1.465 ;
      RECT  0.55 1.465 0.84 1.585 ;
  END
END SEN_AOI21_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_S_2
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_S_2
  CLASS CORE ;
  FOREIGN SEN_AOI21_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0948 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.84 1.44 0.965 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  1.35 0.05 1.46 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.845 0.33 0.965 0.47 ;
      RECT  0.845 0.47 1.73 0.555 ;
      RECT  1.55 0.31 1.73 0.47 ;
      RECT  0.845 0.555 1.65 0.56 ;
      RECT  1.55 0.56 1.65 1.18 ;
      RECT  1.34 1.18 1.65 1.3 ;
    END
    ANTENNADIFFAREA 0.239 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.15 1.225 0.24 ;
      RECT  1.105 0.24 1.225 0.38 ;
      RECT  0.585 0.24 0.705 0.47 ;
      RECT  0.065 0.26 0.185 0.47 ;
      RECT  0.065 0.47 0.705 0.56 ;
      RECT  0.065 1.23 1.225 1.35 ;
      RECT  0.065 1.35 0.185 1.45 ;
      RECT  1.105 1.35 1.225 1.52 ;
      RECT  1.105 1.52 1.75 1.61 ;
      RECT  1.625 1.41 1.75 1.52 ;
  END
END SEN_AOI21_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_S_4
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_S_4
  CLASS CORE ;
  FOREIGN SEN_AOI21_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.695 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2133 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.695 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2133 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.73 0.695 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1896 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.36 1.41 1.49 1.75 ;
      RECT  1.88 1.41 2.01 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  2.39 0.05 2.52 0.39 ;
      RECT  2.91 0.05 3.04 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.885 0.325 2.005 0.495 ;
      RECT  1.885 0.495 2.775 0.505 ;
      RECT  2.655 0.215 2.775 0.495 ;
      RECT  1.365 0.33 1.485 0.505 ;
      RECT  1.365 0.505 3.295 0.595 ;
      RECT  3.15 0.22 3.295 0.505 ;
      RECT  2.35 0.595 2.45 1.11 ;
      RECT  2.35 1.11 3.05 1.29 ;
    END
    ANTENNADIFFAREA 0.447 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.145 2.265 0.235 ;
      RECT  1.625 0.235 1.745 0.39 ;
      RECT  2.145 0.235 2.265 0.39 ;
      RECT  1.105 0.235 1.225 0.475 ;
      RECT  0.065 0.26 0.185 0.475 ;
      RECT  0.065 0.475 1.225 0.575 ;
      RECT  0.585 0.26 0.705 0.475 ;
      RECT  0.065 1.21 2.26 1.32 ;
      RECT  2.145 1.32 2.26 1.38 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  2.145 1.38 3.305 1.5 ;
      RECT  3.185 1.5 3.305 1.6 ;
  END
END SEN_AOI21_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_S_8
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_S_8
  CLASS CORE ;
  FOREIGN SEN_AOI21_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4275 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4275 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.81 0.71 6.45 0.89 ;
      RECT  6.35 0.89 6.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3792 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.845 1.255 0.965 1.75 ;
      RECT  1.365 1.255 1.485 1.75 ;
      RECT  1.885 1.255 2.005 1.75 ;
      RECT  2.405 1.255 2.525 1.75 ;
      RECT  2.925 1.255 3.045 1.75 ;
      RECT  3.445 1.255 3.565 1.75 ;
      RECT  3.96 1.44 4.085 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  4.45 0.05 4.62 0.335 ;
      RECT  4.97 0.05 5.14 0.34 ;
      RECT  5.49 0.05 5.66 0.34 ;
      RECT  6.01 0.05 6.18 0.34 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      RECT  1.88 0.05 2.01 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.71 0.3 4.88 0.43 ;
      RECT  4.71 0.43 6.45 0.45 ;
      RECT  5.23 0.3 5.4 0.43 ;
      RECT  5.75 0.3 5.92 0.43 ;
      RECT  6.295 0.21 6.45 0.43 ;
      RECT  2.38 0.37 2.55 0.41 ;
      RECT  2.38 0.41 4.11 0.45 ;
      RECT  2.9 0.37 3.07 0.41 ;
      RECT  3.42 0.37 3.59 0.41 ;
      RECT  3.94 0.37 4.11 0.41 ;
      RECT  2.38 0.45 6.45 0.57 ;
      RECT  2.38 0.57 4.72 0.58 ;
      RECT  4.0 0.58 4.72 0.62 ;
      RECT  4.55 0.62 4.72 1.11 ;
      RECT  4.55 1.11 6.165 1.18 ;
      RECT  4.46 1.18 6.165 1.29 ;
    END
    ANTENNADIFFAREA 0.877 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.13 0.14 4.36 0.28 ;
      RECT  2.64 0.28 2.81 0.32 ;
      RECT  3.16 0.28 3.33 0.32 ;
      RECT  3.68 0.28 3.85 0.32 ;
      RECT  4.215 0.28 4.36 0.36 ;
      RECT  2.13 0.28 2.28 0.48 ;
      RECT  0.065 0.26 0.185 0.48 ;
      RECT  0.065 0.48 2.28 0.62 ;
      RECT  0.585 0.26 0.705 0.48 ;
      RECT  1.105 0.26 1.225 0.48 ;
      RECT  1.625 0.26 1.745 0.48 ;
      RECT  0.54 1.005 3.85 1.165 ;
      RECT  3.68 1.165 3.85 1.18 ;
      RECT  0.54 1.165 0.665 1.21 ;
      RECT  3.68 1.18 4.37 1.35 ;
      RECT  0.065 1.21 0.665 1.325 ;
      RECT  0.065 1.325 0.185 1.43 ;
      RECT  4.2 1.35 4.37 1.44 ;
      RECT  4.2 1.44 6.48 1.6 ;
  END
END SEN_AOI21_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_0P75
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_0P75
  CLASS CORE ;
  FOREIGN SEN_AOI21_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.425 1.05 0.98 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.465 0.47 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.84 0.05 1.01 0.335 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.69 0.485 ;
      RECT  0.55 0.485 0.85 0.575 ;
      RECT  0.75 0.575 0.85 1.11 ;
      RECT  0.75 1.11 1.05 1.21 ;
      RECT  0.855 1.21 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.141 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.285 0.695 1.375 ;
      RECT  0.07 1.375 0.18 1.505 ;
      RECT  0.595 1.375 0.695 1.51 ;
  END
END SEN_AOI21_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_0P5
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.5 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.9 ;
      RECT  0.35 0.9 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.035 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.475 0.47 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.885 0.05 1.015 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.23 0.69 0.48 ;
      RECT  0.55 0.48 0.85 0.58 ;
      RECT  0.75 0.58 0.85 1.125 ;
      RECT  0.75 1.125 1.05 1.215 ;
      RECT  0.87 1.215 1.05 1.53 ;
    END
    ANTENNADIFFAREA 0.101 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.295 0.705 1.385 ;
      RECT  0.585 1.385 0.705 1.515 ;
      RECT  0.065 1.385 0.185 1.52 ;
  END
END SEN_AOI21_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_1
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_1
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.82 1.48 0.99 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.28 0.05 0.42 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.27 1.05 1.055 ;
      RECT  0.95 1.055 1.485 1.145 ;
      RECT  1.35 1.145 1.485 1.49 ;
    END
    ANTENNADIFFAREA 0.308 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.255 1.22 1.375 ;
      RECT  0.065 1.375 0.185 1.485 ;
      RECT  1.105 1.375 1.22 1.485 ;
  END
END SEN_AOI21_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_12
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_12
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.55 0.69 11.65 0.89 ;
      RECT  11.55 0.89 11.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2096 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.69 ;
      RECT  0.15 0.69 4.51 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2096 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.945 0.71 14.25 0.89 ;
      RECT  14.15 0.89 14.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.756 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.27 0.47 1.75 ;
      RECT  0.0 1.75 14.4 1.85 ;
      RECT  0.82 1.27 0.99 1.75 ;
      RECT  1.34 1.27 1.51 1.75 ;
      RECT  1.86 1.27 2.03 1.75 ;
      RECT  2.38 1.44 2.55 1.75 ;
      RECT  2.9 1.435 3.07 1.75 ;
      RECT  3.42 1.44 3.59 1.75 ;
      RECT  3.94 1.44 4.11 1.75 ;
      RECT  4.46 1.44 4.63 1.75 ;
      RECT  4.98 1.44 5.15 1.75 ;
      RECT  5.5 1.44 5.67 1.75 ;
      RECT  6.02 1.44 6.19 1.75 ;
      RECT  6.54 1.44 6.71 1.75 ;
      RECT  7.06 1.44 7.23 1.75 ;
      RECT  7.58 1.44 7.75 1.75 ;
      RECT  8.1 1.44 8.27 1.75 ;
      RECT  8.62 1.44 8.79 1.75 ;
      RECT  9.14 1.44 9.31 1.75 ;
      RECT  9.66 1.46 9.83 1.75 ;
      RECT  10.18 1.46 10.35 1.75 ;
      RECT  10.7 1.46 10.87 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 14.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 14.4 0.05 ;
      RECT  11.33 0.05 11.5 0.32 ;
      RECT  11.85 0.05 12.02 0.32 ;
      RECT  12.37 0.05 12.54 0.32 ;
      RECT  12.89 0.05 13.06 0.32 ;
      RECT  13.41 0.05 13.58 0.32 ;
      RECT  13.93 0.05 14.1 0.32 ;
      RECT  0.56 0.05 0.73 0.335 ;
      RECT  1.08 0.05 1.25 0.335 ;
      RECT  1.6 0.05 1.77 0.335 ;
      RECT  2.12 0.05 2.29 0.335 ;
      RECT  2.64 0.05 2.81 0.335 ;
      RECT  3.16 0.05 3.33 0.335 ;
      RECT  3.68 0.05 3.85 0.335 ;
      RECT  4.2 0.05 4.37 0.335 ;
      RECT  4.72 0.05 4.89 0.335 ;
      RECT  5.24 0.05 5.41 0.335 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 14.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.88 0.395 9.05 0.445 ;
      RECT  8.88 0.445 14.335 0.465 ;
      RECT  9.4 0.395 9.57 0.445 ;
      RECT  9.92 0.395 10.09 0.445 ;
      RECT  10.44 0.395 10.61 0.445 ;
      RECT  10.97 0.24 11.12 0.445 ;
      RECT  11.61 0.305 11.74 0.445 ;
      RECT  12.125 0.305 12.27 0.445 ;
      RECT  14.215 0.33 14.335 0.445 ;
      RECT  7.345 0.355 7.45 0.465 ;
      RECT  7.345 0.465 14.335 0.555 ;
      RECT  7.83 0.35 8.01 0.465 ;
      RECT  8.35 0.35 8.53 0.465 ;
      RECT  7.345 0.555 12.79 0.565 ;
      RECT  7.345 0.565 7.45 0.6 ;
      RECT  12.15 0.565 12.79 0.69 ;
      RECT  5.75 0.385 5.93 0.6 ;
      RECT  5.75 0.6 7.45 0.7 ;
      RECT  6.28 0.395 6.45 0.6 ;
      RECT  6.8 0.395 6.97 0.6 ;
      RECT  12.15 0.69 12.45 1.11 ;
      RECT  11.75 1.11 14.06 1.18 ;
      RECT  11.35 1.015 11.46 1.18 ;
      RECT  11.35 1.18 14.06 1.29 ;
      LAYER M2 ;
      RECT  7.83 0.35 12.295 0.45 ;
      LAYER V1 ;
      RECT  7.87 0.35 7.97 0.45 ;
      RECT  8.39 0.35 8.49 0.45 ;
      RECT  10.995 0.35 11.095 0.45 ;
      RECT  11.625 0.35 11.725 0.45 ;
      RECT  12.15 0.35 12.25 0.45 ;
    END
    ANTENNADIFFAREA 1.906 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.51 0.15 10.88 0.26 ;
      RECT  5.51 0.26 7.23 0.285 ;
      RECT  9.14 0.26 10.88 0.285 ;
      RECT  7.61 0.26 7.72 0.375 ;
      RECT  8.13 0.26 8.24 0.375 ;
      RECT  8.645 0.26 8.765 0.375 ;
      RECT  5.51 0.285 5.66 0.425 ;
      RECT  6.56 0.285 6.69 0.49 ;
      RECT  7.06 0.285 7.23 0.49 ;
      RECT  6.05 0.285 6.16 0.495 ;
      RECT  10.7 0.285 10.88 0.335 ;
      RECT  9.14 0.285 9.31 0.35 ;
      RECT  9.66 0.285 9.83 0.355 ;
      RECT  10.18 0.285 10.35 0.355 ;
      RECT  0.34 0.28 0.44 0.425 ;
      RECT  0.34 0.425 5.66 0.575 ;
      RECT  0.85 0.28 0.96 0.425 ;
      RECT  1.37 0.28 1.48 0.425 ;
      RECT  1.89 0.28 2.0 0.425 ;
      RECT  2.41 0.28 2.52 0.425 ;
      RECT  2.93 0.28 3.04 0.425 ;
      RECT  3.45 0.28 3.56 0.425 ;
      RECT  3.97 0.28 4.08 0.425 ;
      RECT  4.49 0.28 4.6 0.425 ;
      RECT  5.01 0.28 5.12 0.425 ;
      RECT  0.065 1.0 11.255 1.17 ;
      RECT  0.065 1.17 0.185 1.23 ;
      RECT  2.355 1.17 11.255 1.25 ;
      RECT  10.98 1.25 11.255 1.4 ;
      RECT  10.98 1.4 14.32 1.64 ;
      LAYER M2 ;
      RECT  3.94 0.35 7.235 0.45 ;
      LAYER V1 ;
      RECT  3.98 0.35 4.08 0.45 ;
      RECT  4.5 0.35 4.6 0.45 ;
      RECT  5.015 0.35 5.115 0.45 ;
      RECT  5.55 0.35 5.65 0.45 ;
      RECT  6.055 0.35 6.155 0.45 ;
      RECT  6.575 0.35 6.675 0.45 ;
      RECT  7.095 0.35 7.195 0.45 ;
  END
END SEN_AOI21_T_12
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_1P5
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_1P5
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1506 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.31 0.25 0.71 ;
      RECT  0.15 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1506 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  1.94 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.43 0.45 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.84 1.43 0.97 1.75 ;
      RECT  1.34 1.475 1.51 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.56 0.05 0.73 0.335 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.145 0.05 2.275 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.9 0.3 2.05 0.45 ;
      RECT  1.065 0.45 2.05 0.54 ;
      RECT  1.065 0.54 1.85 0.56 ;
      RECT  1.75 0.56 1.85 1.01 ;
      RECT  1.75 1.01 2.05 1.1 ;
      RECT  1.875 1.1 2.05 1.375 ;
    END
    ANTENNADIFFAREA 0.234 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.85 0.22 1.53 0.33 ;
      RECT  0.85 0.33 0.96 0.445 ;
      RECT  0.34 0.325 0.445 0.445 ;
      RECT  0.34 0.445 0.96 0.545 ;
      RECT  0.07 1.205 1.74 1.325 ;
      RECT  0.07 1.325 0.185 1.43 ;
      RECT  1.63 1.325 1.74 1.505 ;
      RECT  1.63 1.505 2.265 1.595 ;
      RECT  2.155 1.375 2.265 1.505 ;
  END
END SEN_AOI21_T_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_2
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_2
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.665 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.85 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.44 0.71 2.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.24 0.45 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.845 1.24 0.97 1.75 ;
      RECT  1.365 1.225 1.495 1.75 ;
      RECT  1.86 1.495 2.03 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  2.145 0.05 2.265 0.36 ;
      RECT  0.83 0.05 0.98 0.385 ;
      RECT  2.665 0.05 2.785 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.405 0.19 2.525 0.45 ;
      RECT  1.485 0.45 2.525 0.55 ;
      RECT  2.15 0.55 2.25 1.055 ;
      RECT  2.15 1.055 2.65 1.165 ;
      RECT  2.55 1.165 2.65 1.29 ;
    END
    ANTENNADIFFAREA 0.436 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.11 0.215 2.04 0.335 ;
      RECT  1.11 0.335 1.22 0.53 ;
      RECT  0.585 0.44 0.71 0.53 ;
      RECT  0.585 0.53 1.22 0.62 ;
      RECT  0.065 0.995 1.745 1.125 ;
      RECT  1.625 1.125 1.745 1.28 ;
      RECT  0.065 1.125 0.18 1.285 ;
      RECT  1.625 1.28 2.26 1.37 ;
      RECT  2.15 1.37 2.26 1.425 ;
      RECT  2.15 1.425 2.81 1.545 ;
  END
END SEN_AOI21_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_3
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_3
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.205 0.61 2.85 0.725 ;
      RECT  2.75 0.725 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3024 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.305 0.45 0.71 ;
      RECT  0.35 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3024 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.65 0.93 ;
      RECT  3.55 0.93 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.189 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.57 1.44 0.72 1.75 ;
      RECT  1.09 1.44 1.24 1.75 ;
      RECT  1.61 1.44 1.76 1.75 ;
      RECT  2.13 1.44 2.28 1.75 ;
      RECT  2.64 1.47 2.81 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.83 0.05 1.0 0.33 ;
      RECT  3.17 0.05 3.34 0.33 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.74 0.05 3.86 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.34 0.32 1.51 0.42 ;
      RECT  1.34 0.42 3.6 0.51 ;
      RECT  1.86 0.32 2.03 0.42 ;
      RECT  2.38 0.32 2.55 0.42 ;
      RECT  2.93 0.24 3.05 0.42 ;
      RECT  3.15 0.51 3.6 0.54 ;
      RECT  3.15 0.54 3.25 1.24 ;
      RECT  3.15 1.24 3.85 1.355 ;
      RECT  3.715 1.355 3.85 1.5 ;
    END
    ANTENNADIFFAREA 0.524 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.12 0.14 2.81 0.23 ;
      RECT  1.6 0.23 1.77 0.33 ;
      RECT  2.12 0.23 2.29 0.33 ;
      RECT  2.64 0.23 2.81 0.33 ;
      RECT  1.12 0.23 1.23 0.45 ;
      RECT  0.54 0.45 1.23 0.575 ;
      RECT  0.3 1.22 3.055 1.34 ;
      RECT  2.935 1.34 3.055 1.465 ;
      RECT  2.935 1.465 3.615 1.585 ;
  END
END SEN_AOI21_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_4
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_4
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.63 3.65 0.74 ;
      RECT  3.55 0.74 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.65 1.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.85 0.89 ;
      RECT  4.75 0.89 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.465 0.47 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.82 1.24 0.99 1.75 ;
      RECT  1.34 1.24 1.51 1.75 ;
      RECT  1.86 1.24 2.03 1.75 ;
      RECT  2.38 1.24 2.55 1.75 ;
      RECT  2.9 1.235 3.07 1.75 ;
      RECT  3.42 1.465 3.59 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  3.94 0.05 4.11 0.33 ;
      RECT  4.46 0.05 4.63 0.33 ;
      RECT  0.56 0.05 0.73 0.335 ;
      RECT  1.08 0.05 1.25 0.335 ;
      RECT  1.6 0.05 1.77 0.335 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.12 0.335 2.29 0.42 ;
      RECT  2.12 0.42 4.865 0.515 ;
      RECT  2.64 0.335 2.81 0.42 ;
      RECT  3.16 0.335 3.33 0.42 ;
      RECT  3.705 0.24 3.85 0.42 ;
      RECT  4.745 0.3 4.865 0.42 ;
      RECT  3.95 0.515 4.865 0.55 ;
      RECT  3.95 0.55 4.05 1.11 ;
      RECT  3.95 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.642 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.885 0.145 3.59 0.245 ;
      RECT  2.9 0.245 3.07 0.305 ;
      RECT  3.42 0.245 3.59 0.305 ;
      RECT  2.38 0.245 2.55 0.32 ;
      RECT  1.885 0.245 2.005 0.425 ;
      RECT  0.32 0.25 0.45 0.425 ;
      RECT  0.32 0.425 2.005 0.515 ;
      RECT  0.84 0.25 0.97 0.425 ;
      RECT  1.36 0.24 1.49 0.425 ;
      RECT  0.585 1.0 3.3 1.12 ;
      RECT  0.585 1.12 0.705 1.2 ;
      RECT  3.185 1.12 3.3 1.23 ;
      RECT  0.065 1.2 0.705 1.295 ;
      RECT  3.185 1.23 3.82 1.32 ;
      RECT  0.065 1.295 0.185 1.42 ;
      RECT  3.705 1.32 3.82 1.465 ;
      RECT  3.705 1.465 4.865 1.585 ;
      RECT  4.745 1.365 4.865 1.465 ;
  END
END SEN_AOI21_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_6
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_6
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.7 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 2.25 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6048 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.38 0.71 7.45 0.89 ;
      RECT  7.35 0.89 7.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.47 0.47 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  0.82 1.24 0.99 1.75 ;
      RECT  1.34 1.24 1.51 1.75 ;
      RECT  1.86 1.24 2.03 1.75 ;
      RECT  2.38 1.24 2.55 1.75 ;
      RECT  2.9 1.24 3.07 1.75 ;
      RECT  3.42 1.24 3.59 1.75 ;
      RECT  3.94 1.24 4.11 1.75 ;
      RECT  4.46 1.24 4.63 1.75 ;
      RECT  4.98 1.24 5.15 1.75 ;
      RECT  5.5 1.465 5.67 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  6.02 0.05 6.19 0.33 ;
      RECT  6.54 0.05 6.71 0.33 ;
      RECT  7.06 0.05 7.23 0.33 ;
      RECT  0.56 0.05 0.73 0.34 ;
      RECT  1.08 0.05 1.25 0.34 ;
      RECT  1.6 0.05 1.77 0.34 ;
      RECT  2.12 0.05 2.29 0.34 ;
      RECT  2.64 0.05 2.81 0.34 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.16 0.355 3.33 0.45 ;
      RECT  3.16 0.45 7.505 0.58 ;
      RECT  3.68 0.355 3.85 0.45 ;
      RECT  4.2 0.355 4.37 0.45 ;
      RECT  4.72 0.355 4.89 0.45 ;
      RECT  5.24 0.355 5.41 0.45 ;
      RECT  5.785 0.22 5.9 0.45 ;
      RECT  3.16 0.58 6.28 0.585 ;
      RECT  6.15 0.585 6.28 1.11 ;
      RECT  6.035 1.11 7.25 1.29 ;
    END
    ANTENNADIFFAREA 0.948 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.92 0.145 5.67 0.265 ;
      RECT  3.42 0.265 3.59 0.305 ;
      RECT  3.94 0.265 4.11 0.305 ;
      RECT  4.46 0.265 4.63 0.305 ;
      RECT  4.98 0.265 5.15 0.305 ;
      RECT  5.5 0.265 5.67 0.305 ;
      RECT  2.92 0.265 3.05 0.46 ;
      RECT  0.325 0.23 0.445 0.46 ;
      RECT  0.325 0.46 3.05 0.59 ;
      RECT  0.845 0.23 0.965 0.46 ;
      RECT  1.365 0.23 1.485 0.46 ;
      RECT  1.885 0.23 2.005 0.46 ;
      RECT  2.405 0.23 2.525 0.46 ;
      RECT  0.585 1.02 5.415 1.15 ;
      RECT  5.285 1.15 5.415 1.18 ;
      RECT  0.585 1.15 0.705 1.29 ;
      RECT  5.285 1.18 5.915 1.31 ;
      RECT  0.065 1.29 0.705 1.38 ;
      RECT  5.785 1.31 5.915 1.44 ;
      RECT  0.065 1.38 0.185 1.51 ;
      RECT  5.785 1.44 7.505 1.575 ;
  END
END SEN_AOI21_T_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_T_8
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_T_8
  CLASS CORE ;
  FOREIGN SEN_AOI21_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.02 0.71 7.65 0.89 ;
      RECT  7.55 0.89 7.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 2.54 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.06 0.71 9.85 0.89 ;
      RECT  9.75 0.89 9.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.465 0.47 1.75 ;
      RECT  0.0 1.75 10.0 1.85 ;
      RECT  0.82 1.24 0.99 1.75 ;
      RECT  1.34 1.24 1.51 1.75 ;
      RECT  1.86 1.24 2.03 1.75 ;
      RECT  2.38 1.24 2.55 1.75 ;
      RECT  2.9 1.24 3.07 1.75 ;
      RECT  3.42 1.24 3.59 1.75 ;
      RECT  3.94 1.24 4.11 1.75 ;
      RECT  4.46 1.24 4.63 1.75 ;
      RECT  4.98 1.24 5.15 1.75 ;
      RECT  5.5 1.24 5.67 1.75 ;
      RECT  6.02 1.24 6.19 1.75 ;
      RECT  6.54 1.25 6.71 1.75 ;
      RECT  7.06 1.47 7.23 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.0 0.05 ;
      RECT  7.615 0.05 7.745 0.36 ;
      RECT  8.135 0.05 8.265 0.36 ;
      RECT  8.655 0.05 8.785 0.36 ;
      RECT  9.175 0.05 9.305 0.36 ;
      RECT  0.3 0.05 0.47 0.37 ;
      RECT  0.82 0.05 0.99 0.37 ;
      RECT  1.34 0.05 1.51 0.37 ;
      RECT  1.86 0.05 2.03 0.37 ;
      RECT  2.38 0.05 2.55 0.37 ;
      RECT  2.9 0.05 3.07 0.37 ;
      RECT  3.42 0.05 3.59 0.37 ;
      RECT  9.72 0.05 9.84 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.06 0.41 7.23 0.45 ;
      RECT  7.06 0.45 9.575 0.47 ;
      RECT  3.94 0.43 4.11 0.47 ;
      RECT  3.94 0.47 9.575 0.62 ;
      RECT  4.46 0.43 4.63 0.47 ;
      RECT  4.98 0.43 5.15 0.47 ;
      RECT  5.5 0.43 5.67 0.47 ;
      RECT  6.02 0.43 6.19 0.47 ;
      RECT  6.54 0.41 6.71 0.47 ;
      RECT  3.94 0.62 4.85 0.69 ;
      RECT  7.75 0.62 7.92 1.11 ;
      RECT  7.75 1.11 9.65 1.29 ;
    END
    ANTENNADIFFAREA 1.224 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.68 0.16 7.49 0.32 ;
      RECT  4.2 0.32 4.37 0.36 ;
      RECT  4.72 0.32 4.89 0.36 ;
      RECT  5.24 0.32 5.41 0.36 ;
      RECT  5.76 0.32 5.93 0.36 ;
      RECT  6.28 0.32 6.45 0.36 ;
      RECT  6.8 0.32 6.97 0.36 ;
      RECT  7.32 0.32 7.49 0.36 ;
      RECT  3.68 0.32 3.85 0.46 ;
      RECT  0.065 0.26 0.185 0.46 ;
      RECT  0.065 0.46 3.85 0.59 ;
      RECT  0.585 0.27 0.705 0.46 ;
      RECT  1.105 0.3 1.225 0.46 ;
      RECT  1.625 0.3 1.745 0.46 ;
      RECT  2.145 0.3 2.265 0.46 ;
      RECT  2.665 0.3 2.785 0.46 ;
      RECT  3.185 0.3 3.305 0.46 ;
      RECT  0.585 0.98 7.0 1.15 ;
      RECT  6.83 1.15 7.0 1.18 ;
      RECT  0.585 1.15 0.7 1.21 ;
      RECT  6.83 1.18 7.495 1.35 ;
      RECT  0.065 1.21 0.7 1.315 ;
      RECT  0.065 1.315 0.185 1.43 ;
      RECT  7.32 1.35 7.495 1.415 ;
      RECT  7.32 1.415 9.82 1.585 ;
  END
END SEN_AOI21_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_G_0P5
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_G_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI21_G_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.66 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.255 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.255 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.985 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.485 0.545 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.115 0.05 0.245 0.39 ;
      RECT  0.945 0.05 1.075 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.615 0.215 0.85 0.335 ;
      RECT  0.75 0.335 0.85 1.075 ;
      RECT  0.75 1.075 1.05 1.185 ;
      RECT  0.93 1.185 1.05 1.53 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.135 1.305 0.785 1.395 ;
      RECT  0.135 1.395 0.26 1.53 ;
      RECT  0.665 1.395 0.785 1.53 ;
  END
END SEN_AOI21_G_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_G_0P75
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_G_0P75
  CLASS CORE ;
  FOREIGN SEN_AOI21_G_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.66 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.255 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.48 0.545 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.115 0.05 0.245 0.39 ;
      RECT  0.945 0.05 1.075 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.61 0.22 0.85 0.33 ;
      RECT  0.75 0.33 0.85 1.095 ;
      RECT  0.75 1.095 1.05 1.185 ;
      RECT  0.93 1.185 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.143 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.09 1.275 0.83 1.385 ;
  END
END SEN_AOI21_G_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_G_1
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_G_1
  CLASS CORE ;
  FOREIGN SEN_AOI21_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.66 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.51 0.255 0.71 ;
      RECT  0.145 0.71 0.45 0.9 ;
      RECT  0.145 0.9 0.255 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.51 1.05 0.93 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.465 0.545 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.115 0.05 0.245 0.39 ;
      RECT  0.955 0.05 1.085 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.605 0.24 0.85 0.36 ;
      RECT  0.75 0.36 0.85 1.025 ;
      RECT  0.75 1.025 1.05 1.115 ;
      RECT  0.925 1.115 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.095 1.255 0.835 1.375 ;
  END
END SEN_AOI21_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_G_2
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_G_2
  CLASS CORE ;
  FOREIGN SEN_AOI21_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.66 0.865 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.535 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.21 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.415 0.435 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.835 1.415 0.955 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.315 0.05 0.435 0.36 ;
      RECT  1.815 0.05 1.935 0.36 ;
      RECT  1.295 0.05 1.415 0.69 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.53 0.45 1.85 0.57 ;
      RECT  1.75 0.57 1.85 1.3 ;
      RECT  0.81 0.45 1.15 0.57 ;
      RECT  1.05 0.57 1.15 0.855 ;
      RECT  1.05 0.855 1.46 0.945 ;
      RECT  1.35 0.945 1.46 1.3 ;
      RECT  1.35 1.3 1.85 1.39 ;
    END
    ANTENNADIFFAREA 0.312 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.575 0.18 1.205 0.27 ;
      RECT  1.095 0.27 1.205 0.36 ;
      RECT  0.575 0.27 0.695 0.47 ;
      RECT  0.055 0.17 0.175 0.47 ;
      RECT  0.055 0.47 0.695 0.56 ;
      RECT  0.055 1.205 1.21 1.325 ;
      RECT  1.1 1.325 1.21 1.48 ;
      RECT  0.055 1.325 0.175 1.6 ;
      RECT  1.1 1.48 1.785 1.6 ;
  END
END SEN_AOI21_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_G_3
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_G_3
  CLASS CORE ;
  FOREIGN SEN_AOI21_G_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.9 ;
      RECT  1.55 0.9 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.9 ;
      RECT  0.55 0.9 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.5 2.45 0.71 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.36 1.41 1.49 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.88 0.05 2.01 0.36 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  2.395 0.05 2.53 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.145 0.3 2.25 0.47 ;
      RECT  1.055 0.47 2.25 0.59 ;
      RECT  1.95 0.59 2.05 1.11 ;
      RECT  1.86 1.11 2.25 1.215 ;
      RECT  1.86 1.215 2.525 1.315 ;
      RECT  2.405 1.315 2.525 1.465 ;
    END
    ANTENNADIFFAREA 0.504 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.255 1.535 0.375 ;
      RECT  0.845 0.375 0.965 0.5 ;
      RECT  0.325 0.37 0.445 0.5 ;
      RECT  0.325 0.5 0.965 0.59 ;
      RECT  0.065 1.21 1.745 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  1.625 1.32 1.745 1.48 ;
      RECT  1.625 1.48 2.315 1.6 ;
  END
END SEN_AOI21_G_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21_G_4
#      Description : "One 2-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21_G_4
  CLASS CORE ;
  FOREIGN SEN_AOI21_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.9 ;
      RECT  2.15 0.9 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.9 ;
      RECT  0.75 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.45 0.9 ;
      RECT  3.335 0.9 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.41 0.49 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.91 1.41 1.04 1.75 ;
      RECT  1.6 1.41 1.73 1.75 ;
      RECT  2.12 1.41 2.25 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.31 0.05 0.44 0.39 ;
      RECT  0.83 0.05 0.96 0.39 ;
      RECT  2.385 0.05 2.51 0.39 ;
      RECT  2.9 0.05 3.03 0.39 ;
      RECT  3.42 0.05 3.545 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.305 0.48 3.33 0.59 ;
      RECT  2.75 0.59 2.85 1.11 ;
      RECT  2.645 1.11 3.05 1.205 ;
      RECT  2.645 1.205 3.285 1.295 ;
      RECT  3.165 1.295 3.285 1.425 ;
    END
    ANTENNADIFFAREA 0.624 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.095 0.235 2.295 0.355 ;
      RECT  1.095 0.355 1.215 0.48 ;
      RECT  0.055 0.19 0.175 0.48 ;
      RECT  0.055 0.48 1.215 0.59 ;
      RECT  0.055 1.21 2.505 1.31 ;
      RECT  2.385 1.31 2.505 1.57 ;
      RECT  0.055 1.31 0.175 1.61 ;
      RECT  2.385 1.57 3.545 1.66 ;
      RECT  2.905 1.41 3.025 1.57 ;
      RECT  3.425 1.41 3.545 1.57 ;
  END
END SEN_AOI21_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21B_0P5
#      Description : "One 2-input AND into 2-input NOR (other input inverted)"
#      Equation    : X=!((A1&A2)|!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21B_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI21B_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 1.045 ;
      RECT  0.35 1.045 0.58 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.69 1.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.455 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.415 1.41 1.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  0.845 0.05 0.975 0.42 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.735 0.49 ;
      RECT  0.55 0.49 0.65 0.82 ;
      RECT  0.55 0.82 1.05 0.91 ;
      RECT  0.95 0.91 1.05 1.31 ;
      RECT  0.85 1.31 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.108 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.14 0.18 1.26 0.62 ;
      RECT  0.74 0.62 1.26 0.73 ;
      RECT  1.14 0.73 1.26 1.63 ;
      RECT  0.07 1.26 0.71 1.35 ;
      RECT  0.07 1.35 0.19 1.53 ;
      RECT  0.59 1.35 0.71 1.53 ;
  END
END SEN_AOI21B_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21B_1
#      Description : "One 2-input AND into 2-input NOR (other input inverted)"
#      Equation    : X=!((A1&A2)|!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21B_1
  CLASS CORE ;
  FOREIGN SEN_AOI21B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.505 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.35 1.41 0.495 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.39 1.435 1.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.095 0.05 0.215 0.39 ;
      RECT  1.0 0.05 1.16 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.58 0.24 0.85 0.36 ;
      RECT  0.75 0.36 0.85 1.0 ;
      RECT  0.75 1.0 1.05 1.09 ;
      RECT  0.89 1.09 1.05 1.3 ;
    END
    ANTENNADIFFAREA 0.192 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.41 0.22 1.51 0.5 ;
      RECT  1.155 0.5 1.51 0.59 ;
      RECT  1.155 0.59 1.255 0.79 ;
      RECT  0.99 0.79 1.255 0.89 ;
      RECT  1.15 0.89 1.255 1.55 ;
      RECT  0.09 1.21 0.76 1.3 ;
      RECT  0.09 1.3 0.22 1.43 ;
      RECT  0.63 1.3 0.76 1.43 ;
  END
END SEN_AOI21B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21B_2
#      Description : "One 2-input AND into 2-input NOR (other input inverted)"
#      Equation    : X=!((A1&A2)|!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21B_2
  CLASS CORE ;
  FOREIGN SEN_AOI21B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.475 0.47 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.82 1.475 0.99 1.75 ;
      RECT  2.245 1.41 2.355 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.85 0.05 2.02 0.35 ;
      RECT  1.35 0.05 1.475 0.37 ;
      RECT  2.4 0.05 2.515 0.39 ;
      RECT  0.3 0.05 0.47 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.82 0.465 1.76 0.59 ;
      RECT  1.35 0.59 1.45 1.0 ;
      RECT  1.35 1.0 1.485 1.17 ;
    END
    ANTENNADIFFAREA 0.312 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.16 1.21 0.25 ;
      RECT  1.105 0.25 1.21 0.375 ;
      RECT  0.585 0.25 0.705 0.5 ;
      RECT  0.06 0.37 0.19 0.5 ;
      RECT  0.06 0.5 0.705 0.59 ;
      RECT  2.13 0.22 2.25 0.5 ;
      RECT  1.86 0.5 2.25 0.59 ;
      RECT  1.86 0.59 1.95 0.79 ;
      RECT  1.605 0.79 1.95 0.9 ;
      RECT  1.86 0.9 1.95 1.155 ;
      RECT  1.86 1.155 1.995 1.33 ;
      RECT  0.065 1.26 1.77 1.375 ;
      RECT  0.065 1.375 0.185 1.48 ;
  END
END SEN_AOI21B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21B_3
#      Description : "One 2-input AND into 2-input NOR (other input inverted)"
#      Equation    : X=!((A1&A2)|!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21B_3
  CLASS CORE ;
  FOREIGN SEN_AOI21B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.695 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 0.71 ;
      RECT  2.87 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.45 0.47 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.82 1.45 0.99 1.75 ;
      RECT  1.34 1.45 1.51 1.75 ;
      RECT  2.555 1.45 2.745 1.75 ;
      RECT  3.125 1.235 3.245 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  1.87 0.05 2.015 0.345 ;
      RECT  0.58 0.05 0.71 0.375 ;
      RECT  3.115 0.05 3.25 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  2.45 0.05 2.57 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.08 0.44 2.32 0.56 ;
      RECT  1.95 0.56 2.05 1.11 ;
      RECT  1.89 1.11 2.55 1.29 ;
    END
    ANTENNADIFFAREA 0.488 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.225 1.54 0.345 ;
      RECT  0.845 0.345 0.965 0.465 ;
      RECT  0.3 0.465 0.965 0.585 ;
      RECT  2.67 0.43 3.0 0.55 ;
      RECT  2.67 0.55 2.77 0.79 ;
      RECT  2.165 0.79 2.77 0.89 ;
      RECT  2.67 0.89 2.77 1.24 ;
      RECT  2.67 1.24 2.995 1.355 ;
      RECT  0.065 1.24 1.74 1.36 ;
      RECT  1.63 1.36 1.74 1.445 ;
      RECT  0.065 1.36 0.185 1.46 ;
      RECT  1.63 1.445 2.32 1.555 ;
  END
END SEN_AOI21B_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21B_4
#      Description : "One 2-input AND into 2-input NOR (other input inverted)"
#      Equation    : X=!((A1&A2)|!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21B_4
  CLASS CORE ;
  FOREIGN SEN_AOI21B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.93 0.71 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1251 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.445 0.445 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.845 1.445 0.965 1.75 ;
      RECT  1.365 1.445 1.485 1.75 ;
      RECT  1.885 1.445 2.005 1.75 ;
      RECT  3.445 1.2 3.57 1.75 ;
      RECT  4.04 1.21 4.16 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.315 0.05 0.455 0.35 ;
      RECT  0.845 0.05 0.965 0.35 ;
      RECT  2.915 0.05 3.035 0.355 ;
      RECT  2.395 0.05 2.51 0.365 ;
      RECT  3.95 0.05 4.075 0.375 ;
      RECT  3.435 0.05 3.555 0.555 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.34 0.455 3.32 0.575 ;
      RECT  2.55 0.575 2.65 1.11 ;
      RECT  2.405 1.11 3.05 1.29 ;
    END
    ANTENNADIFFAREA 0.624 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.235 2.29 0.35 ;
      RECT  1.105 0.35 1.225 0.445 ;
      RECT  0.07 0.33 0.19 0.445 ;
      RECT  0.07 0.445 1.225 0.555 ;
      RECT  3.705 0.31 3.81 0.48 ;
      RECT  3.705 0.48 4.335 0.57 ;
      RECT  4.215 0.31 4.335 0.48 ;
      RECT  3.705 0.57 3.805 0.775 ;
      RECT  2.74 0.775 3.805 0.895 ;
      RECT  3.715 0.895 3.805 1.24 ;
      RECT  3.715 1.24 3.92 1.36 ;
      RECT  0.065 1.245 2.265 1.355 ;
      RECT  2.145 1.355 2.265 1.46 ;
      RECT  0.065 1.355 0.185 1.47 ;
      RECT  2.145 1.46 3.305 1.57 ;
      RECT  3.185 1.35 3.305 1.46 ;
  END
END SEN_AOI21B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI21B_8
#      Description : "One 2-input AND into 2-input NOR (other input inverted)"
#      Equation    : X=!((A1&A2)|!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI21B_8
  CLASS CORE ;
  FOREIGN SEN_AOI21B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.655 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.71 7.25 0.89 ;
      RECT  7.15 0.89 7.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.45 0.45 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  0.84 1.45 0.97 1.75 ;
      RECT  1.36 1.45 1.49 1.75 ;
      RECT  1.88 1.45 2.01 1.75 ;
      RECT  2.4 1.45 2.53 1.75 ;
      RECT  2.92 1.45 3.05 1.75 ;
      RECT  3.44 1.45 3.57 1.75 ;
      RECT  3.96 1.45 4.09 1.75 ;
      RECT  6.81 1.45 6.94 1.75 ;
      RECT  7.36 1.21 7.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  0.32 0.05 0.45 0.35 ;
      RECT  0.84 0.05 0.97 0.35 ;
      RECT  1.36 0.05 1.49 0.35 ;
      RECT  1.88 0.05 2.01 0.35 ;
      RECT  6.55 0.05 6.68 0.35 ;
      RECT  7.07 0.05 7.2 0.35 ;
      RECT  4.47 0.05 4.6 0.38 ;
      RECT  4.99 0.05 5.12 0.38 ;
      RECT  5.51 0.05 5.64 0.38 ;
      RECT  6.03 0.05 6.16 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.38 0.47 4.15 0.505 ;
      RECT  2.38 0.505 6.45 0.6 ;
      RECT  3.75 0.6 6.45 0.69 ;
      RECT  4.74 0.69 4.91 1.11 ;
      RECT  4.485 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.12 0.19 4.37 0.32 ;
      RECT  2.12 0.32 3.25 0.36 ;
      RECT  2.12 0.36 2.29 0.44 ;
      RECT  0.065 0.35 0.185 0.44 ;
      RECT  0.065 0.44 2.29 0.57 ;
      RECT  1.61 0.57 2.29 0.61 ;
      RECT  6.555 0.44 7.51 0.56 ;
      RECT  6.555 0.56 6.66 0.785 ;
      RECT  5.02 0.785 6.66 0.895 ;
      RECT  6.555 0.895 6.66 1.24 ;
      RECT  6.555 1.24 7.25 1.36 ;
      RECT  1.55 1.19 4.37 1.24 ;
      RECT  0.065 1.24 4.37 1.36 ;
      RECT  4.2 1.36 4.37 1.44 ;
      RECT  0.065 1.36 0.185 1.46 ;
      RECT  4.2 1.44 6.475 1.57 ;
      RECT  4.2 1.57 4.85 1.61 ;
  END
END SEN_AOI21B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI221_0P5
#      Description : "Two 2-input ANDs into 3-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI221_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI221_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0297 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0297 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0297 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0297 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.13 0.05 1.26 0.38 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.235 1.585 0.355 ;
      RECT  1.35 0.355 1.45 0.47 ;
      RECT  0.535 0.235 1.04 0.355 ;
      RECT  0.94 0.355 1.04 0.47 ;
      RECT  0.94 0.47 1.45 0.56 ;
      RECT  1.35 0.56 1.45 1.2 ;
      RECT  1.35 1.2 1.735 1.29 ;
      RECT  1.615 1.29 1.735 1.53 ;
    END
    ANTENNADIFFAREA 0.126 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.26 1.225 1.35 ;
      RECT  1.105 1.35 1.225 1.48 ;
      RECT  0.065 1.35 0.185 1.53 ;
      RECT  0.585 1.35 0.705 1.53 ;
      RECT  0.845 1.44 0.965 1.57 ;
      RECT  0.845 1.57 1.475 1.66 ;
      RECT  1.355 1.395 1.475 1.57 ;
  END
END SEN_AOI221_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI221_1
#      Description : "Two 2-input ANDs into 3-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI221_1
  CLASS CORE ;
  FOREIGN SEN_AOI221_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.41 0.445 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.195 0.05 1.365 0.235 ;
      RECT  0.065 0.05 0.185 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.56 0.24 1.1 0.325 ;
      RECT  0.56 0.325 1.735 0.36 ;
      RECT  1.615 0.2 1.735 0.325 ;
      RECT  1.01 0.36 1.735 0.42 ;
      RECT  1.35 0.42 1.45 1.3 ;
      RECT  1.35 1.3 1.735 1.39 ;
      RECT  1.615 1.39 1.735 1.52 ;
    END
    ANTENNADIFFAREA 0.269 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.21 1.225 1.32 ;
      RECT  1.105 1.32 1.225 1.39 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  0.79 1.48 1.5 1.6 ;
  END
END SEN_AOI221_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI221_2
#      Description : "Two 2-input ANDs into 3-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI221_2
  CLASS CORE ;
  FOREIGN SEN_AOI221_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.66 0.9 ;
      RECT  1.35 0.9 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.91 2.65 1.09 ;
      RECT  2.55 1.09 2.65 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.9 ;
      RECT  0.75 0.9 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.45 0.91 ;
      RECT  0.15 0.91 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.94 0.7 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.43 0.445 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.845 1.43 0.965 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.325 0.05 0.445 0.365 ;
      RECT  2.68 0.05 2.8 0.37 ;
      RECT  2.165 0.05 2.285 0.385 ;
      RECT  3.205 0.05 3.325 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.945 0.31 3.065 0.51 ;
      RECT  2.75 0.51 3.065 0.61 ;
      RECT  2.75 0.61 2.85 0.69 ;
      RECT  0.82 0.46 1.855 0.58 ;
      RECT  1.75 0.58 1.855 0.69 ;
      RECT  1.75 0.69 2.85 0.78 ;
      RECT  2.75 0.78 2.85 1.11 ;
      RECT  2.75 1.11 3.06 1.29 ;
    END
    ANTENNADIFFAREA 0.408 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.24 1.25 0.36 ;
      RECT  0.585 0.36 0.705 0.47 ;
      RECT  0.065 0.37 0.185 0.47 ;
      RECT  0.065 0.47 0.705 0.59 ;
      RECT  1.36 0.245 2.075 0.365 ;
      RECT  1.985 0.365 2.075 0.475 ;
      RECT  1.985 0.475 2.6 0.595 ;
      RECT  0.065 1.22 2.46 1.34 ;
      RECT  2.34 1.34 2.46 1.39 ;
      RECT  0.065 1.34 0.185 1.44 ;
      RECT  3.19 1.41 3.325 1.48 ;
      RECT  1.51 1.48 3.325 1.6 ;
  END
END SEN_AOI221_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI221_4
#      Description : "Two 2-input ANDs into 3-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI221_4
  CLASS CORE ;
  FOREIGN SEN_AOI221_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.9 ;
      RECT  2.95 0.9 3.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.91 4.85 1.09 ;
      RECT  4.75 1.09 4.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.85 0.89 ;
      RECT  5.75 0.89 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.845 1.44 0.965 1.75 ;
      RECT  1.55 1.44 1.67 1.75 ;
      RECT  2.07 1.44 2.19 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  3.545 0.05 3.715 0.305 ;
      RECT  4.08 0.05 4.25 0.305 ;
      RECT  0.3 0.05 0.47 0.375 ;
      RECT  0.82 0.05 0.99 0.375 ;
      RECT  5.2 0.05 5.32 0.395 ;
      RECT  4.655 0.05 4.775 0.56 ;
      RECT  5.74 0.05 5.86 0.595 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.94 0.485 5.63 0.6 ;
      RECT  4.94 0.6 5.06 0.655 ;
      RECT  1.24 0.225 2.45 0.345 ;
      RECT  2.33 0.345 2.45 0.47 ;
      RECT  2.33 0.47 3.25 0.575 ;
      RECT  2.33 0.575 3.515 0.59 ;
      RECT  3.15 0.59 3.515 0.655 ;
      RECT  3.15 0.655 5.06 0.765 ;
      RECT  4.94 0.765 5.06 1.11 ;
      RECT  4.94 1.11 5.65 1.29 ;
    END
    ANTENNADIFFAREA 0.845 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.56 0.23 3.455 0.36 ;
      RECT  3.365 0.36 3.455 0.395 ;
      RECT  3.365 0.395 4.545 0.485 ;
      RECT  0.065 0.36 0.19 0.47 ;
      RECT  0.065 0.47 2.22 0.58 ;
      RECT  0.065 1.23 4.59 1.35 ;
      RECT  0.065 1.35 0.185 1.45 ;
      RECT  5.73 1.34 5.85 1.44 ;
      RECT  2.54 1.44 5.85 1.56 ;
  END
END SEN_AOI221_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI222_1
#      Description : "Three 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|(C1&C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI222_1
  CLASS CORE ;
  FOREIGN SEN_AOI222_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.3 1.65 0.71 ;
      RECT  1.35 0.71 1.65 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.48 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.71 1.06 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.44 0.45 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.815 0.05 1.935 0.37 ;
      RECT  1.12 0.05 1.23 0.385 ;
      RECT  0.07 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.24 1.03 0.36 ;
      RECT  0.94 0.36 1.03 0.495 ;
      RECT  0.94 0.495 1.45 0.59 ;
      RECT  1.15 0.59 1.45 0.615 ;
      RECT  1.15 0.615 1.25 1.015 ;
      RECT  1.15 1.015 1.45 1.135 ;
      RECT  1.35 1.135 1.45 1.21 ;
      RECT  1.35 1.21 1.935 1.32 ;
      RECT  1.815 1.32 1.935 1.43 ;
    END
    ANTENNADIFFAREA 0.315 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.23 1.23 1.35 ;
      RECT  1.11 1.35 1.23 1.405 ;
      RECT  0.07 1.35 0.19 1.45 ;
      RECT  0.8 1.495 1.725 1.6 ;
  END
END SEN_AOI222_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI222_2
#      Description : "Three 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|(C1&C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI222_2
  CLASS CORE ;
  FOREIGN SEN_AOI222_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.7 3.65 0.89 ;
      RECT  3.55 0.89 3.65 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.32 0.71 2.45 0.83 ;
      RECT  2.02 0.83 2.45 0.93 ;
      RECT  2.35 0.93 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.83 1.65 1.09 ;
      RECT  1.35 1.09 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.99 0.87 ;
      RECT  0.75 0.87 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.42 0.445 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.845 1.425 0.965 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  1.555 0.05 1.675 0.36 ;
      RECT  3.345 0.05 3.465 0.38 ;
      RECT  0.325 0.05 0.445 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.025 0.49 2.97 0.595 ;
      RECT  2.55 0.595 2.97 0.61 ;
      RECT  2.025 0.595 2.115 0.65 ;
      RECT  2.55 0.61 2.65 1.01 ;
      RECT  0.815 0.47 1.18 0.59 ;
      RECT  1.09 0.59 1.18 0.65 ;
      RECT  1.09 0.65 2.115 0.74 ;
      RECT  2.55 1.01 2.85 1.1 ;
      RECT  2.75 1.1 2.85 1.27 ;
      RECT  2.75 1.27 3.46 1.39 ;
      RECT  3.345 1.1 3.46 1.27 ;
    END
    ANTENNADIFFAREA 0.498 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.215 1.28 0.335 ;
      RECT  0.585 0.335 0.705 0.475 ;
      RECT  0.065 0.36 0.185 0.475 ;
      RECT  0.065 0.475 0.705 0.58 ;
      RECT  1.815 0.23 2.455 0.35 ;
      RECT  2.335 0.35 2.455 0.4 ;
      RECT  1.815 0.35 1.935 0.45 ;
      RECT  1.27 0.45 1.935 0.56 ;
      RECT  2.565 0.23 3.21 0.35 ;
      RECT  2.565 0.35 2.685 0.4 ;
      RECT  3.08 0.35 3.21 0.47 ;
      RECT  3.08 0.47 3.725 0.59 ;
      RECT  3.605 0.37 3.725 0.47 ;
      RECT  0.065 1.21 1.26 1.33 ;
      RECT  0.065 1.33 0.185 1.43 ;
      RECT  1.145 1.33 1.26 1.48 ;
      RECT  1.145 1.48 2.45 1.6 ;
      RECT  2.335 1.43 2.45 1.48 ;
      RECT  1.555 1.22 2.66 1.34 ;
      RECT  1.555 1.34 1.675 1.39 ;
      RECT  2.54 1.34 2.66 1.48 ;
      RECT  2.54 1.48 3.725 1.61 ;
      RECT  3.605 1.41 3.725 1.48 ;
  END
END SEN_AOI222_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI222_4
#      Description : "Three 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|(C1&C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI222_4
  CLASS CORE ;
  FOREIGN SEN_AOI222_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.7 5.45 0.895 ;
      RECT  4.95 0.895 5.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.71 6.85 0.89 ;
      RECT  6.75 0.89 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.975 ;
      RECT  2.55 0.975 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.825 4.65 1.09 ;
      RECT  4.55 1.09 4.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 2.05 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.9 ;
      RECT  0.35 0.9 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.18 0.185 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.585 1.42 0.705 1.75 ;
      RECT  1.105 1.42 1.225 1.75 ;
      RECT  1.625 1.42 1.745 1.75 ;
      RECT  2.145 1.42 2.265 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  3.68 0.05 3.85 0.315 ;
      RECT  4.2 0.05 4.37 0.315 ;
      RECT  0.325 0.05 0.445 0.37 ;
      RECT  0.845 0.05 0.965 0.37 ;
      RECT  6.035 0.05 6.155 0.375 ;
      RECT  6.555 0.05 6.675 0.375 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.465 5.65 0.585 ;
      RECT  4.75 0.585 4.85 0.6 ;
      RECT  5.55 0.585 5.65 1.11 ;
      RECT  1.335 0.46 3.33 0.58 ;
      RECT  3.15 0.58 3.33 0.6 ;
      RECT  3.15 0.6 4.85 0.69 ;
      RECT  5.55 1.11 6.66 1.24 ;
      RECT  4.95 1.24 6.66 1.29 ;
      RECT  4.95 1.29 5.655 1.36 ;
    END
    ANTENNADIFFAREA 0.996 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.7 0.2 5.9 0.305 ;
      RECT  4.7 0.305 4.85 0.375 ;
      RECT  5.775 0.305 5.9 0.47 ;
      RECT  5.775 0.47 6.935 0.59 ;
      RECT  6.81 0.37 6.935 0.47 ;
      RECT  1.105 0.2 2.265 0.32 ;
      RECT  2.145 0.32 2.265 0.37 ;
      RECT  1.105 0.32 1.225 0.46 ;
      RECT  0.065 0.36 0.185 0.46 ;
      RECT  0.065 0.46 1.225 0.58 ;
      RECT  2.375 0.23 3.565 0.35 ;
      RECT  3.445 0.35 3.565 0.405 ;
      RECT  3.445 0.405 4.605 0.51 ;
      RECT  4.485 0.29 4.605 0.405 ;
      RECT  0.295 1.21 4.4 1.33 ;
      RECT  2.405 1.425 2.525 1.48 ;
      RECT  2.405 1.48 6.935 1.6 ;
      RECT  3.94 1.45 5.405 1.48 ;
      RECT  6.815 1.38 6.935 1.48 ;
  END
END SEN_AOI222_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI222_0P5
#      Description : "Three 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|(C1&C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI222_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI222_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.92 ;
      RECT  0.95 0.92 1.06 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.85 0.695 ;
      RECT  1.75 0.695 1.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.45 0.69 ;
      RECT  1.35 0.69 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.365 1.005 1.93 1.125 ;
      RECT  1.815 1.125 1.93 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.155 0.05 1.325 0.2 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.815 0.2 1.935 0.3 ;
      RECT  0.35 0.3 1.935 0.42 ;
      RECT  0.35 0.42 0.45 1.31 ;
      RECT  0.32 1.31 0.45 1.48 ;
    END
    ANTENNADIFFAREA 0.145 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.155 0.915 1.26 1.24 ;
      RECT  1.155 1.24 1.675 1.27 ;
      RECT  0.85 1.27 1.675 1.36 ;
      RECT  0.85 1.36 1.02 1.44 ;
      RECT  1.555 1.36 1.675 1.48 ;
      RECT  1.11 1.45 1.305 1.565 ;
      RECT  1.11 1.565 1.2 1.57 ;
      RECT  0.065 1.375 0.185 1.57 ;
      RECT  0.065 1.57 1.2 1.66 ;
      RECT  0.59 1.385 0.7 1.57 ;
  END
END SEN_AOI222_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI222_3
#      Description : "Three 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|(C1&C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI222_3
  CLASS CORE ;
  FOREIGN SEN_AOI222_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.171 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.171 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.171 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.171 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.171 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 5.05 0.89 ;
      RECT  4.95 0.89 5.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.171 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  3.46 1.44 3.59 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  3.96 1.47 4.13 1.75 ;
      RECT  4.48 1.47 4.65 1.75 ;
      RECT  5.02 1.41 5.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.65 0.05 2.82 0.24 ;
      RECT  3.19 0.05 3.36 0.24 ;
      RECT  0.56 0.05 0.73 0.41 ;
      RECT  4.48 0.05 4.65 0.43 ;
      RECT  5.02 0.05 5.145 0.47 ;
      RECT  0.06 0.05 0.19 0.525 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.625 0.18 2.22 0.28 ;
      RECT  2.12 0.28 2.22 0.33 ;
      RECT  1.625 0.28 1.745 0.49 ;
      RECT  2.12 0.33 4.16 0.42 ;
      RECT  1.07 0.49 1.745 0.58 ;
      RECT  1.07 0.58 1.65 0.605 ;
      RECT  1.55 0.605 1.65 1.26 ;
      RECT  0.275 1.26 1.65 1.375 ;
    END
    ANTENNADIFFAREA 0.696 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.295 1.535 0.4 ;
      RECT  0.845 0.4 0.96 0.5 ;
      RECT  0.325 0.38 0.445 0.5 ;
      RECT  0.325 0.5 0.96 0.6 ;
      RECT  1.885 0.39 2.005 0.51 ;
      RECT  1.885 0.51 3.115 0.615 ;
      RECT  3.655 0.52 4.94 0.62 ;
      RECT  1.835 1.24 4.935 1.35 ;
      RECT  0.065 1.37 0.185 1.465 ;
      RECT  0.065 1.465 3.37 1.59 ;
  END
END SEN_AOI222_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI222_8
#      Description : "Three 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2)|(C1&C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI222_8
  CLASS CORE ;
  FOREIGN SEN_AOI222_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.35 0.51 8.45 0.71 ;
      RECT  8.35 0.71 9.98 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4554 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.35 0.51 12.45 0.71 ;
      RECT  10.95 0.71 12.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4554 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 5.725 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4554 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.51 8.25 0.71 ;
      RECT  7.28 0.71 8.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4554 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.695 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4554 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.35 0.71 1.48 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4554 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  0.555 1.445 0.73 1.75 ;
      RECT  1.08 1.445 1.25 1.75 ;
      RECT  1.6 1.445 1.77 1.75 ;
      RECT  2.12 1.445 2.29 1.75 ;
      RECT  2.64 1.445 2.81 1.75 ;
      RECT  3.16 1.445 3.33 1.75 ;
      RECT  3.68 1.445 3.85 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  6.53 0.05 6.7 0.32 ;
      RECT  7.05 0.05 7.22 0.32 ;
      RECT  7.57 0.05 7.74 0.32 ;
      RECT  10.69 0.05 10.86 0.32 ;
      RECT  11.21 0.05 11.38 0.32 ;
      RECT  11.73 0.05 11.9 0.32 ;
      RECT  0.82 0.05 0.99 0.325 ;
      RECT  1.34 0.05 1.51 0.325 ;
      RECT  1.86 0.05 2.03 0.325 ;
      RECT  0.28 0.05 0.42 0.39 ;
      RECT  8.13 0.05 8.26 0.39 ;
      RECT  12.295 0.05 12.425 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.63 0.31 8.78 0.45 ;
      RECT  8.63 0.45 10.34 0.62 ;
      RECT  10.15 0.62 10.34 1.11 ;
      RECT  3.94 0.155 4.65 0.175 ;
      RECT  2.35 0.175 4.65 0.325 ;
      RECT  4.47 0.325 4.65 0.45 ;
      RECT  4.47 0.45 6.18 0.62 ;
      RECT  5.95 0.62 6.18 0.71 ;
      RECT  5.95 0.71 7.12 0.89 ;
      RECT  6.95 0.89 7.12 0.99 ;
      RECT  6.95 0.99 8.625 1.11 ;
      RECT  6.95 1.11 12.45 1.16 ;
      RECT  8.445 1.16 12.45 1.29 ;
    END
    ANTENNADIFFAREA 1.855 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.75 0.19 6.44 0.36 ;
      RECT  6.27 0.36 6.44 0.41 ;
      RECT  6.27 0.41 7.99 0.585 ;
      RECT  8.89 0.19 10.6 0.36 ;
      RECT  10.43 0.36 10.6 0.43 ;
      RECT  10.43 0.43 12.14 0.62 ;
      RECT  0.58 0.37 0.705 0.45 ;
      RECT  0.58 0.45 4.38 0.515 ;
      RECT  2.095 0.415 4.38 0.45 ;
      RECT  0.58 0.515 3.85 0.585 ;
      RECT  0.58 0.585 2.205 0.62 ;
      RECT  0.325 1.18 6.73 1.255 ;
      RECT  0.325 1.255 8.285 1.35 ;
      RECT  12.53 1.385 12.655 1.47 ;
      RECT  4.19 1.47 12.655 1.64 ;
  END
END SEN_AOI222_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_0P5
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI22_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.3 1.05 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.88 1.415 1.0 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.07 0.05 0.19 0.39 ;
      RECT  1.165 0.05 1.285 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.27 0.81 0.39 ;
      RECT  0.35 0.39 0.46 1.46 ;
    END
    ANTENNADIFFAREA 0.11 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.615 1.235 1.26 1.325 ;
      RECT  1.14 1.325 1.26 1.53 ;
      RECT  0.615 1.325 0.735 1.555 ;
      RECT  0.09 1.41 0.21 1.555 ;
      RECT  0.09 1.555 0.735 1.645 ;
  END
END SEN_AOI22_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_1
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_1
  CLASS CORE ;
  FOREIGN SEN_AOI22_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.925 ;
      RECT  0.75 0.925 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.88 1.415 1.0 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.17 0.05 1.29 0.39 ;
      RECT  0.08 0.05 0.2 0.57 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.24 0.81 0.36 ;
      RECT  0.35 0.36 0.45 1.29 ;
    END
    ANTENNADIFFAREA 0.224 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.61 1.21 1.25 1.31 ;
      RECT  0.61 1.31 0.73 1.41 ;
      RECT  1.14 1.31 1.25 1.43 ;
      RECT  0.085 1.41 0.73 1.525 ;
      RECT  0.085 1.525 0.205 1.63 ;
  END
END SEN_AOI22_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_2
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_2
  CLASS CORE ;
  FOREIGN SEN_AOI22_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.71 0.855 0.89 ;
      RECT  0.75 0.89 0.855 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.54 1.415 1.66 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  2.155 1.415 2.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.325 0.05 0.445 0.39 ;
      RECT  2.155 0.05 2.275 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.835 0.47 1.785 0.59 ;
      RECT  0.95 0.59 1.05 1.23 ;
      RECT  0.34 1.11 0.45 1.23 ;
      RECT  0.34 1.23 1.05 1.35 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.535 0.205 1.24 0.325 ;
      RECT  1.12 0.325 1.24 0.375 ;
      RECT  0.535 0.325 0.625 0.5 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 0.625 0.59 ;
      RECT  1.35 0.24 2.015 0.36 ;
      RECT  1.895 0.36 2.015 0.5 ;
      RECT  1.895 0.5 2.535 0.59 ;
      RECT  2.415 0.37 2.535 0.5 ;
      RECT  1.18 1.21 2.535 1.32 ;
      RECT  2.415 1.32 2.535 1.43 ;
      RECT  1.18 1.32 1.31 1.45 ;
      RECT  0.065 1.4 0.185 1.45 ;
      RECT  0.065 1.45 1.31 1.57 ;
  END
END SEN_AOI22_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_3
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_3
  CLASS CORE ;
  FOREIGN SEN_AOI22_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.925 ;
      RECT  1.55 0.925 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.9 ;
      RECT  0.35 0.9 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.45 0.9 ;
      RECT  1.95 0.9 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.9 1.415 2.02 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  2.42 1.43 2.54 1.75 ;
      RECT  2.94 1.43 3.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.6 0.05 0.72 0.37 ;
      RECT  2.68 0.05 2.8 0.375 ;
      RECT  3.215 0.05 3.335 0.575 ;
      RECT  0.08 0.05 0.2 0.58 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.12 0.44 2.305 0.56 ;
      RECT  1.12 0.56 1.25 0.61 ;
      RECT  1.15 0.61 1.25 1.24 ;
      RECT  0.31 1.24 1.53 1.36 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.86 0.225 1.525 0.345 ;
      RECT  0.86 0.345 0.98 0.46 ;
      RECT  0.315 0.46 0.98 0.58 ;
      RECT  1.875 0.225 2.54 0.345 ;
      RECT  2.42 0.345 2.54 0.47 ;
      RECT  2.42 0.47 3.085 0.59 ;
      RECT  1.64 1.21 3.32 1.3 ;
      RECT  3.2 1.3 3.32 1.42 ;
      RECT  1.64 1.3 1.76 1.455 ;
      RECT  0.08 1.35 0.2 1.455 ;
      RECT  0.08 1.455 1.76 1.575 ;
  END
END SEN_AOI22_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_4
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_4
  CLASS CORE ;
  FOREIGN SEN_AOI22_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.895 ;
      RECT  1.95 0.895 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.7 4.25 0.9 ;
      RECT  4.15 0.9 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.57 1.41 2.69 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  3.23 1.41 3.35 1.75 ;
      RECT  3.785 1.41 3.905 1.75 ;
      RECT  4.34 1.41 4.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.325 0.05 0.445 0.37 ;
      RECT  0.845 0.05 0.965 0.37 ;
      RECT  3.785 0.05 3.905 0.37 ;
      RECT  4.34 0.05 4.46 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.34 0.47 3.395 0.59 ;
      RECT  1.34 0.59 1.45 1.215 ;
      RECT  0.295 1.215 2.06 1.335 ;
    END
    ANTENNADIFFAREA 0.872 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.24 2.29 0.36 ;
      RECT  1.105 0.36 1.225 0.46 ;
      RECT  0.065 0.36 0.185 0.46 ;
      RECT  0.065 0.46 1.225 0.58 ;
      RECT  2.42 0.24 3.62 0.36 ;
      RECT  3.5 0.36 3.62 0.47 ;
      RECT  3.5 0.47 4.735 0.59 ;
      RECT  4.615 0.37 4.735 0.47 ;
      RECT  2.19 1.21 4.735 1.32 ;
      RECT  4.615 1.32 4.735 1.43 ;
      RECT  2.19 1.32 2.31 1.44 ;
      RECT  0.065 1.34 0.185 1.44 ;
      RECT  0.065 1.44 2.31 1.56 ;
  END
END SEN_AOI22_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_12
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_12
  CLASS CORE ;
  FOREIGN SEN_AOI22_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.215 0.51 12.375 0.925 ;
      RECT  10.755 0.51 11.055 0.69 ;
      RECT  10.965 0.69 11.055 0.925 ;
      RECT  9.77 0.51 10.07 0.69 ;
      RECT  9.97 0.69 10.07 0.935 ;
      RECT  8.81 0.51 9.11 0.69 ;
      RECT  9.02 0.69 9.11 0.925 ;
      RECT  7.08 0.51 8.15 0.6 ;
      RECT  7.85 0.6 8.15 0.69 ;
      RECT  7.08 0.6 7.25 0.925 ;
      RECT  8.055 0.69 8.15 0.925 ;
      LAYER M2 ;
      RECT  7.81 0.55 12.36 0.65 ;
      LAYER V1 ;
      RECT  12.215 0.55 12.315 0.65 ;
      RECT  10.755 0.55 10.855 0.65 ;
      RECT  10.955 0.55 11.055 0.65 ;
      RECT  9.77 0.55 9.87 0.65 ;
      RECT  9.97 0.55 10.07 0.65 ;
      RECT  8.81 0.55 8.91 0.65 ;
      RECT  9.01 0.55 9.11 0.65 ;
      RECT  7.85 0.55 7.95 0.65 ;
      RECT  8.05 0.55 8.15 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.55 0.51 12.65 1.09 ;
      RECT  11.615 0.71 11.945 0.9 ;
      RECT  10.365 0.71 10.665 0.9 ;
      RECT  9.38 0.71 9.68 0.9 ;
      RECT  8.42 0.71 8.72 0.9 ;
      RECT  7.46 0.71 7.76 0.9 ;
      RECT  6.35 0.71 6.49 1.09 ;
      LAYER M2 ;
      RECT  6.345 0.75 12.69 0.85 ;
      LAYER V1 ;
      RECT  12.55 0.75 12.65 0.85 ;
      RECT  11.645 0.75 11.745 0.85 ;
      RECT  11.845 0.75 11.945 0.85 ;
      RECT  10.365 0.75 10.465 0.85 ;
      RECT  10.565 0.75 10.665 0.85 ;
      RECT  9.38 0.75 9.48 0.85 ;
      RECT  9.58 0.75 9.68 0.85 ;
      RECT  8.42 0.75 8.52 0.85 ;
      RECT  8.62 0.75 8.72 0.85 ;
      RECT  7.46 0.75 7.56 0.85 ;
      RECT  7.66 0.75 7.76 0.85 ;
      RECT  6.385 0.75 6.485 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.71 6.05 0.9 ;
      RECT  4.79 0.71 5.165 0.9 ;
      RECT  3.755 0.71 4.125 0.9 ;
      RECT  2.74 0.71 3.085 0.9 ;
      RECT  1.625 0.71 2.045 0.9 ;
      RECT  0.455 0.71 1.14 0.9 ;
      LAYER M2 ;
      RECT  0.795 0.75 6.09 0.85 ;
      LAYER V1 ;
      RECT  5.75 0.75 5.85 0.85 ;
      RECT  5.95 0.75 6.05 0.85 ;
      RECT  4.865 0.75 4.965 0.85 ;
      RECT  5.065 0.75 5.165 0.85 ;
      RECT  3.825 0.75 3.925 0.85 ;
      RECT  4.025 0.75 4.125 0.85 ;
      RECT  2.785 0.75 2.885 0.85 ;
      RECT  2.985 0.75 3.085 0.85 ;
      RECT  1.745 0.75 1.845 0.85 ;
      RECT  1.945 0.75 2.045 0.85 ;
      RECT  0.835 0.75 0.935 0.85 ;
      RECT  1.035 0.75 1.135 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.305 0.755 5.45 0.91 ;
      RECT  5.305 0.91 5.65 0.99 ;
      RECT  3.275 0.755 3.365 0.91 ;
      RECT  3.275 0.91 3.65 0.99 ;
      RECT  2.15 0.755 2.385 0.91 ;
      RECT  2.15 0.91 2.65 0.99 ;
      RECT  1.23 0.755 1.45 0.99 ;
      RECT  1.23 0.99 6.255 1.0 ;
      RECT  4.345 0.735 4.65 0.99 ;
      RECT  6.15 0.71 6.255 0.99 ;
      RECT  0.15 0.71 0.25 1.0 ;
      RECT  0.15 1.0 6.255 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.45 0.475 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  0.82 1.45 0.99 1.75 ;
      RECT  1.34 1.45 1.51 1.75 ;
      RECT  1.86 1.45 2.03 1.75 ;
      RECT  2.38 1.45 2.55 1.75 ;
      RECT  2.9 1.45 3.07 1.75 ;
      RECT  3.42 1.45 3.59 1.75 ;
      RECT  3.94 1.45 4.11 1.75 ;
      RECT  4.46 1.45 4.63 1.75 ;
      RECT  4.98 1.45 5.15 1.75 ;
      RECT  5.5 1.45 5.67 1.75 ;
      RECT  6.045 1.44 6.15 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  1.08 0.05 1.25 0.305 ;
      RECT  2.12 0.05 2.29 0.305 ;
      RECT  3.16 0.05 3.33 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  5.24 0.05 5.41 0.305 ;
      RECT  6.28 0.05 6.45 0.305 ;
      RECT  7.39 0.05 7.56 0.32 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  12.61 0.05 12.74 0.39 ;
      RECT  8.455 0.05 8.575 0.62 ;
      RECT  9.495 0.05 9.615 0.62 ;
      RECT  10.535 0.05 10.655 0.62 ;
      RECT  11.575 0.05 11.69 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  12.035 0.275 12.265 0.395 ;
      RECT  12.035 0.395 12.125 1.03 ;
      RECT  11.0 0.3 11.25 0.42 ;
      RECT  11.145 0.42 11.25 1.03 ;
      RECT  10.03 0.25 10.25 0.42 ;
      RECT  10.16 0.42 10.25 1.03 ;
      RECT  8.915 0.24 9.29 0.36 ;
      RECT  9.2 0.36 9.29 1.03 ;
      RECT  7.88 0.25 8.33 0.37 ;
      RECT  8.24 0.37 8.33 1.03 ;
      RECT  6.75 0.19 7.0 0.31 ;
      RECT  6.55 0.31 7.0 0.36 ;
      RECT  6.55 0.36 6.89 0.415 ;
      RECT  3.55 0.31 3.85 0.415 ;
      RECT  0.53 0.415 6.89 0.585 ;
      RECT  4.665 0.305 4.97 0.415 ;
      RECT  6.64 0.585 6.89 1.03 ;
      RECT  6.64 1.03 12.46 1.29 ;
      LAYER M2 ;
      RECT  3.51 0.35 6.89 0.45 ;
      LAYER V1 ;
      RECT  3.55 0.35 3.65 0.45 ;
      RECT  3.75 0.35 3.85 0.45 ;
      RECT  4.665 0.35 4.765 0.45 ;
      RECT  4.865 0.35 4.965 0.45 ;
      RECT  6.55 0.35 6.65 0.45 ;
      RECT  6.75 0.35 6.85 0.45 ;
    END
    ANTENNADIFFAREA 2.634 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 1.18 6.49 1.35 ;
      RECT  6.24 1.35 6.49 1.415 ;
      RECT  3.71 1.35 3.81 1.49 ;
      RECT  4.24 1.35 4.34 1.49 ;
      RECT  6.24 1.415 12.72 1.64 ;
      LAYER M2 ;
      RECT  3.67 1.35 6.385 1.45 ;
      LAYER V1 ;
      RECT  3.71 1.35 3.81 1.45 ;
      RECT  4.24 1.35 4.34 1.45 ;
      RECT  6.245 1.35 6.345 1.45 ;
  END
END SEN_AOI22_12
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_6
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_6
  CLASS CORE ;
  FOREIGN SEN_AOI22_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.565 0.51 5.865 0.69 ;
      RECT  5.775 0.69 5.865 0.935 ;
      RECT  4.605 0.51 4.905 0.69 ;
      RECT  4.645 0.69 4.785 0.925 ;
      RECT  3.795 0.51 4.125 0.69 ;
      RECT  3.795 0.69 3.885 0.925 ;
      LAYER M2 ;
      RECT  3.785 0.55 5.905 0.65 ;
      LAYER V1 ;
      RECT  5.565 0.55 5.665 0.65 ;
      RECT  5.765 0.55 5.865 0.65 ;
      RECT  4.605 0.55 4.705 0.65 ;
      RECT  4.805 0.55 4.905 0.65 ;
      RECT  3.825 0.55 3.925 0.65 ;
      RECT  4.025 0.55 4.125 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.51 6.34 0.925 ;
      RECT  5.235 0.71 5.42 1.0 ;
      RECT  4.215 0.71 4.515 0.9 ;
      RECT  3.26 0.71 3.42 0.995 ;
      LAYER M2 ;
      RECT  3.26 0.75 6.29 0.85 ;
      LAYER V1 ;
      RECT  6.15 0.75 6.25 0.85 ;
      RECT  5.235 0.75 5.335 0.85 ;
      RECT  4.215 0.75 4.315 0.85 ;
      RECT  4.415 0.75 4.515 0.85 ;
      RECT  3.3 0.75 3.4 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.9 ;
      RECT  1.6 0.71 1.955 0.9 ;
      RECT  0.63 0.71 1.135 0.9 ;
      LAYER M2 ;
      RECT  0.795 0.75 2.89 0.85 ;
      LAYER V1 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.655 0.75 1.755 0.85 ;
      RECT  1.855 0.75 1.955 0.85 ;
      RECT  0.835 0.75 0.935 0.85 ;
      RECT  1.035 0.75 1.135 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.035 0.755 3.145 0.91 ;
      RECT  2.95 0.91 3.145 1.02 ;
      RECT  2.265 0.755 2.45 0.91 ;
      RECT  2.15 0.91 2.45 1.02 ;
      RECT  1.225 0.75 1.315 0.91 ;
      RECT  1.225 0.91 1.45 1.02 ;
      RECT  0.15 0.71 0.275 0.91 ;
      RECT  0.15 0.91 0.45 1.02 ;
      RECT  0.15 1.02 3.145 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.82 1.48 0.99 1.75 ;
      RECT  1.34 1.48 1.51 1.75 ;
      RECT  1.86 1.48 2.03 1.75 ;
      RECT  2.38 1.48 2.55 1.75 ;
      RECT  2.9 1.48 3.07 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.08 0.05 1.25 0.32 ;
      RECT  2.12 0.05 2.29 0.32 ;
      RECT  3.16 0.05 3.33 0.32 ;
      RECT  5.25 0.05 5.4 0.36 ;
      RECT  0.06 0.05 0.19 0.385 ;
      RECT  4.21 0.05 4.36 0.385 ;
      RECT  6.325 0.05 6.455 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.8 0.25 6.05 0.42 ;
      RECT  5.96 0.42 6.05 1.11 ;
      RECT  4.72 0.23 5.11 0.355 ;
      RECT  5.015 0.355 5.11 0.91 ;
      RECT  4.95 0.91 5.11 1.11 ;
      RECT  3.55 0.25 3.81 0.42 ;
      RECT  3.55 0.42 3.68 0.435 ;
      RECT  0.53 0.435 3.68 0.565 ;
      RECT  3.55 0.565 3.68 1.11 ;
      RECT  3.445 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.215 3.315 1.345 ;
      RECT  3.17 1.345 3.315 1.415 ;
      RECT  0.065 1.345 0.185 1.44 ;
      RECT  3.17 1.415 6.45 1.545 ;
  END
END SEN_AOI22_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_8
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_8
  CLASS CORE ;
  FOREIGN SEN_AOI22_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.51 8.06 0.94 ;
      RECT  6.655 0.51 6.825 0.69 ;
      RECT  6.735 0.69 6.825 0.925 ;
      RECT  5.535 0.51 5.835 0.69 ;
      RECT  5.745 0.69 5.835 0.925 ;
      RECT  4.88 0.51 5.02 0.94 ;
      LAYER M2 ;
      RECT  4.88 0.55 8.09 0.65 ;
      LAYER V1 ;
      RECT  7.95 0.55 8.05 0.65 ;
      RECT  6.725 0.55 6.825 0.65 ;
      RECT  5.535 0.55 5.635 0.65 ;
      RECT  5.735 0.55 5.835 0.65 ;
      RECT  4.92 0.55 5.02 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.71 8.39 0.935 ;
      RECT  7.215 0.71 7.645 0.9 ;
      RECT  6.14 0.71 6.45 0.9 ;
      RECT  5.145 0.71 5.445 0.9 ;
      RECT  4.27 0.71 4.45 0.93 ;
      RECT  4.27 0.93 4.37 1.08 ;
      LAYER M2 ;
      RECT  4.31 0.75 8.29 0.85 ;
      LAYER V1 ;
      RECT  8.15 0.75 8.25 0.85 ;
      RECT  7.33 0.75 7.43 0.85 ;
      RECT  7.53 0.75 7.63 0.85 ;
      RECT  6.15 0.75 6.25 0.85 ;
      RECT  6.35 0.75 6.45 0.85 ;
      RECT  5.145 0.75 5.245 0.85 ;
      RECT  5.345 0.75 5.445 0.85 ;
      RECT  4.35 0.75 4.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.695 0.71 3.995 0.9 ;
      RECT  2.71 0.71 3.085 0.9 ;
      RECT  1.67 0.71 2.045 0.9 ;
      RECT  0.635 0.71 1.135 0.9 ;
      LAYER M2 ;
      RECT  0.795 0.75 4.09 0.85 ;
      LAYER V1 ;
      RECT  3.695 0.75 3.795 0.85 ;
      RECT  3.895 0.75 3.995 0.85 ;
      RECT  2.785 0.75 2.885 0.85 ;
      RECT  2.985 0.75 3.085 0.85 ;
      RECT  1.745 0.75 1.845 0.85 ;
      RECT  1.945 0.75 2.045 0.85 ;
      RECT  0.835 0.75 0.935 0.85 ;
      RECT  1.035 0.75 1.135 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.265 0.75 2.355 0.91 ;
      RECT  2.15 0.91 2.355 1.025 ;
      RECT  1.225 0.75 1.315 0.91 ;
      RECT  1.225 0.91 1.45 1.025 ;
      RECT  0.15 0.71 0.275 0.91 ;
      RECT  0.15 0.91 0.45 1.025 ;
      RECT  0.15 1.025 4.175 1.115 ;
      RECT  3.265 0.73 3.45 1.025 ;
      RECT  4.085 0.75 4.175 1.025 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.82 1.48 0.99 1.75 ;
      RECT  1.34 1.48 1.51 1.75 ;
      RECT  1.86 1.48 2.03 1.75 ;
      RECT  2.38 1.48 2.55 1.75 ;
      RECT  2.9 1.48 3.07 1.75 ;
      RECT  3.42 1.48 3.59 1.75 ;
      RECT  3.94 1.48 4.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  1.08 0.05 1.25 0.32 ;
      RECT  2.12 0.05 2.29 0.32 ;
      RECT  3.16 0.05 3.33 0.32 ;
      RECT  4.2 0.05 4.37 0.32 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  8.4 0.05 8.52 0.59 ;
      RECT  5.25 0.05 5.41 0.62 ;
      RECT  6.29 0.05 6.435 0.62 ;
      RECT  7.33 0.05 7.48 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.215 8.035 0.335 ;
      RECT  7.75 0.335 7.86 1.11 ;
      RECT  6.775 0.24 7.05 0.36 ;
      RECT  6.915 0.36 7.05 1.11 ;
      RECT  5.73 0.24 6.05 0.36 ;
      RECT  5.925 0.36 6.05 1.11 ;
      RECT  4.63 0.265 4.935 0.385 ;
      RECT  4.63 0.385 4.75 0.45 ;
      RECT  0.555 0.45 4.75 0.62 ;
      RECT  4.55 0.62 4.75 1.11 ;
      RECT  4.55 1.11 8.25 1.12 ;
      RECT  4.5 1.12 8.25 1.29 ;
    END
    ANTENNADIFFAREA 1.752 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 1.215 4.38 1.385 ;
      RECT  4.2 1.385 4.38 1.415 ;
      RECT  4.2 1.415 8.49 1.585 ;
  END
END SEN_AOI22_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_S_1
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_S_1
  CLASS CORE ;
  FOREIGN SEN_AOI22_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.41 0.455 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  1.145 0.05 1.275 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.265 1.05 0.385 ;
      RECT  0.95 0.385 1.05 1.18 ;
      RECT  0.805 1.18 1.05 1.3 ;
    END
    ANTENNADIFFAREA 0.174 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.21 0.71 1.3 ;
      RECT  0.59 1.3 0.71 1.4 ;
      RECT  0.07 1.3 0.19 1.43 ;
      RECT  0.59 1.4 1.285 1.52 ;
  END
END SEN_AOI22_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_S_1P5
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_S_1P5
  CLASS CORE ;
  FOREIGN SEN_AOI22_S_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.615 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0783 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0783 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0783 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.91 ;
      RECT  1.55 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0783 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.46 1.39 1.58 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  2.025 1.405 2.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  2.025 0.05 2.145 0.4 ;
      RECT  0.06 0.05 0.185 0.58 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.14 1.485 0.2 ;
      RECT  0.54 0.2 1.655 0.23 ;
      RECT  1.395 0.23 1.655 0.32 ;
      RECT  0.54 0.23 0.65 1.205 ;
      RECT  0.275 1.205 1.015 1.325 ;
    END
    ANTENNADIFFAREA 0.303 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.76 0.32 1.305 0.42 ;
      RECT  1.215 0.42 1.305 0.435 ;
      RECT  1.215 0.435 1.885 0.525 ;
      RECT  1.765 0.19 1.885 0.435 ;
      RECT  1.2 1.18 1.935 1.3 ;
      RECT  1.2 1.3 1.31 1.415 ;
      RECT  0.065 1.415 1.31 1.535 ;
      RECT  0.065 1.535 0.185 1.64 ;
  END
END SEN_AOI22_S_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_S_2
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_S_2
  CLASS CORE ;
  FOREIGN SEN_AOI22_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.695 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.585 1.41 0.715 1.75 ;
      RECT  1.105 1.41 1.235 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.325 0.05 0.455 0.39 ;
      RECT  2.135 0.05 2.265 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.85 0.33 0.97 0.47 ;
      RECT  0.85 0.47 1.74 0.56 ;
      RECT  1.62 0.33 1.74 0.47 ;
      RECT  1.35 0.56 1.45 0.99 ;
      RECT  1.35 0.99 1.85 1.105 ;
      RECT  1.75 1.105 1.85 1.185 ;
      RECT  1.75 1.185 2.31 1.305 ;
    END
    ANTENNADIFFAREA 0.348 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.59 0.15 1.23 0.24 ;
      RECT  1.11 0.24 1.23 0.38 ;
      RECT  0.59 0.24 0.71 0.48 ;
      RECT  0.07 0.245 0.19 0.48 ;
      RECT  0.07 0.48 0.71 0.57 ;
      RECT  1.36 0.15 2.0 0.24 ;
      RECT  1.36 0.24 1.48 0.38 ;
      RECT  1.88 0.24 2.0 0.48 ;
      RECT  1.88 0.48 2.52 0.57 ;
      RECT  2.4 0.24 2.52 0.48 ;
      RECT  0.28 1.195 1.48 1.315 ;
      RECT  1.36 1.315 1.48 1.44 ;
      RECT  1.36 1.44 2.52 1.56 ;
      RECT  2.4 1.34 2.52 1.44 ;
  END
END SEN_AOI22_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_S_4
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_S_4
  CLASS CORE ;
  FOREIGN SEN_AOI22_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.71 ;
      RECT  1.35 0.71 1.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.4 1.41 2.53 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  2.92 1.41 3.05 1.75 ;
      RECT  3.44 1.41 3.57 1.75 ;
      RECT  3.96 1.41 4.09 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  3.445 0.05 3.565 0.39 ;
      RECT  4.04 0.05 4.16 0.585 ;
      RECT  0.24 0.05 0.36 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.575 0.435 2.845 0.555 ;
      RECT  1.95 0.555 2.05 1.11 ;
      RECT  0.34 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.702 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.085 0.215 2.06 0.335 ;
      RECT  1.085 0.335 1.195 0.48 ;
      RECT  0.585 0.34 0.705 0.48 ;
      RECT  0.585 0.48 1.195 0.59 ;
      RECT  2.36 0.215 3.25 0.335 ;
      RECT  3.155 0.335 3.25 0.48 ;
      RECT  3.155 0.48 3.825 0.59 ;
      RECT  3.705 0.34 3.825 0.48 ;
      RECT  2.145 1.19 4.345 1.31 ;
      RECT  2.145 1.31 2.265 1.44 ;
      RECT  4.225 1.31 4.345 1.63 ;
      RECT  0.065 1.34 0.185 1.44 ;
      RECT  0.065 1.44 2.265 1.56 ;
  END
END SEN_AOI22_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_S_8
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_S_8
  CLASS CORE ;
  FOREIGN SEN_AOI22_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.465 0.89 ;
      RECT  3.35 0.89 3.465 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 1.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 5.25 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.51 8.05 0.71 ;
      RECT  6.55 0.71 8.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.225 1.44 4.355 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  4.745 1.44 4.875 1.75 ;
      RECT  5.265 1.44 5.395 1.75 ;
      RECT  5.79 1.25 5.91 1.75 ;
      RECT  6.31 1.25 6.43 1.75 ;
      RECT  6.83 1.25 6.95 1.75 ;
      RECT  7.35 1.25 7.47 1.75 ;
      RECT  7.89 1.21 8.01 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  0.765 0.05 0.895 0.355 ;
      RECT  1.285 0.05 1.415 0.355 ;
      RECT  1.795 0.05 1.965 0.355 ;
      RECT  6.28 0.05 6.41 0.36 ;
      RECT  6.825 0.05 6.955 0.36 ;
      RECT  7.345 0.05 7.475 0.36 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  7.895 0.05 8.025 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.385 0.415 5.675 0.585 ;
      RECT  3.68 0.585 3.85 1.18 ;
      RECT  0.07 1.11 3.25 1.18 ;
      RECT  0.07 1.18 3.85 1.29 ;
      RECT  3.115 1.29 3.85 1.35 ;
    END
    ANTENNADIFFAREA 1.446 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.08 0.155 3.855 0.325 ;
      RECT  2.08 0.325 2.25 0.445 ;
      RECT  0.375 0.445 2.25 0.615 ;
      RECT  4.205 0.155 5.94 0.325 ;
      RECT  5.77 0.325 5.94 0.45 ;
      RECT  5.77 0.45 7.78 0.62 ;
      RECT  5.385 0.98 7.73 1.15 ;
      RECT  5.385 1.15 5.555 1.18 ;
      RECT  3.95 1.18 5.555 1.35 ;
      RECT  3.95 1.35 4.115 1.45 ;
      RECT  0.3 1.45 4.115 1.62 ;
  END
END SEN_AOI22_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_0P75
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_0P75
  CLASS CORE ;
  FOREIGN SEN_AOI22_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.505 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.865 1.415 1.0 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.075 0.05 0.205 0.39 ;
      RECT  1.15 0.05 1.28 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.24 0.785 0.355 ;
      RECT  0.35 0.355 0.45 1.385 ;
    END
    ANTENNADIFFAREA 0.166 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.605 1.215 1.255 1.305 ;
      RECT  1.135 1.305 1.255 1.435 ;
      RECT  0.605 1.305 0.73 1.52 ;
      RECT  0.08 1.37 0.2 1.52 ;
      RECT  0.08 1.52 0.73 1.61 ;
  END
END SEN_AOI22_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_5
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_5
  CLASS CORE ;
  FOREIGN SEN_AOI22_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.85 0.9 ;
      RECT  2.75 0.9 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.05 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.055 0.71 3.85 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 5.25 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.915 1.435 3.05 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  3.435 1.435 3.575 1.75 ;
      RECT  3.955 1.435 4.085 1.75 ;
      RECT  4.475 1.435 4.61 1.75 ;
      RECT  4.995 1.435 5.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  4.22 0.05 4.35 0.36 ;
      RECT  4.74 0.05 4.87 0.36 ;
      RECT  0.58 0.05 0.71 0.395 ;
      RECT  1.1 0.05 1.23 0.4 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.3 0.05 5.42 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.575 0.48 3.85 0.595 ;
      RECT  1.74 0.595 1.85 1.11 ;
      RECT  0.34 1.11 2.53 1.29 ;
    END
    ANTENNADIFFAREA 1.08 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.365 0.24 2.58 0.36 ;
      RECT  1.365 0.36 1.485 0.5 ;
      RECT  0.33 0.4 0.44 0.5 ;
      RECT  0.33 0.5 1.485 0.62 ;
      RECT  2.865 0.24 4.09 0.36 ;
      RECT  3.96 0.36 4.09 0.48 ;
      RECT  3.96 0.48 5.16 0.595 ;
      RECT  2.66 1.225 5.435 1.335 ;
      RECT  2.66 1.335 2.79 1.445 ;
      RECT  0.065 1.33 0.185 1.445 ;
      RECT  0.065 1.445 2.79 1.555 ;
  END
END SEN_AOI22_5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_T_0P5
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_T_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI22_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.65 0.69 ;
      RECT  0.55 0.69 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.4 0.445 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.065 0.05 0.19 0.39 ;
      RECT  1.14 0.05 1.27 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.535 0.215 1.05 0.335 ;
      RECT  0.94 0.335 1.05 1.305 ;
      RECT  0.82 1.305 1.05 1.405 ;
    END
    ANTENNADIFFAREA 0.108 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 1.22 0.705 1.31 ;
      RECT  0.065 1.31 0.185 1.44 ;
      RECT  0.585 1.31 0.705 1.495 ;
      RECT  0.585 1.495 1.28 1.6 ;
  END
END SEN_AOI22_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_T_1
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_T_1
  CLASS CORE ;
  FOREIGN SEN_AOI22_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.505 1.05 0.71 ;
      RECT  0.95 0.71 1.45 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.9 ;
      RECT  1.75 0.9 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.445 0.85 0.985 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.495 0.47 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.82 1.495 0.99 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.295 0.05 0.425 0.39 ;
      RECT  1.54 0.05 1.67 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.24 1.11 0.345 ;
      RECT  0.55 0.345 0.65 1.085 ;
      RECT  0.55 1.085 1.54 1.205 ;
    END
    ANTENNADIFFAREA 0.302 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.285 0.36 1.405 0.49 ;
      RECT  1.285 0.49 1.925 0.58 ;
      RECT  1.805 0.36 1.925 0.49 ;
      RECT  0.06 1.295 1.745 1.405 ;
      RECT  0.06 1.405 0.185 1.515 ;
      RECT  1.625 1.405 1.745 1.52 ;
  END
END SEN_AOI22_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_T_1P5
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_T_1P5
  CLASS CORE ;
  FOREIGN SEN_AOI22_T_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.655 0.91 ;
      RECT  1.55 0.91 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.745 0.51 2.85 0.71 ;
      RECT  2.35 0.71 2.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1398 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1506 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1506 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.42 0.45 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.84 1.42 0.97 1.75 ;
      RECT  1.36 1.42 1.49 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  2.14 0.05 2.27 0.39 ;
      RECT  2.695 0.05 2.825 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.795 0.45 1.85 0.545 ;
      RECT  1.75 0.545 1.85 0.71 ;
      RECT  1.75 0.71 2.25 0.8 ;
      RECT  2.15 0.8 2.25 1.11 ;
      RECT  2.15 1.11 2.65 1.185 ;
      RECT  1.845 1.185 2.65 1.29 ;
    END
    ANTENNADIFFAREA 0.324 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.19 1.225 0.28 ;
      RECT  1.105 0.28 1.225 0.36 ;
      RECT  0.585 0.28 0.705 0.45 ;
      RECT  0.065 0.32 0.185 0.45 ;
      RECT  0.065 0.45 0.705 0.54 ;
      RECT  1.315 0.215 2.05 0.335 ;
      RECT  1.95 0.335 2.05 0.48 ;
      RECT  1.95 0.48 2.58 0.59 ;
      RECT  0.065 1.205 1.745 1.325 ;
      RECT  0.065 1.325 0.19 1.43 ;
      RECT  1.625 1.325 1.745 1.45 ;
      RECT  1.625 1.45 2.855 1.57 ;
  END
END SEN_AOI22_T_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_T_2
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_T_2
  CLASS CORE ;
  FOREIGN SEN_AOI22_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1872 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.58 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 0.71 ;
      RECT  1.15 0.71 1.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.305 1.455 0.475 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.825 1.455 0.995 1.75 ;
      RECT  1.415 1.455 1.585 1.75 ;
      RECT  2.065 1.455 2.235 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  2.185 0.05 2.355 0.305 ;
      RECT  2.705 0.05 2.875 0.305 ;
      RECT  1.095 0.05 1.265 0.32 ;
      RECT  1.67 0.05 1.79 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.225 0.46 3.45 0.56 ;
      RECT  3.35 0.56 3.45 1.21 ;
      RECT  0.085 0.315 0.175 0.41 ;
      RECT  0.085 0.41 0.77 0.51 ;
      RECT  0.67 0.51 0.77 0.685 ;
      RECT  0.67 0.685 0.85 0.785 ;
      RECT  0.75 0.785 0.85 1.06 ;
      RECT  0.75 1.06 2.85 1.16 ;
      RECT  2.75 1.16 2.85 1.21 ;
      RECT  2.75 1.21 3.45 1.315 ;
    END
    ANTENNADIFFAREA 0.451 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.305 0.215 0.97 0.305 ;
      RECT  0.86 0.305 0.97 0.41 ;
      RECT  0.86 0.41 1.57 0.515 ;
      RECT  3.0 0.21 3.62 0.305 ;
      RECT  3.52 0.305 3.62 0.385 ;
      RECT  3.0 0.305 3.1 0.42 ;
      RECT  1.96 0.29 2.06 0.42 ;
      RECT  1.96 0.42 3.1 0.53 ;
      RECT  0.08 1.25 2.53 1.35 ;
      RECT  2.42 1.35 2.53 1.415 ;
      RECT  0.08 1.35 0.18 1.49 ;
      RECT  2.42 1.415 3.68 1.525 ;
  END
END SEN_AOI22_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_T_3
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_T_3
  CLASS CORE ;
  FOREIGN SEN_AOI22_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.74 0.71 5.05 0.94 ;
      RECT  4.95 0.94 5.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.835 ;
      RECT  1.75 0.835 2.735 0.89 ;
      RECT  2.12 0.89 2.735 0.935 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3024 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3024 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.455 0.47 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.82 1.455 0.99 1.75 ;
      RECT  1.34 1.455 1.51 1.75 ;
      RECT  1.86 1.455 2.03 1.75 ;
      RECT  2.38 1.455 2.55 1.75 ;
      RECT  2.9 1.455 3.07 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.9 0.05 3.07 0.305 ;
      RECT  3.42 0.05 3.59 0.305 ;
      RECT  3.94 0.05 4.11 0.305 ;
      RECT  2.38 0.05 2.55 0.32 ;
      RECT  0.3 0.05 0.47 0.355 ;
      RECT  0.82 0.05 0.99 0.355 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.01 0.335 5.13 0.445 ;
      RECT  4.43 0.445 5.13 0.56 ;
      RECT  4.55 0.56 4.65 1.21 ;
      RECT  1.315 0.43 2.525 0.54 ;
      RECT  2.425 0.54 2.525 0.63 ;
      RECT  2.425 0.63 3.25 0.73 ;
      RECT  3.15 0.73 3.25 1.02 ;
      RECT  3.15 1.02 3.56 1.12 ;
      RECT  3.45 1.12 3.56 1.21 ;
      RECT  3.45 1.21 4.92 1.325 ;
    END
    ANTENNADIFFAREA 0.835 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.11 0.23 2.29 0.34 ;
      RECT  1.11 0.34 1.22 0.445 ;
      RECT  0.07 0.335 0.18 0.445 ;
      RECT  0.07 0.445 1.22 0.555 ;
      RECT  4.235 0.245 4.92 0.355 ;
      RECT  4.235 0.355 4.335 0.42 ;
      RECT  2.615 0.42 4.335 0.53 ;
      RECT  0.065 1.24 3.3 1.35 ;
      RECT  3.19 1.35 3.3 1.44 ;
      RECT  0.065 1.35 0.19 1.465 ;
      RECT  3.19 1.44 5.13 1.56 ;
      RECT  5.01 1.325 5.13 1.44 ;
  END
END SEN_AOI22_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_T_4
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_T_4
  CLASS CORE ;
  FOREIGN SEN_AOI22_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.3 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.71 6.65 0.91 ;
      RECT  5.15 0.91 6.65 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.675 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.675 ;
      RECT  0.15 0.675 1.7 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.445 0.47 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  0.82 1.445 0.99 1.75 ;
      RECT  1.34 1.445 1.51 1.75 ;
      RECT  1.86 1.445 2.03 1.75 ;
      RECT  2.38 1.445 2.55 1.75 ;
      RECT  2.9 1.445 3.07 1.75 ;
      RECT  3.42 1.445 3.59 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  0.56 0.05 0.73 0.35 ;
      RECT  1.08 0.05 1.25 0.35 ;
      RECT  1.6 0.05 1.77 0.35 ;
      RECT  4.985 0.05 5.155 0.375 ;
      RECT  5.505 0.05 5.675 0.375 ;
      RECT  6.025 0.05 6.195 0.375 ;
      RECT  6.59 0.05 6.71 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.1 0.435 4.65 0.535 ;
      RECT  4.505 0.535 4.65 1.11 ;
      RECT  4.35 1.11 4.65 1.245 ;
      RECT  3.92 1.245 6.69 1.36 ;
      RECT  4.985 1.36 5.155 1.365 ;
      RECT  5.505 1.36 5.675 1.365 ;
      RECT  6.55 1.36 6.69 1.5 ;
    END
    ANTENNADIFFAREA 0.881 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.68 0.225 4.875 0.33 ;
      RECT  4.75 0.33 4.875 0.475 ;
      RECT  4.75 0.475 6.48 0.595 ;
      RECT  1.89 0.225 3.59 0.335 ;
      RECT  1.89 0.335 2.0 0.44 ;
      RECT  0.34 0.32 0.445 0.44 ;
      RECT  0.34 0.44 2.0 0.545 ;
      RECT  0.065 1.21 3.83 1.32 ;
      RECT  0.065 1.32 0.185 1.435 ;
      RECT  3.705 1.32 3.83 1.485 ;
      RECT  3.705 1.485 6.46 1.6 ;
  END
END SEN_AOI22_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_T_6
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_T_6
  CLASS CORE ;
  FOREIGN SEN_AOI22_T_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.71 6.97 0.89 ;
      RECT  5.75 0.89 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.75 0.71 9.85 0.91 ;
      RECT  7.75 0.91 9.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5616 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.695 5.265 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6048 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.695 ;
      RECT  0.35 0.695 2.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6048 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.45 0.47 1.75 ;
      RECT  0.0 1.75 10.2 1.85 ;
      RECT  0.82 1.45 0.99 1.75 ;
      RECT  1.34 1.45 1.51 1.75 ;
      RECT  1.86 1.45 2.03 1.75 ;
      RECT  2.38 1.45 2.55 1.75 ;
      RECT  2.9 1.45 3.07 1.75 ;
      RECT  3.42 1.45 3.59 1.75 ;
      RECT  3.94 1.45 4.11 1.75 ;
      RECT  4.46 1.45 4.63 1.75 ;
      RECT  4.98 1.45 5.15 1.75 ;
      RECT  5.5 1.435 5.67 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      RECT  7.58 0.05 7.75 0.32 ;
      RECT  8.1 0.05 8.27 0.32 ;
      RECT  8.62 0.05 8.79 0.32 ;
      RECT  9.14 0.05 9.31 0.32 ;
      RECT  9.66 0.05 9.83 0.335 ;
      RECT  1.08 0.05 1.25 0.36 ;
      RECT  1.6 0.05 1.77 0.36 ;
      RECT  2.12 0.05 2.29 0.36 ;
      RECT  2.64 0.05 2.81 0.36 ;
      RECT  0.555 0.05 0.685 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.16 0.45 7.25 0.58 ;
      RECT  7.12 0.58 7.25 1.11 ;
      RECT  6.02 1.11 7.25 1.25 ;
      RECT  6.02 1.25 9.83 1.29 ;
      RECT  7.12 1.29 9.83 1.38 ;
      RECT  9.655 1.38 9.83 1.4 ;
    END
    ANTENNADIFFAREA 1.319 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.91 0.21 5.175 0.36 ;
      RECT  2.91 0.36 3.05 0.45 ;
      RECT  0.79 0.45 3.05 0.58 ;
      RECT  5.78 0.19 7.49 0.36 ;
      RECT  7.36 0.36 7.49 0.45 ;
      RECT  7.36 0.45 10.06 0.59 ;
      RECT  9.945 0.365 10.06 0.45 ;
      RECT  0.065 1.21 5.92 1.34 ;
      RECT  0.065 1.34 0.185 1.43 ;
      RECT  5.76 1.34 5.92 1.49 ;
      RECT  5.76 1.49 10.06 1.625 ;
      RECT  9.945 1.37 10.06 1.49 ;
  END
END SEN_AOI22_T_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI22_T_8
#      Description : "Two 2-input ANDs into 2-input NOR"
#      Equation    : X=!((A1&A2)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI22_T_8
  CLASS CORE ;
  FOREIGN SEN_AOI22_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 8.95 0.89 ;
      RECT  7.35 0.89 7.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.75 0.71 12.85 0.91 ;
      RECT  10.75 0.91 12.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7488 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.025 0.71 6.85 0.89 ;
      RECT  6.75 0.89 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.69 ;
      RECT  0.35 0.69 3.565 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.325 0.45 1.75 ;
      RECT  0.0 1.75 13.0 1.85 ;
      RECT  0.84 1.325 0.97 1.75 ;
      RECT  1.36 1.325 1.49 1.75 ;
      RECT  1.88 1.325 2.01 1.75 ;
      RECT  2.4 1.325 2.53 1.75 ;
      RECT  2.92 1.325 3.045 1.75 ;
      RECT  3.44 1.325 3.57 1.75 ;
      RECT  3.96 1.325 4.09 1.75 ;
      RECT  4.48 1.325 4.61 1.75 ;
      RECT  5.0 1.325 5.13 1.75 ;
      RECT  5.52 1.325 5.65 1.75 ;
      RECT  6.02 1.48 6.19 1.75 ;
      RECT  6.54 1.48 6.71 1.75 ;
      RECT  7.06 1.44 7.195 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 13.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
      RECT  11.85 1.75 11.95 1.85 ;
      RECT  12.45 1.75 12.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 13.0 0.05 ;
      RECT  0.815 0.05 0.99 0.36 ;
      RECT  1.34 0.05 1.51 0.36 ;
      RECT  1.86 0.05 2.03 0.36 ;
      RECT  2.38 0.05 2.55 0.36 ;
      RECT  2.9 0.05 3.07 0.36 ;
      RECT  3.42 0.05 3.59 0.36 ;
      RECT  10.18 0.05 10.35 0.395 ;
      RECT  10.7 0.05 10.87 0.395 ;
      RECT  11.22 0.05 11.39 0.395 ;
      RECT  11.74 0.05 11.91 0.395 ;
      RECT  12.26 0.05 12.43 0.395 ;
      RECT  9.68 0.05 9.82 0.41 ;
      RECT  12.805 0.05 12.925 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 13.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
      RECT  11.85 -0.05 11.95 0.05 ;
      RECT  12.45 -0.05 12.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.96 0.45 9.275 0.62 ;
      RECT  6.95 0.62 7.25 0.69 ;
      RECT  9.1 0.62 9.275 1.11 ;
      RECT  7.62 1.11 9.45 1.21 ;
      RECT  7.62 1.21 12.925 1.29 ;
      RECT  9.1 1.29 12.925 1.385 ;
    END
    ANTENNADIFFAREA 1.749 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.68 0.21 7.01 0.36 ;
      RECT  3.68 0.36 3.85 0.45 ;
      RECT  0.565 0.32 0.685 0.45 ;
      RECT  0.565 0.45 3.85 0.58 ;
      RECT  7.36 0.19 9.555 0.36 ;
      RECT  9.385 0.36 9.555 0.52 ;
      RECT  9.385 0.52 12.66 0.69 ;
      RECT  0.08 1.005 5.945 1.175 ;
      RECT  5.775 1.175 5.945 1.18 ;
      RECT  5.775 1.18 7.505 1.35 ;
      RECT  7.305 1.35 7.505 1.495 ;
      RECT  7.305 1.495 12.715 1.64 ;
  END
END SEN_AOI22_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI311_1
#      Description : "One 3-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2&A3)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI311_1
  CLASS CORE ;
  FOREIGN SEN_AOI311_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.71 0.51 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.77 ;
      RECT  0.35 0.77 0.54 0.94 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.34 0.7 1.46 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.06 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.22 0.185 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.595 1.43 0.715 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  1.12 0.05 1.24 0.365 ;
      RECT  0.065 0.05 0.185 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.8 0.24 1.03 0.36 ;
      RECT  0.94 0.36 1.03 0.455 ;
      RECT  0.94 0.455 1.525 0.575 ;
      RECT  1.15 0.575 1.25 1.395 ;
      RECT  1.15 1.395 1.505 1.575 ;
    END
    ANTENNADIFFAREA 0.258 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.295 1.22 1.03 1.34 ;
  END
END SEN_AOI311_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI311_2
#      Description : "One 3-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2&A3)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI311_2
  CLASS CORE ;
  FOREIGN SEN_AOI311_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.59 1.43 0.71 1.75 ;
      RECT  1.11 1.43 1.23 1.75 ;
      RECT  1.63 1.43 1.75 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.33 0.05 0.45 0.37 ;
      RECT  2.715 0.05 2.835 0.37 ;
      RECT  2.185 0.05 2.305 0.375 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.3 3.085 0.465 ;
      RECT  1.365 0.465 3.085 0.585 ;
      RECT  2.55 0.585 2.65 1.11 ;
      RECT  2.55 1.11 2.85 1.29 ;
    END
    ANTENNADIFFAREA 0.467 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.8 0.24 1.82 0.36 ;
      RECT  0.07 0.37 0.19 0.47 ;
      RECT  0.07 0.47 1.255 0.59 ;
      RECT  0.28 1.21 2.35 1.33 ;
      RECT  1.86 1.44 3.125 1.56 ;
  END
END SEN_AOI311_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI311_4
#      Description : "One 3-input AND into 3-input NOR"
#      Equation    : X=!((A1&A2&A3)|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI311_4
  CLASS CORE ;
  FOREIGN SEN_AOI311_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.9 ;
      RECT  2.55 0.9 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.9 ;
      RECT  1.35 0.9 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.9 ;
      RECT  0.35 0.9 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.9 ;
      RECT  3.75 0.9 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.59 1.43 0.71 1.75 ;
      RECT  1.11 1.43 1.23 1.75 ;
      RECT  1.63 1.43 1.75 1.75 ;
      RECT  2.15 1.43 2.27 1.75 ;
      RECT  2.67 1.43 2.79 1.75 ;
      RECT  3.19 1.43 3.31 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  0.33 0.05 0.45 0.37 ;
      RECT  0.85 0.05 0.97 0.37 ;
      RECT  3.73 0.05 3.85 0.37 ;
      RECT  4.25 0.05 4.37 0.37 ;
      RECT  4.77 0.05 4.89 0.37 ;
      RECT  5.295 0.05 5.415 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.405 0.46 5.715 0.58 ;
      RECT  4.75 0.58 4.85 1.11 ;
      RECT  4.75 1.11 5.45 1.29 ;
    END
    ANTENNADIFFAREA 0.851 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.32 0.2 3.38 0.32 ;
      RECT  0.07 0.36 0.19 0.46 ;
      RECT  0.07 0.46 2.295 0.58 ;
      RECT  0.305 1.22 4.42 1.34 ;
      RECT  3.42 1.44 5.705 1.56 ;
  END
END SEN_AOI311_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_0P5
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI31_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.47 1.25 0.93 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.205 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.59 1.42 0.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.14 0.05 1.29 0.38 ;
      RECT  0.06 0.05 0.2 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.855 0.28 1.05 0.4 ;
      RECT  0.95 0.4 1.05 1.04 ;
      RECT  0.95 1.04 1.26 1.13 ;
      RECT  1.14 1.13 1.26 1.565 ;
    END
    ANTENNADIFFAREA 0.105 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 1.24 1.0 1.33 ;
      RECT  0.34 1.33 0.45 1.53 ;
      RECT  0.88 1.33 1.0 1.53 ;
  END
END SEN_AOI31_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_1
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_1
  CLASS CORE ;
  FOREIGN SEN_AOI31_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.49 1.25 0.935 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.59 1.415 0.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.05 0.05 0.2 0.385 ;
      RECT  1.14 0.05 1.28 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.855 0.24 1.05 0.36 ;
      RECT  0.95 0.36 1.05 1.025 ;
      RECT  0.95 1.025 1.26 1.115 ;
      RECT  1.14 1.115 1.26 1.3 ;
    END
    ANTENNADIFFAREA 0.192 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.305 1.205 1.03 1.325 ;
  END
END SEN_AOI31_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_2
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_2
  CLASS CORE ;
  FOREIGN SEN_AOI31_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.9 ;
      RECT  1.75 0.9 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.9 ;
      RECT  0.75 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.9 ;
      RECT  2.35 0.9 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.415 0.465 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.835 1.415 0.985 1.75 ;
      RECT  1.51 1.415 1.66 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  2.135 0.05 2.285 0.37 ;
      RECT  0.315 0.05 0.465 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.36 2.53 0.465 ;
      RECT  1.345 0.465 2.53 0.585 ;
      RECT  1.95 0.585 2.05 1.02 ;
      RECT  1.95 1.02 2.26 1.11 ;
      RECT  2.14 1.11 2.26 1.29 ;
    END
    ANTENNADIFFAREA 0.37 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.79 0.24 1.81 0.36 ;
      RECT  0.07 0.37 0.19 0.48 ;
      RECT  0.07 0.48 1.255 0.59 ;
      RECT  0.07 1.21 2.015 1.32 ;
      RECT  0.07 1.32 0.19 1.43 ;
      RECT  1.885 1.32 2.015 1.51 ;
      RECT  1.885 1.51 2.53 1.63 ;
      RECT  2.41 1.41 2.53 1.51 ;
  END
END SEN_AOI31_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_3
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_3
  CLASS CORE ;
  FOREIGN SEN_AOI31_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.45 0.91 ;
      RECT  1.95 0.91 2.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 0.71 ;
      RECT  2.95 0.71 3.25 0.925 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.57 1.415 0.72 1.75 ;
      RECT  1.09 1.415 1.24 1.75 ;
      RECT  1.61 1.425 1.76 1.75 ;
      RECT  2.15 1.425 2.295 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.57 0.05 0.72 0.385 ;
      RECT  2.68 0.05 2.83 0.385 ;
      RECT  3.2 0.05 3.34 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.945 0.27 3.075 0.44 ;
      RECT  2.945 0.44 3.05 0.475 ;
      RECT  1.86 0.475 3.05 0.59 ;
      RECT  1.86 0.59 2.85 0.595 ;
      RECT  2.75 0.595 2.85 1.105 ;
      RECT  2.695 1.105 2.85 1.11 ;
      RECT  2.695 1.11 3.335 1.29 ;
    END
    ANTENNADIFFAREA 0.504 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.08 0.24 2.305 0.36 ;
      RECT  0.3 0.475 1.51 0.595 ;
      RECT  0.3 1.21 2.56 1.325 ;
      RECT  2.43 1.325 2.56 1.45 ;
      RECT  2.43 1.45 3.13 1.57 ;
  END
END SEN_AOI31_3
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_4
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_4
  CLASS CORE ;
  FOREIGN SEN_AOI31_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.9 ;
      RECT  2.75 0.9 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.9 ;
      RECT  0.35 0.9 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.415 0.465 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.835 1.415 0.985 1.75 ;
      RECT  1.385 1.415 1.535 1.75 ;
      RECT  1.975 1.415 2.125 1.75 ;
      RECT  2.525 1.415 2.675 1.75 ;
      RECT  3.045 1.415 3.195 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  3.62 0.05 3.77 0.375 ;
      RECT  4.14 0.05 4.29 0.375 ;
      RECT  0.315 0.05 0.465 0.41 ;
      RECT  0.835 0.05 0.985 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.29 0.32 2.48 0.425 ;
      RECT  2.385 0.425 2.48 0.47 ;
      RECT  2.385 0.47 4.535 0.59 ;
      RECT  4.415 0.37 4.535 0.47 ;
      RECT  3.55 0.59 3.65 1.11 ;
      RECT  3.55 1.11 4.25 1.29 ;
    END
    ANTENNADIFFAREA 0.667 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.95 0.14 2.7 0.23 ;
      RECT  1.95 0.23 2.07 0.235 ;
      RECT  2.57 0.23 2.7 0.235 ;
      RECT  1.31 0.235 2.07 0.355 ;
      RECT  2.57 0.235 3.29 0.355 ;
      RECT  0.07 0.38 0.19 0.5 ;
      RECT  0.07 0.5 2.175 0.545 ;
      RECT  0.07 0.545 2.295 0.62 ;
      RECT  2.125 0.62 2.295 0.66 ;
      RECT  0.07 1.205 3.445 1.325 ;
      RECT  3.325 1.325 3.445 1.38 ;
      RECT  0.07 1.325 0.19 1.43 ;
      RECT  3.325 1.38 4.51 1.5 ;
  END
END SEN_AOI31_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_12
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_12
  CLASS CORE ;
  FOREIGN SEN_AOI31_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.945 0.71 4.055 0.96 ;
      RECT  3.945 0.96 8.65 1.0 ;
      RECT  5.545 0.78 5.655 0.96 ;
      RECT  7.145 0.78 7.255 0.96 ;
      RECT  8.55 0.78 8.65 0.96 ;
      RECT  2.345 0.71 2.455 0.91 ;
      RECT  2.345 0.91 2.65 1.0 ;
      RECT  0.55 0.31 0.65 0.51 ;
      RECT  0.55 0.51 0.925 0.6 ;
      RECT  0.825 0.6 0.925 0.91 ;
      RECT  0.825 0.91 1.05 1.0 ;
      RECT  0.825 1.0 8.65 1.05 ;
      RECT  0.825 1.05 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.37 0.535 8.85 0.69 ;
      RECT  8.37 0.69 8.46 0.75 ;
      RECT  8.75 0.69 8.85 0.75 ;
      RECT  8.285 0.75 8.46 0.87 ;
      RECT  8.75 0.75 9.125 0.89 ;
      RECT  6.93 0.51 7.45 0.69 ;
      RECT  6.93 0.69 7.05 0.735 ;
      RECT  7.35 0.69 7.45 0.75 ;
      RECT  6.695 0.735 7.05 0.87 ;
      RECT  7.35 0.75 7.595 0.87 ;
      RECT  5.35 0.51 5.85 0.69 ;
      RECT  5.35 0.69 5.45 0.73 ;
      RECT  5.76 0.69 5.85 0.75 ;
      RECT  5.135 0.73 5.45 0.87 ;
      RECT  5.76 0.75 6.035 0.87 ;
      RECT  4.345 0.51 4.445 0.755 ;
      RECT  4.345 0.755 4.53 0.87 ;
      RECT  3.75 0.51 3.85 0.775 ;
      RECT  3.575 0.775 3.85 0.895 ;
      RECT  2.745 0.51 2.85 0.71 ;
      RECT  2.745 0.71 3.05 0.89 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.35 0.71 0.645 0.9 ;
      LAYER M2 ;
      RECT  0.31 0.55 8.79 0.65 ;
      LAYER V1 ;
      RECT  8.45 0.55 8.55 0.65 ;
      RECT  8.65 0.55 8.75 0.65 ;
      RECT  7.05 0.55 7.15 0.65 ;
      RECT  7.25 0.55 7.35 0.65 ;
      RECT  5.45 0.55 5.55 0.65 ;
      RECT  5.65 0.55 5.75 0.65 ;
      RECT  4.345 0.55 4.445 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  2.15 0.55 2.25 0.65 ;
      RECT  1.15 0.55 1.25 0.65 ;
      RECT  0.35 0.55 0.45 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.215 0.75 9.56 0.895 ;
      RECT  7.76 0.75 8.14 0.87 ;
      RECT  6.205 0.735 6.59 0.87 ;
      RECT  4.62 0.735 5.02 0.87 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  0.15 0.51 0.255 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.75 9.395 0.85 ;
      LAYER V1 ;
      RECT  9.255 0.75 9.355 0.85 ;
      RECT  7.8 0.75 7.9 0.85 ;
      RECT  8.0 0.75 8.1 0.85 ;
      RECT  6.25 0.75 6.35 0.85 ;
      RECT  6.45 0.75 6.55 0.85 ;
      RECT  4.66 0.75 4.76 0.85 ;
      RECT  4.86 0.75 4.96 0.85 ;
      RECT  3.15 0.75 3.25 0.85 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.15 0.75 0.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.13 0.71 12.65 0.89 ;
      RECT  12.55 0.89 12.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.756 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  1.36 1.415 1.49 1.75 ;
      RECT  1.88 1.415 2.01 1.75 ;
      RECT  2.4 1.415 2.53 1.75 ;
      RECT  2.92 1.415 3.05 1.75 ;
      RECT  3.44 1.415 3.57 1.75 ;
      RECT  3.96 1.415 4.09 1.75 ;
      RECT  4.48 1.415 4.61 1.75 ;
      RECT  5.0 1.415 5.13 1.75 ;
      RECT  5.52 1.415 5.65 1.75 ;
      RECT  6.04 1.415 6.165 1.75 ;
      RECT  6.54 1.48 6.71 1.75 ;
      RECT  7.06 1.48 7.23 1.75 ;
      RECT  7.58 1.48 7.75 1.75 ;
      RECT  8.1 1.48 8.27 1.75 ;
      RECT  8.62 1.48 8.79 1.75 ;
      RECT  9.14 1.48 9.31 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  9.425 0.05 9.595 0.32 ;
      RECT  9.975 0.05 10.145 0.32 ;
      RECT  10.495 0.05 10.665 0.32 ;
      RECT  7.86 0.05 7.98 0.36 ;
      RECT  11.04 0.05 11.16 0.36 ;
      RECT  11.56 0.05 11.68 0.36 ;
      RECT  12.08 0.05 12.2 0.36 ;
      RECT  1.62 0.05 1.75 0.385 ;
      RECT  3.18 0.05 3.31 0.385 ;
      RECT  4.75 0.05 4.87 0.385 ;
      RECT  6.3 0.05 6.43 0.385 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  12.61 0.05 12.73 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.07 0.175 9.25 0.41 ;
      RECT  8.07 0.41 10.51 0.425 ;
      RECT  8.07 0.425 8.28 0.45 ;
      RECT  8.95 0.425 10.51 0.45 ;
      RECT  6.55 0.175 7.75 0.385 ;
      RECT  7.54 0.385 7.75 0.45 ;
      RECT  6.55 0.385 6.72 0.475 ;
      RECT  7.54 0.45 8.28 0.66 ;
      RECT  8.95 0.45 12.51 0.575 ;
      RECT  5.125 0.215 6.12 0.385 ;
      RECT  5.125 0.385 5.25 0.475 ;
      RECT  5.95 0.385 6.12 0.475 ;
      RECT  3.44 0.235 4.66 0.36 ;
      RECT  3.44 0.36 3.565 0.475 ;
      RECT  4.535 0.36 4.66 0.475 ;
      RECT  1.95 0.24 3.065 0.36 ;
      RECT  1.95 0.36 2.05 0.475 ;
      RECT  2.94 0.36 3.065 0.475 ;
      RECT  0.79 0.24 1.45 0.36 ;
      RECT  1.35 0.36 1.45 0.475 ;
      RECT  1.35 0.475 2.05 0.565 ;
      RECT  2.94 0.475 3.565 0.6 ;
      RECT  4.535 0.475 5.25 0.605 ;
      RECT  5.95 0.475 6.72 0.645 ;
      RECT  8.95 0.575 11.115 0.62 ;
      RECT  8.95 0.62 9.99 0.66 ;
      RECT  9.74 0.66 9.99 1.11 ;
      RECT  9.74 1.11 12.46 1.29 ;
    END
    ANTENNADIFFAREA 1.836 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.15 1.14 6.49 1.16 ;
      RECT  4.15 1.16 9.65 1.205 ;
      RECT  8.275 1.14 9.65 1.16 ;
      RECT  0.065 1.205 9.65 1.325 ;
      RECT  6.255 1.325 9.65 1.39 ;
      RECT  0.065 1.325 0.185 1.43 ;
      RECT  9.4 1.39 9.65 1.4 ;
      RECT  9.4 1.4 12.72 1.52 ;
      RECT  12.6 1.3 12.72 1.4 ;
      RECT  9.4 1.52 11.35 1.58 ;
      RECT  9.4 1.58 10.32 1.615 ;
  END
END SEN_AOI31_12
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_6
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_6
  CLASS CORE ;
  FOREIGN SEN_AOI31_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.51 ;
      RECT  0.55 0.51 0.945 0.6 ;
      RECT  0.835 0.6 0.945 0.91 ;
      RECT  0.835 0.91 1.05 1.0 ;
      RECT  0.835 1.0 4.25 1.09 ;
      RECT  2.345 0.81 2.65 1.0 ;
      RECT  2.95 0.91 3.05 1.0 ;
      RECT  3.945 0.78 4.25 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.51 4.45 0.69 ;
      RECT  3.75 0.69 3.85 0.71 ;
      RECT  4.35 0.69 4.45 0.925 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  2.15 0.51 2.85 0.69 ;
      RECT  2.15 0.69 2.25 0.71 ;
      RECT  2.75 0.69 2.85 0.9 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  0.35 0.51 0.45 0.715 ;
      RECT  0.35 0.715 0.65 0.89 ;
      LAYER M2 ;
      RECT  0.31 0.55 4.29 0.65 ;
      LAYER V1 ;
      RECT  3.95 0.55 4.05 0.65 ;
      RECT  4.15 0.55 4.25 0.65 ;
      RECT  2.35 0.55 2.45 0.65 ;
      RECT  2.55 0.55 2.65 0.65 ;
      RECT  1.15 0.55 1.25 0.65 ;
      RECT  0.35 0.55 0.45 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.85 0.89 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  0.15 0.51 0.25 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.75 4.89 0.85 ;
      LAYER V1 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  3.15 0.75 3.25 0.85 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.15 0.75 0.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.325 0.71 6.45 0.89 ;
      RECT  6.35 0.89 6.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.378 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.455 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.845 1.415 0.975 1.75 ;
      RECT  1.365 1.415 1.495 1.75 ;
      RECT  1.885 1.415 2.015 1.75 ;
      RECT  2.405 1.415 2.535 1.75 ;
      RECT  2.925 1.415 3.055 1.75 ;
      RECT  3.445 1.415 3.575 1.75 ;
      RECT  3.965 1.415 4.095 1.75 ;
      RECT  4.485 1.415 4.615 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.63 0.05 1.755 0.385 ;
      RECT  3.185 0.05 3.315 0.385 ;
      RECT  4.76 0.05 4.89 0.385 ;
      RECT  5.295 0.05 5.425 0.385 ;
      RECT  5.815 0.05 5.945 0.385 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  6.36 0.05 6.48 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.235 4.67 0.365 ;
      RECT  4.54 0.365 4.67 0.475 ;
      RECT  3.55 0.365 3.65 0.49 ;
      RECT  4.54 0.475 6.25 0.605 ;
      RECT  1.95 0.24 3.05 0.36 ;
      RECT  1.95 0.36 2.05 0.49 ;
      RECT  2.95 0.36 3.05 0.49 ;
      RECT  0.795 0.24 1.45 0.36 ;
      RECT  1.35 0.36 1.45 0.49 ;
      RECT  1.35 0.49 2.05 0.58 ;
      RECT  2.95 0.49 3.65 0.58 ;
      RECT  4.95 0.605 5.08 1.11 ;
      RECT  4.95 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 0.918 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.18 4.86 1.31 ;
      RECT  0.07 1.31 0.19 1.4 ;
      RECT  4.73 1.31 4.86 1.435 ;
      RECT  4.73 1.435 6.51 1.565 ;
  END
END SEN_AOI31_6
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_8
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_8
  CLASS CORE ;
  FOREIGN SEN_AOI31_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.51 ;
      RECT  0.55 0.51 0.955 0.6 ;
      RECT  0.845 0.6 0.955 0.91 ;
      RECT  0.845 0.91 1.05 1.0 ;
      RECT  0.845 1.0 5.655 1.09 ;
      RECT  2.345 0.81 2.65 1.0 ;
      RECT  2.95 0.91 3.05 1.0 ;
      RECT  3.945 0.78 4.25 1.0 ;
      RECT  4.55 0.91 4.65 1.0 ;
      RECT  5.545 0.75 5.655 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.51 5.85 0.655 ;
      RECT  5.35 0.655 5.45 0.71 ;
      RECT  5.75 0.655 5.85 0.71 ;
      RECT  5.15 0.71 5.45 0.89 ;
      RECT  5.75 0.71 6.04 0.89 ;
      RECT  3.75 0.51 4.45 0.69 ;
      RECT  3.75 0.69 3.85 0.71 ;
      RECT  4.35 0.69 4.45 0.9 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  2.15 0.51 2.85 0.69 ;
      RECT  2.15 0.69 2.25 0.71 ;
      RECT  2.75 0.69 2.85 0.9 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  0.35 0.51 0.45 0.715 ;
      RECT  0.35 0.715 0.65 0.89 ;
      LAYER M2 ;
      RECT  0.31 0.55 5.79 0.65 ;
      LAYER V1 ;
      RECT  5.45 0.55 5.55 0.65 ;
      RECT  5.65 0.55 5.75 0.65 ;
      RECT  3.95 0.55 4.05 0.65 ;
      RECT  4.15 0.55 4.25 0.65 ;
      RECT  2.35 0.55 2.45 0.65 ;
      RECT  2.55 0.55 2.65 0.65 ;
      RECT  1.15 0.55 1.25 0.65 ;
      RECT  0.35 0.55 0.45 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.45 0.89 ;
      RECT  4.75 0.71 5.05 0.89 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  0.15 0.51 0.25 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.75 6.29 0.85 ;
      LAYER V1 ;
      RECT  6.15 0.75 6.25 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
      RECT  3.15 0.75 3.25 0.85 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.15 0.75 0.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.93 0.71 8.45 0.89 ;
      RECT  8.35 0.89 8.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.4 0.455 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.845 1.4 0.975 1.75 ;
      RECT  1.365 1.4 1.495 1.75 ;
      RECT  1.885 1.4 2.015 1.75 ;
      RECT  2.405 1.4 2.535 1.75 ;
      RECT  2.925 1.415 3.055 1.75 ;
      RECT  3.445 1.44 3.575 1.75 ;
      RECT  3.965 1.44 4.095 1.75 ;
      RECT  4.485 1.44 4.615 1.75 ;
      RECT  5.005 1.44 5.135 1.75 ;
      RECT  5.525 1.44 5.655 1.75 ;
      RECT  6.045 1.44 6.175 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  6.305 0.05 6.435 0.36 ;
      RECT  4.76 0.05 4.875 0.385 ;
      RECT  6.825 0.05 6.955 0.385 ;
      RECT  7.345 0.05 7.475 0.385 ;
      RECT  7.865 0.05 7.995 0.385 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  1.625 0.05 1.755 0.39 ;
      RECT  3.185 0.05 3.315 0.39 ;
      RECT  8.4 0.05 8.52 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.12 0.215 6.135 0.385 ;
      RECT  5.95 0.385 6.135 0.45 ;
      RECT  5.12 0.385 5.25 0.475 ;
      RECT  5.95 0.45 6.72 0.475 ;
      RECT  3.55 0.235 4.67 0.365 ;
      RECT  4.54 0.365 4.67 0.475 ;
      RECT  3.55 0.365 3.65 0.49 ;
      RECT  4.54 0.475 5.25 0.605 ;
      RECT  5.95 0.475 8.3 0.605 ;
      RECT  1.95 0.24 3.05 0.36 ;
      RECT  1.95 0.36 2.05 0.49 ;
      RECT  2.95 0.36 3.05 0.49 ;
      RECT  0.8 0.24 1.45 0.36 ;
      RECT  1.35 0.36 1.45 0.49 ;
      RECT  1.35 0.49 2.05 0.58 ;
      RECT  2.95 0.49 3.65 0.58 ;
      RECT  5.95 0.605 6.72 0.62 ;
      RECT  6.55 0.62 6.72 1.11 ;
      RECT  6.55 1.11 8.25 1.29 ;
    END
    ANTENNADIFFAREA 1.224 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.18 6.455 1.3 ;
      RECT  3.39 1.3 6.455 1.35 ;
      RECT  0.07 1.3 0.19 1.4 ;
      RECT  6.285 1.35 6.455 1.43 ;
      RECT  6.285 1.43 8.51 1.57 ;
      RECT  8.39 1.35 8.51 1.43 ;
  END
END SEN_AOI31_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_G_8
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_G_8
  CLASS CORE ;
  FOREIGN SEN_AOI31_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.51 ;
      RECT  0.55 0.51 0.945 0.6 ;
      RECT  0.835 0.6 0.945 0.91 ;
      RECT  0.835 0.91 1.05 1.0 ;
      RECT  0.835 1.0 5.655 1.09 ;
      RECT  2.345 0.81 2.65 1.0 ;
      RECT  2.95 0.91 3.05 1.0 ;
      RECT  3.945 0.78 4.25 1.0 ;
      RECT  4.55 0.91 4.65 1.0 ;
      RECT  5.545 0.78 5.655 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.51 5.85 0.69 ;
      RECT  5.35 0.69 5.45 0.71 ;
      RECT  5.75 0.69 5.85 0.71 ;
      RECT  5.15 0.71 5.45 0.89 ;
      RECT  5.75 0.71 6.04 0.89 ;
      RECT  3.75 0.51 4.45 0.69 ;
      RECT  3.75 0.69 3.85 0.71 ;
      RECT  4.35 0.69 4.45 0.9 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  2.15 0.51 2.85 0.69 ;
      RECT  2.15 0.69 2.25 0.71 ;
      RECT  2.75 0.69 2.85 0.9 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  0.35 0.51 0.45 0.715 ;
      RECT  0.35 0.715 0.65 0.89 ;
      LAYER M2 ;
      RECT  0.31 0.55 5.79 0.65 ;
      LAYER V1 ;
      RECT  5.45 0.55 5.55 0.65 ;
      RECT  5.65 0.55 5.75 0.65 ;
      RECT  3.95 0.55 4.05 0.65 ;
      RECT  4.15 0.55 4.25 0.65 ;
      RECT  2.35 0.55 2.45 0.65 ;
      RECT  2.55 0.55 2.65 0.65 ;
      RECT  1.15 0.55 1.25 0.65 ;
      RECT  0.35 0.55 0.45 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.45 0.89 ;
      RECT  4.75 0.71 5.05 0.89 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  0.15 0.51 0.25 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.75 6.29 0.85 ;
      LAYER V1 ;
      RECT  6.15 0.75 6.25 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
      RECT  3.15 0.75 3.25 0.85 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.15 0.75 0.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.93 0.71 8.45 0.89 ;
      RECT  8.35 0.89 8.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.455 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.845 1.415 0.975 1.75 ;
      RECT  1.365 1.415 1.495 1.75 ;
      RECT  1.885 1.415 2.015 1.75 ;
      RECT  2.405 1.415 2.535 1.75 ;
      RECT  2.925 1.415 3.055 1.75 ;
      RECT  3.445 1.44 3.575 1.75 ;
      RECT  3.965 1.44 4.095 1.75 ;
      RECT  4.485 1.44 4.615 1.75 ;
      RECT  5.005 1.44 5.135 1.75 ;
      RECT  5.525 1.44 5.655 1.75 ;
      RECT  6.045 1.44 6.175 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  6.305 0.05 6.435 0.36 ;
      RECT  4.76 0.05 4.875 0.385 ;
      RECT  6.825 0.05 6.955 0.385 ;
      RECT  7.345 0.05 7.475 0.385 ;
      RECT  7.865 0.05 7.995 0.385 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  1.625 0.05 1.755 0.39 ;
      RECT  3.185 0.05 3.315 0.39 ;
      RECT  8.4 0.05 8.52 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.12 0.215 6.135 0.385 ;
      RECT  5.95 0.385 6.135 0.45 ;
      RECT  5.12 0.385 5.25 0.475 ;
      RECT  5.95 0.45 6.72 0.475 ;
      RECT  3.55 0.235 4.67 0.365 ;
      RECT  4.54 0.365 4.67 0.475 ;
      RECT  3.55 0.365 3.65 0.49 ;
      RECT  4.54 0.475 5.25 0.605 ;
      RECT  5.95 0.475 8.3 0.605 ;
      RECT  1.95 0.24 3.05 0.36 ;
      RECT  1.95 0.36 2.05 0.49 ;
      RECT  2.95 0.36 3.05 0.49 ;
      RECT  0.79 0.24 1.45 0.36 ;
      RECT  1.35 0.36 1.45 0.49 ;
      RECT  1.35 0.49 2.05 0.58 ;
      RECT  2.95 0.49 3.65 0.58 ;
      RECT  5.95 0.605 6.72 0.62 ;
      RECT  6.55 0.62 6.72 1.11 ;
      RECT  6.55 1.11 8.25 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.18 6.455 1.3 ;
      RECT  3.39 1.3 6.455 1.35 ;
      RECT  0.07 1.3 0.19 1.41 ;
      RECT  6.285 1.35 6.455 1.43 ;
      RECT  6.285 1.43 8.545 1.57 ;
  END
END SEN_AOI31_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_0P75
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_0P75
  CLASS CORE ;
  FOREIGN SEN_AOI31_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.5 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.3 0.65 0.71 ;
      RECT  0.35 0.71 0.65 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.6 1.415 0.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.155 0.05 1.325 0.22 ;
      RECT  0.065 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.825 0.24 1.05 0.36 ;
      RECT  0.95 0.36 1.05 1.01 ;
      RECT  0.95 1.01 1.25 1.1 ;
      RECT  1.15 1.1 1.25 1.49 ;
    END
    ANTENNADIFFAREA 0.141 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 1.205 1.055 1.325 ;
  END
END SEN_AOI31_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_T_0P5
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_T_0P5
  CLASS CORE ;
  FOREIGN SEN_AOI31_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.5 0.86 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.3 0.65 0.71 ;
      RECT  0.35 0.71 0.65 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.59 1.415 0.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.155 0.05 1.325 0.22 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.815 0.24 1.05 0.36 ;
      RECT  0.95 0.36 1.05 1.01 ;
      RECT  0.95 1.01 1.25 1.1 ;
      RECT  1.15 1.1 1.25 1.53 ;
    END
    ANTENNADIFFAREA 0.1 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 1.205 1.05 1.325 ;
  END
END SEN_AOI31_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_T_1
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_T_1
  CLASS CORE ;
  FOREIGN SEN_AOI31_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.5 0.65 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.71 ;
      RECT  1.75 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.455 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  0.845 1.415 0.975 1.75 ;
      RECT  1.39 1.415 1.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  1.955 0.05 2.085 0.39 ;
      RECT  0.3 0.05 0.42 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.85 0.49 ;
      RECT  1.55 0.49 1.65 1.02 ;
      RECT  1.55 1.02 2.06 1.11 ;
      RECT  1.94 1.11 2.06 1.29 ;
    END
    ANTENNADIFFAREA 0.189 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.795 0.23 1.46 0.35 ;
      RECT  0.07 1.205 1.85 1.325 ;
      RECT  0.07 1.325 0.19 1.43 ;
  END
END SEN_AOI31_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_T_2
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_T_2
  CLASS CORE ;
  FOREIGN SEN_AOI31_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.64 2.65 0.89 ;
      RECT  2.15 0.89 2.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.64 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.845 1.415 0.965 1.75 ;
      RECT  1.38 1.415 1.5 1.75 ;
      RECT  1.93 1.415 2.05 1.75 ;
      RECT  2.47 1.415 2.59 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  3.34 0.05 3.46 0.35 ;
      RECT  0.325 0.05 0.445 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.925 0.32 2.095 0.44 ;
      RECT  1.925 0.44 3.745 0.53 ;
      RECT  2.445 0.32 2.615 0.44 ;
      RECT  3.04 0.22 3.16 0.44 ;
      RECT  3.35 0.53 3.745 0.55 ;
      RECT  3.35 0.55 3.45 1.29 ;
    END
    ANTENNADIFFAREA 0.376 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.14 2.85 0.23 ;
      RECT  2.21 0.23 2.33 0.345 ;
      RECT  2.73 0.23 2.85 0.345 ;
      RECT  1.365 0.23 1.485 0.35 ;
      RECT  0.845 0.23 0.965 0.36 ;
      RECT  1.08 0.32 1.25 0.44 ;
      RECT  1.08 0.44 1.77 0.475 ;
      RECT  1.6 0.32 1.77 0.44 ;
      RECT  0.065 0.37 0.185 0.475 ;
      RECT  0.065 0.475 1.77 0.53 ;
      RECT  0.585 0.24 0.705 0.475 ;
      RECT  0.065 0.53 1.25 0.595 ;
      RECT  0.065 1.205 3.06 1.325 ;
      RECT  0.065 1.325 0.185 1.43 ;
      RECT  2.94 1.325 3.06 1.44 ;
      RECT  2.94 1.44 3.745 1.56 ;
  END
END SEN_AOI31_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_T_4
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_T_4
  CLASS CORE ;
  FOREIGN SEN_AOI31_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.655 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.68 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.675 5.85 0.89 ;
      RECT  5.75 0.89 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.365 1.415 1.495 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.885 1.415 2.015 1.75 ;
      RECT  2.405 1.415 2.535 1.75 ;
      RECT  2.925 1.415 3.055 1.75 ;
      RECT  3.465 1.415 3.595 1.75 ;
      RECT  3.985 1.415 4.115 1.75 ;
      RECT  4.51 1.415 4.64 1.75 ;
      RECT  5.04 1.415 5.17 1.75 ;
      RECT  5.56 1.415 5.69 1.75 ;
      RECT  6.08 1.415 6.21 1.75 ;
      RECT  6.605 1.21 6.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  0.825 0.05 0.995 0.315 ;
      RECT  0.325 0.05 0.455 0.385 ;
      RECT  4.78 0.05 4.91 0.385 ;
      RECT  5.3 0.05 5.43 0.385 ;
      RECT  5.82 0.05 5.95 0.385 ;
      RECT  6.37 0.05 6.5 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.07 0.365 0.19 0.475 ;
      RECT  0.07 0.475 2.845 0.52 ;
      RECT  0.95 0.405 2.845 0.475 ;
      RECT  0.07 0.52 1.05 0.595 ;
      RECT  0.95 0.595 1.05 1.11 ;
      RECT  0.34 1.11 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.667 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.31 0.2 4.69 0.315 ;
      RECT  3.195 0.405 4.405 0.475 ;
      RECT  3.195 0.475 6.205 0.52 ;
      RECT  5.045 0.29 5.165 0.475 ;
      RECT  5.565 0.29 5.685 0.475 ;
      RECT  6.085 0.29 6.205 0.475 ;
      RECT  4.305 0.52 6.205 0.565 ;
      RECT  1.155 1.205 6.515 1.325 ;
      RECT  1.155 1.325 1.255 1.44 ;
      RECT  0.07 1.34 0.19 1.44 ;
      RECT  0.07 1.44 1.255 1.56 ;
  END
END SEN_AOI31_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_T_8
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_T_8
  CLASS CORE ;
  FOREIGN SEN_AOI31_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.64 9.45 0.775 ;
      RECT  7.95 0.775 8.25 0.89 ;
      RECT  9.15 0.775 9.45 0.89 ;
      RECT  9.35 0.89 9.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.665 6.05 0.89 ;
      RECT  5.95 0.89 6.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.665 2.45 0.77 ;
      RECT  0.95 0.77 1.25 0.89 ;
      RECT  2.15 0.77 2.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.93 0.71 12.45 0.89 ;
      RECT  12.35 0.89 12.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 12.6 1.85 ;
      RECT  0.58 1.415 0.71 1.75 ;
      RECT  1.1 1.415 1.23 1.75 ;
      RECT  1.62 1.415 1.75 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  2.66 1.44 2.79 1.75 ;
      RECT  3.18 1.44 3.31 1.75 ;
      RECT  3.7 1.44 3.83 1.75 ;
      RECT  4.22 1.44 4.35 1.75 ;
      RECT  4.74 1.44 4.87 1.75 ;
      RECT  5.26 1.44 5.39 1.75 ;
      RECT  5.78 1.44 5.91 1.75 ;
      RECT  6.3 1.44 6.43 1.75 ;
      RECT  6.88 1.44 7.01 1.75 ;
      RECT  7.46 1.44 7.59 1.75 ;
      RECT  7.98 1.44 8.11 1.75 ;
      RECT  8.5 1.44 8.63 1.75 ;
      RECT  9.02 1.44 9.15 1.75 ;
      RECT  9.54 1.44 9.67 1.75 ;
      RECT  10.06 1.44 10.19 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.6 0.05 ;
      RECT  2.64 0.05 2.81 0.315 ;
      RECT  3.16 0.05 3.33 0.315 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  10.58 0.05 10.71 0.365 ;
      RECT  11.1 0.05 11.23 0.365 ;
      RECT  11.62 0.05 11.75 0.365 ;
      RECT  12.14 0.05 12.27 0.365 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.1 0.05 1.23 0.385 ;
      RECT  1.62 0.05 1.75 0.385 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.26 0.375 9.43 0.4 ;
      RECT  9.26 0.4 10.45 0.425 ;
      RECT  9.78 0.375 9.95 0.4 ;
      RECT  10.32 0.255 10.45 0.4 ;
      RECT  8.74 0.375 8.91 0.425 ;
      RECT  8.74 0.425 10.45 0.45 ;
      RECT  8.22 0.375 8.39 0.45 ;
      RECT  8.22 0.45 10.45 0.455 ;
      RECT  8.22 0.455 12.525 0.46 ;
      RECT  12.405 0.375 12.525 0.455 ;
      RECT  7.18 0.38 7.35 0.46 ;
      RECT  7.18 0.46 12.525 0.55 ;
      RECT  7.7 0.38 7.87 0.46 ;
      RECT  10.15 0.55 12.525 0.595 ;
      RECT  10.15 0.595 10.72 0.69 ;
      RECT  10.55 0.69 10.72 1.11 ;
      RECT  10.55 1.11 12.26 1.29 ;
    END
    ANTENNADIFFAREA 1.26 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.68 0.14 10.21 0.23 ;
      RECT  4.72 0.23 9.17 0.24 ;
      RECT  9.52 0.23 9.69 0.31 ;
      RECT  10.04 0.23 10.21 0.31 ;
      RECT  3.68 0.23 3.85 0.315 ;
      RECT  4.2 0.23 4.37 0.315 ;
      RECT  5.24 0.24 8.65 0.265 ;
      RECT  4.72 0.24 4.89 0.32 ;
      RECT  9.0 0.24 9.17 0.32 ;
      RECT  5.76 0.265 8.13 0.29 ;
      RECT  5.24 0.265 5.41 0.32 ;
      RECT  8.48 0.265 8.65 0.32 ;
      RECT  6.77 0.29 7.12 0.31 ;
      RECT  5.76 0.29 5.93 0.32 ;
      RECT  6.28 0.29 6.45 0.32 ;
      RECT  7.44 0.29 7.61 0.32 ;
      RECT  7.96 0.29 8.13 0.32 ;
      RECT  2.405 0.26 2.525 0.405 ;
      RECT  2.405 0.405 4.63 0.43 ;
      RECT  2.925 0.265 3.045 0.405 ;
      RECT  3.445 0.26 3.565 0.405 ;
      RECT  3.94 0.375 4.11 0.405 ;
      RECT  4.46 0.375 4.63 0.405 ;
      RECT  2.405 0.43 5.15 0.44 ;
      RECT  4.98 0.375 5.15 0.43 ;
      RECT  2.405 0.44 6.71 0.45 ;
      RECT  5.5 0.375 5.67 0.44 ;
      RECT  6.02 0.38 6.19 0.44 ;
      RECT  6.54 0.38 6.71 0.44 ;
      RECT  1.885 0.26 2.005 0.45 ;
      RECT  1.885 0.45 6.71 0.475 ;
      RECT  1.365 0.26 1.485 0.475 ;
      RECT  1.365 0.475 6.71 0.485 ;
      RECT  0.325 0.26 0.445 0.485 ;
      RECT  0.325 0.485 6.71 0.53 ;
      RECT  0.845 0.26 0.965 0.485 ;
      RECT  0.325 0.53 4.63 0.575 ;
      RECT  0.3 1.18 10.46 1.305 ;
      RECT  2.15 1.305 10.46 1.35 ;
      RECT  10.29 1.35 10.46 1.43 ;
      RECT  10.29 1.43 12.525 1.57 ;
      RECT  12.405 1.35 12.525 1.43 ;
  END
END SEN_AOI31_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_G_1
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_G_1
  CLASS CORE ;
  FOREIGN SEN_AOI31_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.5 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.3 0.65 0.71 ;
      RECT  0.35 0.71 0.65 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.925 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.6 1.41 0.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.155 0.05 1.325 0.22 ;
      RECT  0.065 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.83 0.24 1.05 0.36 ;
      RECT  0.95 0.36 1.05 1.035 ;
      RECT  0.95 1.035 1.25 1.125 ;
      RECT  1.15 1.125 1.25 1.49 ;
    END
    ANTENNADIFFAREA 0.192 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 1.22 1.0 1.32 ;
      RECT  0.88 1.32 1.0 1.44 ;
  END
END SEN_AOI31_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_G_2
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_G_2
  CLASS CORE ;
  FOREIGN SEN_AOI31_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.585 1.415 0.715 1.75 ;
      RECT  1.105 1.415 1.235 1.75 ;
      RECT  1.625 1.415 1.755 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.325 0.05 0.455 0.385 ;
      RECT  2.145 0.05 2.275 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.37 2.53 0.475 ;
      RECT  1.345 0.475 2.53 0.595 ;
      RECT  1.95 0.595 2.05 1.02 ;
      RECT  1.95 1.02 2.26 1.11 ;
      RECT  2.15 1.11 2.26 1.29 ;
    END
    ANTENNADIFFAREA 0.37 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.795 0.23 1.805 0.35 ;
      RECT  0.07 0.365 0.19 0.475 ;
      RECT  0.07 0.475 1.255 0.595 ;
      RECT  0.28 1.205 2.01 1.325 ;
      RECT  1.89 1.325 2.01 1.44 ;
      RECT  1.89 1.44 2.53 1.56 ;
      RECT  2.41 1.335 2.53 1.44 ;
  END
END SEN_AOI31_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI31_G_4
#      Description : "One 3-input AND into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI31_G_4
  CLASS CORE ;
  FOREIGN SEN_AOI31_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  2.75 0.89 2.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.05 0.89 ;
      RECT  0.55 0.89 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.7 4.65 0.89 ;
      RECT  4.55 0.89 4.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.14 1.21 0.26 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.655 1.415 0.785 1.75 ;
      RECT  1.175 1.415 1.305 1.75 ;
      RECT  1.695 1.415 1.825 1.75 ;
      RECT  2.215 1.415 2.345 1.75 ;
      RECT  2.755 1.415 2.885 1.75 ;
      RECT  3.275 1.415 3.405 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.395 0.05 0.525 0.385 ;
      RECT  0.915 0.05 1.045 0.385 ;
      RECT  3.795 0.05 3.925 0.385 ;
      RECT  4.315 0.05 4.445 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.31 4.7 0.475 ;
      RECT  2.475 0.475 4.7 0.595 ;
      RECT  3.35 0.595 3.85 0.69 ;
      RECT  3.75 0.69 3.85 1.11 ;
      RECT  3.75 1.11 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.682 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.39 0.24 3.45 0.36 ;
      RECT  0.09 0.475 2.365 0.595 ;
      RECT  0.35 1.205 3.66 1.325 ;
      RECT  3.54 1.325 3.66 1.44 ;
      RECT  3.54 1.44 4.7 1.56 ;
      RECT  4.58 1.335 4.7 1.44 ;
  END
END SEN_AOI31_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI32_1
#      Description : "One 3-input AND one 2-input AND into into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI32_1
  CLASS CORE ;
  FOREIGN SEN_AOI32_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.725 0.51 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.79 ;
      RECT  0.35 0.79 0.575 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.5 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.5 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.58 1.41 0.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.05 0.05 0.2 0.39 ;
      RECT  1.395 0.05 1.545 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.82 0.24 1.26 0.36 ;
      RECT  1.14 0.36 1.26 1.3 ;
    END
    ANTENNADIFFAREA 0.224 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.3 1.2 1.0 1.32 ;
      RECT  0.87 1.32 1.0 1.515 ;
      RECT  0.87 1.515 1.52 1.63 ;
      RECT  1.4 1.41 1.52 1.515 ;
  END
END SEN_AOI32_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI32_2
#      Description : "One 3-input AND one 2-input AND into into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI32_2
  CLASS CORE ;
  FOREIGN SEN_AOI32_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.9 ;
      RECT  1.55 0.9 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.9 ;
      RECT  0.95 0.9 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.7 2.65 0.9 ;
      RECT  2.55 0.9 2.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.7 3.25 0.9 ;
      RECT  3.15 0.9 3.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.47 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  1.015 1.41 1.165 1.75 ;
      RECT  1.7 1.41 1.85 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.05 0.05 0.2 0.39 ;
      RECT  0.59 0.05 0.74 0.39 ;
      RECT  2.92 0.05 3.07 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.58 0.47 2.58 0.59 ;
      RECT  2.15 0.59 2.25 1.225 ;
      RECT  2.15 1.225 3.05 1.345 ;
      RECT  2.94 1.11 3.05 1.225 ;
    END
    ANTENNADIFFAREA 0.458 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.83 0.24 2.04 0.36 ;
      RECT  2.13 0.24 2.795 0.36 ;
      RECT  2.675 0.36 2.795 0.48 ;
      RECT  2.675 0.48 3.315 0.59 ;
      RECT  3.195 0.37 3.315 0.48 ;
      RECT  0.28 0.48 1.29 0.59 ;
      RECT  0.065 1.21 2.06 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  1.94 1.32 2.06 1.44 ;
      RECT  1.94 1.44 3.315 1.55 ;
      RECT  3.195 1.33 3.315 1.44 ;
  END
END SEN_AOI32_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI32_4
#      Description : "One 3-input AND one 2-input AND into into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI32_4
  CLASS CORE ;
  FOREIGN SEN_AOI32_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.9 ;
      RECT  2.75 0.9 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.7 2.05 0.9 ;
      RECT  1.55 0.9 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.45 0.9 ;
      RECT  3.75 0.9 3.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.71 5.85 0.9 ;
      RECT  5.75 0.9 5.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.355 1.415 0.505 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.925 1.415 1.07 1.75 ;
      RECT  1.505 1.425 1.655 1.75 ;
      RECT  2.09 1.415 2.24 1.75 ;
      RECT  2.715 1.415 2.865 1.75 ;
      RECT  3.365 1.415 3.515 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  0.065 0.05 0.215 0.385 ;
      RECT  0.585 0.05 0.735 0.385 ;
      RECT  1.105 0.05 1.255 0.385 ;
      RECT  4.995 0.05 5.145 0.385 ;
      RECT  5.515 0.05 5.665 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.645 0.47 4.66 0.59 ;
      RECT  4.55 0.59 4.66 1.11 ;
      RECT  3.945 1.11 5.655 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.345 0.23 3.595 0.35 ;
      RECT  3.685 0.23 4.87 0.35 ;
      RECT  4.75 0.35 4.87 0.485 ;
      RECT  4.75 0.485 5.91 0.605 ;
      RECT  5.79 0.38 5.91 0.485 ;
      RECT  0.28 0.49 2.295 0.61 ;
      RECT  0.08 1.205 3.84 1.325 ;
      RECT  0.08 1.325 0.2 1.43 ;
      RECT  3.69 1.325 3.84 1.44 ;
      RECT  3.69 1.44 5.935 1.56 ;
  END
END SEN_AOI32_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI32_8
#      Description : "One 3-input AND one 2-input AND into into 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|(B1&B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI32_8
  CLASS CORE ;
  FOREIGN SEN_AOI32_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.05 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.65 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.71 7.945 0.89 ;
      RECT  6.55 0.89 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.545 0.71 10.85 0.89 ;
      RECT  10.75 0.89 10.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 11.2 1.85 ;
      RECT  0.59 1.44 0.72 1.75 ;
      RECT  1.11 1.44 1.24 1.75 ;
      RECT  1.63 1.44 1.76 1.75 ;
      RECT  2.15 1.44 2.28 1.75 ;
      RECT  2.67 1.44 2.8 1.75 ;
      RECT  3.19 1.44 3.32 1.75 ;
      RECT  3.71 1.44 3.84 1.75 ;
      RECT  4.23 1.44 4.36 1.75 ;
      RECT  4.75 1.44 4.88 1.75 ;
      RECT  5.27 1.44 5.4 1.75 ;
      RECT  5.79 1.44 5.92 1.75 ;
      RECT  6.31 1.44 6.44 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.2 0.05 ;
      RECT  0.33 0.05 0.46 0.36 ;
      RECT  0.85 0.05 0.98 0.36 ;
      RECT  1.37 0.05 1.5 0.36 ;
      RECT  1.89 0.05 2.02 0.36 ;
      RECT  9.16 0.05 9.29 0.385 ;
      RECT  9.68 0.05 9.81 0.385 ;
      RECT  10.2 0.05 10.33 0.385 ;
      RECT  10.72 0.05 10.85 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.47 0.45 8.8 0.57 ;
      RECT  4.47 0.57 8.25 0.59 ;
      RECT  6.55 0.59 8.25 0.62 ;
      RECT  8.08 0.62 8.25 1.11 ;
      RECT  6.82 1.11 10.65 1.18 ;
      RECT  6.82 1.18 10.9 1.29 ;
    END
    ANTENNADIFFAREA 1.786 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.36 0.19 6.49 0.32 ;
      RECT  3.755 0.32 5.07 0.36 ;
      RECT  6.78 0.19 9.06 0.32 ;
      RECT  8.14 0.32 9.06 0.36 ;
      RECT  8.89 0.36 9.06 0.475 ;
      RECT  8.89 0.475 11.105 0.615 ;
      RECT  10.985 0.39 11.105 0.475 ;
      RECT  0.075 0.34 0.195 0.45 ;
      RECT  0.075 0.45 4.38 0.57 ;
      RECT  1.465 0.57 3.065 0.62 ;
      RECT  1.74 1.18 6.72 1.22 ;
      RECT  0.285 1.22 6.72 1.35 ;
      RECT  4.51 1.35 4.6 1.355 ;
      RECT  6.55 1.35 6.72 1.415 ;
      RECT  6.55 1.415 9.685 1.465 ;
      RECT  6.55 1.465 11.105 1.585 ;
      RECT  10.985 1.36 11.105 1.465 ;
  END
END SEN_AOI32_8
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI33_1
#      Description : "Two 3-input ANDs into a 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|(B1&B2&B3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI33_1
  CLASS CORE ;
  FOREIGN SEN_AOI33_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.755 ;
      RECT  0.69 0.755 0.85 0.925 ;
      RECT  0.75 0.925 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.755 ;
      RECT  0.35 0.755 0.51 0.925 ;
      RECT  0.35 0.925 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.755 ;
      RECT  1.15 0.755 1.28 0.925 ;
      RECT  1.15 0.925 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.575 1.415 0.705 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.06 0.05 0.185 0.39 ;
      RECT  1.62 0.05 1.745 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.785 0.24 1.46 0.36 ;
      RECT  1.35 0.36 1.46 0.69 ;
      RECT  1.37 0.69 1.46 1.0 ;
      RECT  1.35 1.0 1.46 1.23 ;
      RECT  1.05 1.23 1.745 1.35 ;
      RECT  1.63 1.35 1.745 1.61 ;
    END
    ANTENNADIFFAREA 0.297 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.265 1.205 0.96 1.325 ;
      RECT  0.84 1.325 0.96 1.44 ;
      RECT  0.84 1.44 1.535 1.56 ;
  END
END SEN_AOI33_1
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI33_2
#      Description : "Two 3-input ANDs into a 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|(B1&B2&B3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI33_2
  CLASS CORE ;
  FOREIGN SEN_AOI33_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.45 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.05 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.65 0.89 ;
      RECT  3.55 0.89 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.215 0.19 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.59 1.415 0.71 1.75 ;
      RECT  1.11 1.415 1.23 1.75 ;
      RECT  1.6 1.415 1.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.33 0.05 0.45 0.385 ;
      RECT  3.355 0.05 3.475 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.355 0.32 2.525 0.42 ;
      RECT  2.355 0.42 2.475 0.44 ;
      RECT  1.35 0.44 2.475 0.56 ;
      RECT  1.35 0.56 1.45 0.69 ;
      RECT  2.15 0.56 2.25 1.16 ;
      RECT  2.135 1.16 2.25 1.245 ;
      RECT  2.135 1.245 3.5 1.365 ;
    END
    ANTENNADIFFAREA 0.595 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.12 0.14 2.955 0.23 ;
      RECT  2.12 0.23 2.24 0.35 ;
      RECT  2.835 0.23 2.955 0.4 ;
      RECT  0.825 0.23 1.745 0.35 ;
      RECT  3.615 0.38 3.735 0.495 ;
      RECT  2.58 0.495 3.735 0.615 ;
      RECT  2.58 0.615 2.695 0.705 ;
      RECT  0.045 0.475 1.23 0.595 ;
      RECT  1.125 0.595 1.23 0.655 ;
      RECT  0.305 1.205 1.98 1.325 ;
      RECT  1.86 1.325 1.98 1.48 ;
      RECT  1.86 1.48 3.735 1.6 ;
      RECT  3.615 1.36 3.735 1.48 ;
  END
END SEN_AOI33_2
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI33_4
#      Description : "Two 3-input ANDs into a 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|(B1&B2&B3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI33_4
  CLASS CORE ;
  FOREIGN SEN_AOI33_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.85 0.89 ;
      RECT  6.75 0.89 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.585 1.415 0.715 1.75 ;
      RECT  1.105 1.415 1.235 1.75 ;
      RECT  1.625 1.415 1.755 1.75 ;
      RECT  2.145 1.415 2.275 1.75 ;
      RECT  2.655 1.415 2.785 1.75 ;
      RECT  3.175 1.415 3.305 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  0.325 0.05 0.455 0.385 ;
      RECT  0.845 0.05 0.975 0.385 ;
      RECT  6.025 0.05 6.155 0.385 ;
      RECT  6.545 0.05 6.675 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.36 0.47 4.64 0.59 ;
      RECT  4.35 0.59 4.45 1.11 ;
      RECT  3.95 1.11 5.455 1.18 ;
      RECT  3.65 1.18 6.66 1.29 ;
      RECT  5.75 1.11 6.66 1.18 ;
    END
    ANTENNADIFFAREA 1.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.32 0.235 3.355 0.355 ;
      RECT  3.645 0.24 5.655 0.36 ;
      RECT  0.07 0.37 0.19 0.475 ;
      RECT  0.07 0.475 2.27 0.595 ;
      RECT  2.15 0.595 2.27 0.675 ;
      RECT  6.81 0.365 6.93 0.475 ;
      RECT  4.73 0.475 6.93 0.595 ;
      RECT  4.73 0.595 4.85 0.67 ;
      RECT  0.28 1.205 3.56 1.325 ;
      RECT  3.44 1.325 3.56 1.44 ;
      RECT  3.44 1.44 6.93 1.56 ;
      RECT  6.81 1.335 6.93 1.44 ;
  END
END SEN_AOI33_4
#-----------------------------------------------------------------------
#      Cell        : SEN_AOI33_6
#      Description : "Two 3-input ANDs into a 2-input NOR"
#      Equation    : X=!((A1&A2&A3)|(B1&B2&B3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_AOI33_6
  CLASS CORE ;
  FOREIGN SEN_AOI33_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.65 0.89 ;
      RECT  4.55 0.89 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.71 6.28 0.89 ;
      RECT  5.35 0.89 5.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 8.05 0.89 ;
      RECT  7.95 0.89 8.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.95 0.71 10.05 0.89 ;
      RECT  9.95 0.89 10.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 10.2 1.85 ;
      RECT  0.59 1.415 0.72 1.75 ;
      RECT  1.11 1.415 1.24 1.75 ;
      RECT  1.63 1.415 1.76 1.75 ;
      RECT  2.15 1.415 2.28 1.75 ;
      RECT  2.67 1.415 2.8 1.75 ;
      RECT  3.19 1.415 3.32 1.75 ;
      RECT  3.715 1.415 3.845 1.75 ;
      RECT  4.235 1.415 4.365 1.75 ;
      RECT  4.755 1.415 4.885 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      RECT  8.655 0.05 8.785 0.375 ;
      RECT  9.175 0.05 9.305 0.375 ;
      RECT  9.695 0.05 9.825 0.375 ;
      RECT  0.33 0.05 0.46 0.385 ;
      RECT  0.85 0.05 0.98 0.385 ;
      RECT  1.37 0.05 1.5 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.435 0.46 6.725 0.595 ;
      RECT  6.52 0.595 6.65 1.11 ;
      RECT  5.55 1.11 7.855 1.18 ;
      RECT  5.55 1.18 9.85 1.19 ;
      RECT  8.15 1.11 9.85 1.18 ;
      RECT  5.235 1.19 9.85 1.31 ;
    END
    ANTENNADIFFAREA 1.714 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.84 0.23 4.935 0.36 ;
      RECT  5.225 0.23 8.315 0.36 ;
      RECT  9.96 0.37 10.08 0.465 ;
      RECT  6.815 0.465 10.08 0.595 ;
      RECT  0.075 0.38 0.195 0.475 ;
      RECT  0.075 0.475 3.34 0.605 ;
      RECT  0.285 1.195 5.145 1.325 ;
      RECT  5.015 1.325 5.145 1.435 ;
      RECT  5.015 1.435 10.08 1.565 ;
      RECT  9.96 1.335 10.08 1.435 ;
  END
END SEN_AOI33_6
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_1
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_1
  CLASS CORE ;
  FOREIGN SEN_BUF_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.655 0.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.44 0.46 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.335 0.05 0.46 0.375 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.73 0.69 ;
      RECT  0.64 0.69 0.73 1.075 ;
      RECT  0.55 1.075 0.73 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.17 0.185 0.465 ;
      RECT  0.07 0.465 0.445 0.555 ;
      RECT  0.355 0.555 0.445 0.79 ;
      RECT  0.355 0.79 0.55 0.89 ;
      RECT  0.355 0.89 0.445 1.26 ;
      RECT  0.07 1.26 0.445 1.35 ;
      RECT  0.07 1.35 0.19 1.6 ;
  END
END SEN_BUF_1
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_12
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_12
  CLASS CORE ;
  FOREIGN SEN_BUF_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.18 1.41 3.31 1.75 ;
      RECT  3.7 1.41 3.83 1.75 ;
      RECT  4.22 1.41 4.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  1.62 0.05 1.75 0.39 ;
      RECT  2.145 0.05 2.27 0.39 ;
      RECT  2.66 0.05 2.79 0.39 ;
      RECT  3.18 0.05 3.31 0.39 ;
      RECT  3.7 0.05 3.83 0.39 ;
      RECT  4.22 0.05 4.345 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.34 0.51 4.25 0.69 ;
      RECT  3.4 0.69 3.65 1.11 ;
      RECT  1.34 1.11 4.25 1.29 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.3 0.48 1.045 0.59 ;
      RECT  0.955 0.59 1.045 0.79 ;
      RECT  0.955 0.79 3.29 0.89 ;
      RECT  0.955 0.89 1.045 1.21 ;
      RECT  0.3 1.21 1.045 1.32 ;
  END
END SEN_BUF_12
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_16
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_16
  CLASS CORE ;
  FOREIGN SEN_BUF_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.25 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3456 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.595 1.42 0.725 1.75 ;
      RECT  1.115 1.42 1.245 1.75 ;
      RECT  1.64 1.21 1.76 1.75 ;
      RECT  2.16 1.435 2.28 1.75 ;
      RECT  2.675 1.41 2.805 1.75 ;
      RECT  3.195 1.41 3.325 1.75 ;
      RECT  3.715 1.41 3.845 1.75 ;
      RECT  4.235 1.41 4.365 1.75 ;
      RECT  4.755 1.41 4.885 1.75 ;
      RECT  5.275 1.41 5.405 1.75 ;
      RECT  5.815 1.21 5.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  4.235 0.05 4.365 0.37 ;
      RECT  4.755 0.05 4.885 0.37 ;
      RECT  0.595 0.05 0.725 0.38 ;
      RECT  1.115 0.05 1.245 0.38 ;
      RECT  2.155 0.05 2.285 0.39 ;
      RECT  2.675 0.05 2.805 0.39 ;
      RECT  3.195 0.05 3.325 0.39 ;
      RECT  3.715 0.05 3.87 0.39 ;
      RECT  5.275 0.05 5.405 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.64 0.05 1.76 0.59 ;
      RECT  5.815 0.05 5.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.04 0.46 4.85 0.51 ;
      RECT  1.865 0.51 5.685 0.69 ;
      RECT  4.53 0.69 4.85 1.07 ;
      RECT  1.865 1.07 4.85 1.11 ;
      RECT  1.865 1.11 5.685 1.29 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.31 0.47 1.525 0.59 ;
      RECT  1.395 0.59 1.525 0.78 ;
      RECT  1.395 0.78 4.42 0.91 ;
      RECT  1.395 0.91 1.525 1.21 ;
      RECT  0.315 1.21 1.525 1.33 ;
  END
END SEN_BUF_16
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_2
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_2
  CLASS CORE ;
  FOREIGN SEN_BUF_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0432 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.345 1.575 0.515 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.96 1.21 1.08 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.365 0.05 0.495 0.39 ;
      RECT  0.96 0.05 1.08 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.85 0.69 ;
      RECT  0.75 0.69 0.85 1.11 ;
      RECT  0.55 1.11 0.85 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.29 0.19 0.5 ;
      RECT  0.07 0.5 0.45 0.59 ;
      RECT  0.36 0.59 0.45 0.785 ;
      RECT  0.36 0.785 0.66 0.895 ;
      RECT  0.36 0.895 0.45 1.395 ;
      RECT  0.07 1.395 0.45 1.485 ;
      RECT  0.07 1.485 0.2 1.62 ;
  END
END SEN_BUF_2
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_24
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_24
  CLASS CORE ;
  FOREIGN SEN_BUF_24 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.595 1.43 0.725 1.75 ;
      RECT  1.115 1.43 1.245 1.75 ;
      RECT  1.635 1.43 1.77 1.75 ;
      RECT  2.155 1.41 2.285 1.75 ;
      RECT  2.675 1.435 2.805 1.75 ;
      RECT  3.195 1.435 3.325 1.75 ;
      RECT  3.715 1.435 3.845 1.75 ;
      RECT  4.235 1.435 4.365 1.75 ;
      RECT  4.755 1.435 4.885 1.75 ;
      RECT  5.275 1.435 5.405 1.75 ;
      RECT  5.795 1.435 5.925 1.75 ;
      RECT  6.315 1.435 6.445 1.75 ;
      RECT  6.835 1.435 6.965 1.75 ;
      RECT  7.355 1.435 7.485 1.75 ;
      RECT  7.875 1.435 8.005 1.75 ;
      RECT  8.41 1.21 8.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  5.255 0.05 5.425 0.325 ;
      RECT  5.775 0.05 5.945 0.325 ;
      RECT  4.755 0.05 4.885 0.355 ;
      RECT  0.595 0.05 0.725 0.37 ;
      RECT  1.115 0.05 1.245 0.37 ;
      RECT  1.635 0.05 1.765 0.37 ;
      RECT  2.675 0.05 2.805 0.37 ;
      RECT  3.195 0.05 3.325 0.37 ;
      RECT  3.715 0.05 3.845 0.37 ;
      RECT  4.24 0.05 4.36 0.37 ;
      RECT  6.315 0.05 6.445 0.375 ;
      RECT  6.835 0.05 6.965 0.375 ;
      RECT  7.355 0.05 7.485 0.375 ;
      RECT  7.875 0.05 8.005 0.375 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  2.16 0.05 2.28 0.59 ;
      RECT  8.41 0.05 8.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.055 0.415 6.06 0.445 ;
      RECT  4.505 0.445 6.06 0.495 ;
      RECT  2.395 0.495 8.29 0.64 ;
      RECT  2.395 0.64 7.45 0.665 ;
      RECT  5.55 0.665 7.45 0.69 ;
      RECT  5.55 0.69 6.05 1.055 ;
      RECT  5.015 1.055 6.05 1.085 ;
      RECT  2.35 1.085 6.05 1.11 ;
      RECT  2.35 1.11 8.285 1.305 ;
    END
    ANTENNADIFFAREA 2.592 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.31 0.46 2.05 0.59 ;
      RECT  1.87 0.59 2.05 0.75 ;
      RECT  1.87 0.75 2.3 0.775 ;
      RECT  1.87 0.775 5.44 0.895 ;
      RECT  1.87 0.895 2.05 1.21 ;
      RECT  0.315 1.21 2.05 1.34 ;
      RECT  7.575 0.75 8.13 0.785 ;
      RECT  6.16 0.785 8.13 0.895 ;
      LAYER M2 ;
      RECT  1.91 0.75 8.115 0.85 ;
      LAYER V1 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  7.645 0.75 7.745 0.85 ;
      RECT  7.975 0.75 8.075 0.85 ;
  END
END SEN_BUF_24
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_3
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_3
  CLASS CORE ;
  FOREIGN SEN_BUF_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.175 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.395 1.455 0.525 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.94 1.41 1.07 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.945 0.05 1.075 0.375 ;
      RECT  0.395 0.05 0.525 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.22 0.37 1.335 0.48 ;
      RECT  0.95 0.48 1.335 0.51 ;
      RECT  0.55 0.51 1.335 0.59 ;
      RECT  0.55 0.59 1.05 0.69 ;
      RECT  0.95 0.69 1.05 1.11 ;
      RECT  0.55 1.11 1.335 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.125 0.37 0.235 0.49 ;
      RECT  0.125 0.49 0.44 0.59 ;
      RECT  0.35 0.59 0.44 0.785 ;
      RECT  0.35 0.785 0.86 0.895 ;
      RECT  0.35 0.895 0.44 1.265 ;
      RECT  0.12 1.265 0.44 1.365 ;
      RECT  0.12 1.365 0.24 1.5 ;
  END
END SEN_BUF_3
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_4
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_4
  CLASS CORE ;
  FOREIGN SEN_BUF_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0864 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.58 1.425 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.56 0.05 0.73 0.305 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  1.625 0.05 1.745 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.82 0.51 1.65 0.69 ;
      RECT  1.35 0.69 1.45 1.105 ;
      RECT  0.75 1.105 1.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.3 0.41 0.645 0.515 ;
      RECT  0.555 0.515 0.645 0.785 ;
      RECT  0.555 0.785 1.24 0.895 ;
      RECT  0.555 0.895 0.645 1.215 ;
      RECT  0.3 1.215 0.645 1.335 ;
  END
END SEN_BUF_4
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_6
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_6
  CLASS CORE ;
  FOREIGN SEN_BUF_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      RECT  1.115 1.415 1.245 1.75 ;
      RECT  1.635 1.41 1.765 1.75 ;
      RECT  2.18 1.21 2.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      RECT  1.115 0.05 1.245 0.39 ;
      RECT  1.635 0.05 1.765 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  2.18 0.05 2.3 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 2.05 0.69 ;
      RECT  1.92 0.69 2.05 1.11 ;
      RECT  0.75 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.315 0.48 0.645 0.59 ;
      RECT  0.55 0.59 0.645 0.79 ;
      RECT  0.55 0.79 1.81 0.9 ;
      RECT  0.55 0.9 0.645 1.21 ;
      RECT  0.315 1.21 0.645 1.32 ;
  END
END SEN_BUF_6
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_8
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_8
  CLASS CORE ;
  FOREIGN SEN_BUF_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1728 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.36 1.41 1.49 1.75 ;
      RECT  1.895 1.41 2.025 1.75 ;
      RECT  2.45 1.41 2.58 1.75 ;
      RECT  3.01 1.21 3.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      RECT  1.895 0.05 2.025 0.39 ;
      RECT  2.455 0.05 2.585 0.39 ;
      RECT  3.01 0.05 3.13 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 2.88 0.69 ;
      RECT  2.28 0.69 2.45 1.105 ;
      RECT  0.95 1.105 2.88 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 0.845 0.59 ;
      RECT  0.75 0.59 0.845 0.79 ;
      RECT  0.75 0.79 2.17 0.89 ;
      RECT  0.75 0.89 0.845 1.21 ;
      RECT  0.065 1.21 0.845 1.31 ;
      RECT  0.065 1.31 0.185 1.43 ;
  END
END SEN_BUF_8
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_0P5
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_0P5
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.275 0.185 0.71 ;
      RECT  0.065 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNADIFFAREA 0.06 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.55 1.44 0.66 1.75 ;
      RECT  0.0 1.75 1.0 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      RECT  0.55 0.05 0.68 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.825 0.18 0.935 0.71 ;
      RECT  0.75 0.71 0.935 0.8 ;
      RECT  0.75 0.8 0.85 1.31 ;
      RECT  0.75 1.31 0.935 1.49 ;
    END
    ANTENNADIFFAREA 0.076 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.295 0.18 0.415 0.45 ;
      RECT  0.295 0.45 0.735 0.54 ;
      RECT  0.555 0.54 0.735 0.62 ;
      RECT  0.555 0.62 0.66 1.26 ;
      RECT  0.295 1.26 0.66 1.35 ;
      RECT  0.295 1.35 0.415 1.63 ;
  END
END SEN_BUF_AS_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_1
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_1
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.835 ;
      RECT  0.15 0.835 0.475 0.95 ;
      RECT  0.15 0.95 0.25 1.09 ;
    END
    ANTENNADIFFAREA 0.096 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0327 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.485 1.415 0.615 1.75 ;
      RECT  0.0 1.75 1.0 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      RECT  0.55 0.05 0.66 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.205 0.935 0.49 ;
      RECT  0.835 0.49 0.935 1.04 ;
      RECT  0.75 1.04 0.935 1.49 ;
    END
    ANTENNADIFFAREA 0.146 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.295 0.2 0.43 0.4 ;
      RECT  0.34 0.4 0.43 0.54 ;
      RECT  0.34 0.54 0.66 0.63 ;
      RECT  0.565 0.63 0.66 0.675 ;
      RECT  0.565 0.675 0.745 0.845 ;
      RECT  0.565 0.845 0.66 1.21 ;
      RECT  0.145 1.21 0.66 1.3 ;
      RECT  0.145 1.3 0.265 1.49 ;
  END
END SEN_BUF_AS_1
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_10
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_10
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.09 0.27 0.25 0.71 ;
      RECT  0.09 0.71 1.25 0.89 ;
    END
    ANTENNADIFFAREA 0.06 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.48 1.25 0.6 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  1.08 1.25 1.2 1.75 ;
      RECT  1.64 1.21 1.76 1.75 ;
      RECT  2.16 1.21 2.28 1.75 ;
      RECT  2.68 1.21 2.8 1.75 ;
      RECT  3.2 1.215 3.32 1.75 ;
      RECT  3.72 1.21 3.84 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  2.155 0.05 2.285 0.345 ;
      RECT  2.675 0.05 2.805 0.345 ;
      RECT  3.195 0.05 3.325 0.345 ;
      RECT  3.715 0.05 3.845 0.345 ;
      RECT  0.595 0.05 0.725 0.35 ;
      RECT  1.115 0.05 1.245 0.35 ;
      RECT  1.64 0.05 1.76 0.57 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.29 4.1 0.435 ;
      RECT  1.85 0.435 4.1 0.565 ;
      RECT  3.44 0.565 3.65 0.91 ;
      RECT  1.9 0.91 4.1 1.09 ;
      RECT  1.9 1.09 2.05 1.29 ;
      RECT  3.95 1.09 4.1 1.29 ;
    END
    ANTENNADIFFAREA 0.991 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.34 0.46 0.44 ;
      RECT  0.34 0.44 1.55 0.56 ;
      RECT  1.44 0.56 1.55 0.685 ;
      RECT  1.44 0.685 3.35 0.795 ;
      RECT  1.44 0.795 1.55 1.04 ;
      RECT  0.13 1.04 1.55 1.16 ;
  END
END SEN_BUF_AS_10
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_12
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_12
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.12 0.31 0.25 0.71 ;
      RECT  0.12 0.71 1.45 0.89 ;
    END
    ANTENNADIFFAREA 0.099 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3933 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.41 0.505 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.975 1.41 1.105 1.75 ;
      RECT  1.575 1.41 1.705 1.75 ;
      RECT  2.16 1.21 2.28 1.75 ;
      RECT  2.7 1.21 2.82 1.75 ;
      RECT  3.22 1.21 3.34 1.75 ;
      RECT  3.74 1.21 3.86 1.75 ;
      RECT  4.26 1.21 4.38 1.75 ;
      RECT  4.79 1.21 4.91 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  2.415 0.05 2.585 0.315 ;
      RECT  2.935 0.05 3.105 0.315 ;
      RECT  3.455 0.05 3.625 0.315 ;
      RECT  3.975 0.05 4.145 0.315 ;
      RECT  4.495 0.05 4.68 0.315 ;
      RECT  0.875 0.05 1.005 0.38 ;
      RECT  1.395 0.05 1.525 0.38 ;
      RECT  1.92 0.05 2.04 0.545 ;
      RECT  0.36 0.05 0.48 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.155 0.405 4.925 0.53 ;
      RECT  4.0 0.53 4.925 0.54 ;
      RECT  4.0 0.54 4.25 0.91 ;
      RECT  2.35 0.91 4.65 1.09 ;
      RECT  4.52 1.09 4.65 1.29 ;
    END
    ANTENNADIFFAREA 1.113 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.66 0.36 1.78 0.47 ;
      RECT  0.595 0.47 1.78 0.59 ;
      RECT  1.65 0.59 1.78 0.635 ;
      RECT  1.65 0.635 3.89 0.765 ;
      RECT  1.65 0.765 1.78 1.21 ;
      RECT  0.08 1.21 2.035 1.32 ;
      RECT  0.08 1.32 0.2 1.43 ;
  END
END SEN_BUF_AS_12
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_16
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_16
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.205 0.255 0.71 ;
      RECT  0.15 0.71 1.65 0.89 ;
    END
    ANTENNADIFFAREA 0.108 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5244 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.385 1.43 0.515 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.935 1.43 1.065 1.75 ;
      RECT  1.485 1.43 1.615 1.75 ;
      RECT  2.025 1.43 2.165 1.75 ;
      RECT  2.575 1.21 2.695 1.75 ;
      RECT  3.095 1.21 3.215 1.75 ;
      RECT  3.615 1.21 3.735 1.75 ;
      RECT  4.135 1.21 4.255 1.75 ;
      RECT  4.655 1.21 4.775 1.75 ;
      RECT  5.175 1.21 5.295 1.75 ;
      RECT  5.695 1.21 5.815 1.75 ;
      RECT  6.215 1.21 6.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  3.59 0.05 3.76 0.31 ;
      RECT  4.11 0.05 4.28 0.31 ;
      RECT  4.63 0.05 4.8 0.31 ;
      RECT  5.15 0.05 5.32 0.31 ;
      RECT  5.67 0.05 5.84 0.31 ;
      RECT  3.07 0.05 3.24 0.315 ;
      RECT  1.52 0.05 1.65 0.35 ;
      RECT  2.045 0.05 2.175 0.35 ;
      RECT  1.0 0.05 1.13 0.355 ;
      RECT  2.575 0.05 2.695 0.545 ;
      RECT  0.465 0.05 0.585 0.59 ;
      RECT  6.22 0.05 6.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.81 0.41 6.1 0.53 ;
      RECT  2.81 0.53 5.25 0.545 ;
      RECT  4.93 0.545 5.25 0.91 ;
      RECT  2.75 0.91 6.075 1.1 ;
      RECT  5.95 1.1 6.075 1.29 ;
    END
    ANTENNADIFFAREA 1.466 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.72 0.46 2.46 0.59 ;
      RECT  2.275 0.59 2.46 0.635 ;
      RECT  2.275 0.635 4.82 0.82 ;
      RECT  2.275 0.82 2.46 1.115 ;
      RECT  0.09 1.115 2.46 1.285 ;
  END
END SEN_BUF_AS_16
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_1P5
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_1P5
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.275 0.185 0.71 ;
      RECT  0.065 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNADIFFAREA 0.06 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0498 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.49 1.4 0.62 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.16 1.21 1.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.57 0.05 0.7 0.39 ;
      RECT  1.11 0.05 1.24 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.845 0.21 0.955 0.47 ;
      RECT  0.845 0.47 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.31 ;
      RECT  0.75 1.31 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.138 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.315 0.3 0.435 0.48 ;
      RECT  0.315 0.48 0.65 0.57 ;
      RECT  0.55 0.57 0.65 0.745 ;
      RECT  0.55 0.745 0.86 0.855 ;
      RECT  0.55 0.855 0.65 1.22 ;
      RECT  0.155 1.22 0.65 1.31 ;
      RECT  0.155 1.31 0.275 1.46 ;
  END
END SEN_BUF_AS_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_2
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_2
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.24 0.25 0.91 ;
      RECT  0.15 0.91 0.65 1.09 ;
    END
    ANTENNADIFFAREA 0.108 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0654 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.1 1.36 0.225 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.65 1.41 0.78 1.75 ;
      RECT  1.215 1.21 1.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.21 0.05 1.34 0.39 ;
      RECT  0.665 0.05 0.785 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.295 1.055 0.5 ;
      RECT  0.94 0.5 1.25 0.59 ;
      RECT  1.15 0.59 1.25 1.01 ;
      RECT  0.95 1.01 1.25 1.11 ;
      RECT  0.95 1.11 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.4 0.38 0.525 0.71 ;
      RECT  0.4 0.71 1.04 0.8 ;
      RECT  0.75 0.8 1.04 0.82 ;
      RECT  0.75 0.82 0.86 1.21 ;
      RECT  0.37 1.21 0.86 1.31 ;
      RECT  0.37 1.31 0.5 1.49 ;
  END
END SEN_BUF_AS_2
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_3
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_3
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.12 0.205 0.26 0.71 ;
      RECT  0.12 0.71 0.48 0.89 ;
    END
    ANTENNADIFFAREA 0.099 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0978 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.62 1.21 0.74 1.75 ;
      RECT  1.135 1.41 1.265 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.355 0.05 0.485 0.39 ;
      RECT  0.875 0.05 1.005 0.39 ;
      RECT  1.415 0.05 1.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.3 1.25 1.11 ;
      RECT  0.875 1.11 1.525 1.29 ;
    END
    ANTENNADIFFAREA 0.313 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.625 0.27 0.735 0.785 ;
      RECT  0.625 0.785 1.06 0.895 ;
      RECT  0.625 0.895 0.735 1.01 ;
      RECT  0.36 1.01 0.735 1.11 ;
      RECT  0.36 1.11 0.47 1.32 ;
  END
END SEN_BUF_AS_3
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_4
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_4
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.24 0.25 0.71 ;
      RECT  0.15 0.71 0.735 0.89 ;
    END
    ANTENNADIFFAREA 0.108 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1311 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.38 1.21 0.5 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  0.9 1.21 1.02 1.75 ;
      RECT  1.415 1.41 1.545 1.75 ;
      RECT  1.96 1.21 2.08 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  1.63 0.05 1.79 0.37 ;
      RECT  0.42 0.05 0.545 0.59 ;
      RECT  1.045 0.05 1.165 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.33 0.475 2.085 0.575 ;
      RECT  1.75 0.575 1.85 1.11 ;
      RECT  1.15 1.11 1.85 1.29 ;
    END
    ANTENNADIFFAREA 0.4 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.665 0.34 0.955 0.455 ;
      RECT  0.845 0.455 0.955 0.755 ;
      RECT  0.845 0.755 1.64 0.86 ;
      RECT  0.845 0.86 0.955 1.01 ;
      RECT  0.11 1.01 0.955 1.11 ;
      RECT  0.11 1.11 0.23 1.38 ;
      RECT  0.64 1.11 0.76 1.38 ;
  END
END SEN_BUF_AS_4
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_5
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_5
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.27 0.25 0.71 ;
      RECT  0.08 0.71 1.05 0.89 ;
    END
    ANTENNADIFFAREA 0.06 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1665 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.445 1.295 0.615 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.005 1.295 1.175 1.75 ;
      RECT  1.625 1.41 1.755 1.75 ;
      RECT  2.145 1.41 2.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.625 0.05 1.755 0.345 ;
      RECT  2.235 0.05 2.365 0.345 ;
      RECT  0.585 0.05 0.715 0.35 ;
      RECT  1.105 0.05 1.235 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.345 0.435 2.45 0.565 ;
      RECT  2.35 0.565 2.45 1.11 ;
      RECT  1.35 1.11 2.53 1.29 ;
    END
    ANTENNADIFFAREA 0.5 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.37 0.45 0.44 ;
      RECT  0.34 0.44 1.25 0.56 ;
      RECT  1.14 0.56 1.25 0.755 ;
      RECT  1.14 0.755 2.14 0.865 ;
      RECT  1.14 0.865 1.25 1.09 ;
      RECT  0.145 1.09 1.25 1.205 ;
  END
END SEN_BUF_AS_5
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_6
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_6
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.105 0.17 0.25 0.71 ;
      RECT  0.105 0.71 0.68 0.89 ;
    END
    ANTENNADIFFAREA 0.082 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.215 0.455 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.865 1.21 0.985 1.75 ;
      RECT  1.38 1.41 1.51 1.75 ;
      RECT  1.9 1.41 2.03 1.75 ;
      RECT  2.42 1.41 2.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.345 0.05 0.485 0.39 ;
      RECT  0.86 0.05 0.99 0.39 ;
      RECT  1.9 0.05 2.03 0.39 ;
      RECT  2.42 0.05 2.545 0.39 ;
      RECT  1.385 0.05 1.505 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.62 0.51 2.45 0.69 ;
      RECT  1.92 0.69 2.05 1.11 ;
      RECT  1.13 1.11 2.45 1.29 ;
    END
    ANTENNADIFFAREA 0.548 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.605 0.24 0.72 0.51 ;
      RECT  0.605 0.51 1.24 0.62 ;
      RECT  1.135 0.29 1.24 0.51 ;
      RECT  1.12 0.62 1.24 0.8 ;
      RECT  1.12 0.8 1.81 0.81 ;
      RECT  0.925 0.81 1.81 0.92 ;
      RECT  0.925 0.92 1.04 1.01 ;
      RECT  0.065 1.01 1.04 1.12 ;
      RECT  0.065 1.12 0.185 1.23 ;
  END
END SEN_BUF_AS_6
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_AS_8
#      Description : "Symmetric rise/fall time buffer, antenna diode on input"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_AS_8
  CLASS CORE ;
  FOREIGN SEN_BUF_AS_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.24 0.25 0.71 ;
      RECT  0.15 0.71 1.41 0.89 ;
    END
    ANTENNADIFFAREA 0.156 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2619 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.45 1.255 0.565 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  1.005 1.255 1.12 1.75 ;
      RECT  1.525 1.255 1.64 1.75 ;
      RECT  2.035 1.415 2.165 1.75 ;
      RECT  2.555 1.415 2.685 1.75 ;
      RECT  3.075 1.415 3.205 1.75 ;
      RECT  3.615 1.21 3.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  2.555 0.05 2.685 0.37 ;
      RECT  3.075 0.05 3.205 0.37 ;
      RECT  0.475 0.05 0.605 0.39 ;
      RECT  0.985 0.05 1.125 0.39 ;
      RECT  1.515 0.05 1.645 0.39 ;
      RECT  2.035 0.05 2.165 0.39 ;
      RECT  3.615 0.05 3.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.275 0.46 3.505 0.57 ;
      RECT  3.08 0.57 3.505 0.575 ;
      RECT  3.08 0.575 3.25 1.11 ;
      RECT  1.75 1.11 3.46 1.29 ;
    END
    ANTENNADIFFAREA 0.732 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.74 0.24 0.86 0.5 ;
      RECT  0.74 0.5 1.61 0.59 ;
      RECT  1.265 0.24 1.375 0.5 ;
      RECT  1.52 0.59 1.61 0.755 ;
      RECT  1.52 0.755 2.98 0.865 ;
      RECT  1.79 0.24 1.895 0.755 ;
      RECT  1.52 0.865 1.61 1.055 ;
      RECT  0.15 1.055 1.61 1.165 ;
      RECT  0.15 1.165 0.27 1.29 ;
  END
END SEN_BUF_AS_8
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_D_1
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_D_1
  CLASS CORE ;
  FOREIGN SEN_BUF_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.635 0.25 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.32 0.05 0.45 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.69 0.49 ;
      RECT  0.6 0.49 0.69 1.11 ;
      RECT  0.55 1.11 0.69 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.2 0.185 0.455 ;
      RECT  0.065 0.455 0.445 0.545 ;
      RECT  0.355 0.545 0.445 0.755 ;
      RECT  0.355 0.755 0.51 0.925 ;
      RECT  0.355 0.925 0.445 1.26 ;
      RECT  0.065 1.26 0.445 1.35 ;
      RECT  0.065 1.35 0.185 1.61 ;
  END
END SEN_BUF_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_D_12
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_D_12
  CLASS CORE ;
  FOREIGN SEN_BUF_D_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  1.36 1.41 1.49 1.75 ;
      RECT  1.88 1.41 2.01 1.75 ;
      RECT  2.4 1.41 2.53 1.75 ;
      RECT  2.92 1.41 3.05 1.75 ;
      RECT  3.44 1.41 3.57 1.75 ;
      RECT  3.98 1.21 4.1 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  1.34 0.05 1.51 0.325 ;
      RECT  1.86 0.05 2.03 0.325 ;
      RECT  2.38 0.05 2.55 0.325 ;
      RECT  2.9 0.05 3.07 0.325 ;
      RECT  3.42 0.05 3.59 0.325 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  3.98 0.05 4.1 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.065 0.415 3.875 0.535 ;
      RECT  1.95 0.535 3.25 0.585 ;
      RECT  3.0 0.585 3.25 1.11 ;
      RECT  1.055 1.11 3.85 1.29 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.38 0.185 0.475 ;
      RECT  0.065 0.475 0.965 0.595 ;
      RECT  0.86 0.595 0.965 0.77 ;
      RECT  0.86 0.77 2.91 0.895 ;
      RECT  0.86 0.895 0.965 1.205 ;
      RECT  0.065 1.205 0.965 1.325 ;
      RECT  0.065 1.325 0.185 1.425 ;
  END
END SEN_BUF_D_12
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_D_16
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_D_16
  CLASS CORE ;
  FOREIGN SEN_BUF_D_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.58 1.435 0.71 1.75 ;
      RECT  1.105 1.21 1.225 1.75 ;
      RECT  1.62 1.44 1.75 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  2.66 1.44 2.79 1.75 ;
      RECT  3.18 1.44 3.31 1.75 ;
      RECT  3.7 1.44 3.83 1.75 ;
      RECT  4.22 1.44 4.35 1.75 ;
      RECT  4.74 1.41 4.87 1.75 ;
      RECT  5.295 1.21 5.415 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  1.6 0.05 1.77 0.325 ;
      RECT  2.12 0.05 2.29 0.325 ;
      RECT  2.64 0.05 2.81 0.325 ;
      RECT  3.16 0.05 3.33 0.325 ;
      RECT  3.68 0.05 3.85 0.325 ;
      RECT  4.2 0.05 4.37 0.325 ;
      RECT  4.72 0.05 4.89 0.325 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.105 0.05 1.225 0.59 ;
      RECT  5.3 0.05 5.42 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.32 0.415 5.175 0.535 ;
      RECT  2.35 0.535 4.25 0.585 ;
      RECT  3.425 0.585 4.25 0.635 ;
      RECT  3.93 0.635 4.25 1.11 ;
      RECT  2.35 1.11 5.15 1.23 ;
      RECT  1.315 1.23 5.15 1.29 ;
      RECT  1.315 1.29 4.21 1.35 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.3 0.48 0.99 0.59 ;
      RECT  0.9 0.59 0.99 0.77 ;
      RECT  0.9 0.77 3.76 0.895 ;
      RECT  0.9 0.895 0.99 1.23 ;
      RECT  0.3 1.23 0.99 1.345 ;
  END
END SEN_BUF_D_16
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_D_2
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_D_2
  CLASS CORE ;
  FOREIGN SEN_BUF_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.64 0.25 1.175 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.445 0.45 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.865 1.41 0.995 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.32 0.05 0.45 0.365 ;
      RECT  0.865 0.05 0.995 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.56 0.475 0.85 0.595 ;
      RECT  0.75 0.595 0.85 1.11 ;
      RECT  0.55 1.11 0.85 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.21 0.185 0.455 ;
      RECT  0.065 0.455 0.445 0.545 ;
      RECT  0.35 0.545 0.445 0.785 ;
      RECT  0.35 0.785 0.66 0.895 ;
      RECT  0.35 0.895 0.45 1.265 ;
      RECT  0.065 1.265 0.45 1.355 ;
      RECT  0.065 1.355 0.185 1.53 ;
  END
END SEN_BUF_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_D_3
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_D_3
  CLASS CORE ;
  FOREIGN SEN_BUF_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.635 0.25 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.32 0.05 0.45 0.365 ;
      RECT  0.84 0.05 0.97 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.535 0.455 1.275 0.575 ;
      RECT  0.95 0.575 1.05 1.11 ;
      RECT  0.55 1.11 1.25 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.32 0.185 0.455 ;
      RECT  0.065 0.455 0.445 0.545 ;
      RECT  0.355 0.545 0.445 0.795 ;
      RECT  0.355 0.795 0.86 0.885 ;
      RECT  0.355 0.885 0.445 1.26 ;
      RECT  0.065 1.26 0.445 1.35 ;
      RECT  0.065 1.35 0.185 1.48 ;
  END
END SEN_BUF_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_D_4
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_D_4
  CLASS CORE ;
  FOREIGN SEN_BUF_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.635 0.25 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.38 1.21 1.5 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.32 0.05 0.45 0.365 ;
      RECT  0.84 0.05 0.97 0.365 ;
      RECT  1.38 0.05 1.5 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.455 1.275 0.575 ;
      RECT  0.95 0.575 1.05 1.11 ;
      RECT  0.55 1.11 1.25 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.325 0.185 0.455 ;
      RECT  0.065 0.455 0.445 0.545 ;
      RECT  0.355 0.545 0.445 0.795 ;
      RECT  0.355 0.795 0.86 0.885 ;
      RECT  0.355 0.885 0.445 1.26 ;
      RECT  0.065 1.26 0.445 1.35 ;
      RECT  0.065 1.35 0.185 1.48 ;
  END
END SEN_BUF_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_D_6
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_D_6
  CLASS CORE ;
  FOREIGN SEN_BUF_D_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.18 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.16 1.21 2.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  1.62 0.05 1.75 0.39 ;
      RECT  2.16 0.05 2.28 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.82 0.51 2.05 0.69 ;
      RECT  1.92 0.69 2.05 1.11 ;
      RECT  0.845 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.325 0.32 0.445 0.48 ;
      RECT  0.325 0.48 0.645 0.59 ;
      RECT  0.555 0.59 0.645 0.785 ;
      RECT  0.555 0.785 1.83 0.895 ;
      RECT  0.555 0.895 0.645 1.225 ;
      RECT  0.275 1.225 0.645 1.345 ;
  END
END SEN_BUF_D_6
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_D_8
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_D_8
  CLASS CORE ;
  FOREIGN SEN_BUF_D_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.58 1.42 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.69 1.21 2.81 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  0.58 0.05 0.71 0.38 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  1.62 0.05 1.75 0.39 ;
      RECT  2.14 0.05 2.27 0.39 ;
      RECT  0.07 0.05 0.18 0.59 ;
      RECT  2.69 0.05 2.81 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.82 0.51 2.55 0.69 ;
      RECT  2.28 0.69 2.45 1.11 ;
      RECT  0.845 1.11 2.53 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.47 0.645 0.59 ;
      RECT  0.555 0.59 0.645 0.785 ;
      RECT  0.555 0.785 2.17 0.895 ;
      RECT  0.555 0.895 0.645 1.21 ;
      RECT  0.28 1.21 0.645 1.33 ;
  END
END SEN_BUF_D_8
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_S_1
#      Description : "Symmetric rise/fall delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_S_1
  CLASS CORE ;
  FOREIGN SEN_BUF_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.655 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0327 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.41 0.46 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.335 0.05 0.46 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.735 0.69 ;
      RECT  0.645 0.69 0.735 1.07 ;
      RECT  0.55 1.07 0.735 1.25 ;
      RECT  0.55 1.25 0.65 1.49 ;
    END
    ANTENNADIFFAREA 0.146 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.19 0.19 0.475 ;
      RECT  0.07 0.475 0.445 0.565 ;
      RECT  0.355 0.565 0.445 0.78 ;
      RECT  0.355 0.78 0.555 0.95 ;
      RECT  0.355 0.95 0.445 1.21 ;
      RECT  0.07 1.21 0.445 1.3 ;
      RECT  0.07 1.3 0.19 1.49 ;
  END
END SEN_BUF_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_S_12
#      Description : "Symmetric rise/fall delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_S_12
  CLASS CORE ;
  FOREIGN SEN_BUF_S_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.25 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3933 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.355 1.42 0.485 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.875 1.42 1.005 1.75 ;
      RECT  1.395 1.42 1.525 1.75 ;
      RECT  1.92 1.21 2.04 1.75 ;
      RECT  2.43 1.41 2.565 1.75 ;
      RECT  2.955 1.41 3.085 1.75 ;
      RECT  3.475 1.41 3.605 1.75 ;
      RECT  3.995 1.41 4.125 1.75 ;
      RECT  4.55 1.21 4.67 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  2.155 0.05 2.325 0.32 ;
      RECT  2.675 0.05 2.845 0.32 ;
      RECT  3.195 0.05 3.365 0.32 ;
      RECT  3.715 0.05 3.885 0.32 ;
      RECT  4.235 0.05 4.405 0.32 ;
      RECT  0.615 0.05 0.745 0.365 ;
      RECT  1.135 0.05 1.265 0.37 ;
      RECT  1.66 0.05 1.78 0.555 ;
      RECT  0.08 0.05 0.2 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.895 0.43 4.665 0.55 ;
      RECT  1.895 0.55 4.05 0.56 ;
      RECT  3.75 0.56 4.05 1.11 ;
      RECT  2.15 1.11 4.45 1.29 ;
    END
    ANTENNADIFFAREA 1.127 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.4 0.34 1.52 0.47 ;
      RECT  0.335 0.47 1.52 0.59 ;
      RECT  1.37 0.59 1.52 0.65 ;
      RECT  1.37 0.65 3.64 0.8 ;
      RECT  1.37 0.8 1.52 1.21 ;
      RECT  0.075 1.21 1.82 1.33 ;
  END
END SEN_BUF_S_12
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_S_16
#      Description : "Symmetric rise/fall time buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_S_16
  CLASS CORE ;
  FOREIGN SEN_BUF_S_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.85 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5244 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.345 1.44 0.475 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.865 1.44 0.995 1.75 ;
      RECT  1.385 1.44 1.515 1.75 ;
      RECT  1.905 1.44 2.035 1.75 ;
      RECT  2.46 1.21 2.58 1.75 ;
      RECT  3.005 1.41 3.135 1.75 ;
      RECT  3.525 1.41 3.655 1.75 ;
      RECT  4.045 1.41 4.175 1.75 ;
      RECT  4.565 1.41 4.695 1.75 ;
      RECT  5.085 1.41 5.215 1.75 ;
      RECT  5.625 1.41 5.755 1.75 ;
      RECT  6.19 1.21 6.31 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  2.985 0.05 3.155 0.315 ;
      RECT  3.505 0.05 3.675 0.315 ;
      RECT  4.025 0.05 4.195 0.315 ;
      RECT  4.545 0.05 4.715 0.315 ;
      RECT  5.065 0.05 5.235 0.315 ;
      RECT  5.605 0.05 5.775 0.315 ;
      RECT  0.335 0.05 0.465 0.36 ;
      RECT  0.865 0.05 0.995 0.36 ;
      RECT  1.385 0.05 1.515 0.36 ;
      RECT  1.905 0.05 2.035 0.36 ;
      RECT  2.47 0.05 2.59 0.59 ;
      RECT  6.185 0.05 6.305 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.725 0.425 6.065 0.56 ;
      RECT  2.725 0.56 5.46 0.595 ;
      RECT  5.14 0.595 5.46 1.07 ;
      RECT  2.725 1.07 5.46 1.11 ;
      RECT  2.725 1.11 6.05 1.29 ;
    END
    ANTENNADIFFAREA 1.466 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.34 0.195 0.45 ;
      RECT  0.075 0.45 2.315 0.585 ;
      RECT  2.145 0.585 2.315 0.685 ;
      RECT  2.145 0.685 5.03 0.8 ;
      RECT  2.145 0.8 3.935 0.875 ;
      RECT  2.145 0.875 2.335 1.21 ;
      RECT  0.075 1.21 2.335 1.35 ;
      RECT  0.075 1.35 0.195 1.43 ;
  END
END SEN_BUF_S_16
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_S_2
#      Description : "Symmetric rise/fall delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_S_2
  CLASS CORE ;
  FOREIGN SEN_BUF_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0654 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.63 1.41 0.76 1.75 ;
      RECT  1.21 1.21 1.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.63 0.05 0.76 0.39 ;
      RECT  1.205 0.05 1.335 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.29 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.325 0.37 0.445 0.5 ;
      RECT  0.325 0.5 0.645 0.59 ;
      RECT  0.555 0.59 0.645 0.715 ;
      RECT  0.555 0.715 0.86 0.825 ;
      RECT  0.555 0.825 0.645 1.21 ;
      RECT  0.325 1.21 0.645 1.3 ;
      RECT  0.325 1.3 0.445 1.49 ;
  END
END SEN_BUF_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_S_3
#      Description : "Symmetric rise/fall time buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_S_3
  CLASS CORE ;
  FOREIGN SEN_BUF_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.5 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0978 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.1 1.21 0.22 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.63 1.41 0.76 1.75 ;
      RECT  1.15 1.41 1.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.09 0.05 0.21 0.385 ;
      RECT  0.74 0.05 0.86 0.385 ;
      RECT  1.38 0.05 1.5 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.9 0.51 1.25 0.69 ;
      RECT  1.145 0.69 1.25 1.11 ;
      RECT  0.75 1.11 1.535 1.29 ;
    END
    ANTENNADIFFAREA 0.32 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.32 0.29 0.645 0.39 ;
      RECT  0.555 0.39 0.645 0.78 ;
      RECT  0.555 0.78 1.05 0.89 ;
      RECT  0.555 0.89 0.645 1.21 ;
      RECT  0.32 1.21 0.645 1.31 ;
  END
END SEN_BUF_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_S_4
#      Description : "Symmetric rise/fall delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_S_4
  CLASS CORE ;
  FOREIGN SEN_BUF_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 0.71 ;
      RECT  0.15 0.71 0.665 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1311 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.43 0.5 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  0.94 1.23 1.06 1.75 ;
      RECT  1.475 1.43 1.605 1.75 ;
      RECT  2.015 1.225 2.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  1.475 0.05 1.595 0.345 ;
      RECT  0.94 0.05 1.06 0.56 ;
      RECT  0.39 0.05 0.51 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.185 0.45 1.85 0.56 ;
      RECT  1.745 0.56 1.85 1.105 ;
      RECT  1.15 1.105 1.85 1.295 ;
    END
    ANTENNADIFFAREA 0.391 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.62 0.44 0.85 0.56 ;
      RECT  0.755 0.56 0.85 0.755 ;
      RECT  0.755 0.755 1.635 0.865 ;
      RECT  0.755 0.865 0.85 1.225 ;
      RECT  0.07 1.225 0.85 1.34 ;
  END
END SEN_BUF_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_S_6
#      Description : "Symmetric rise/fall time buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_S_6
  CLASS CORE ;
  FOREIGN SEN_BUF_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.295 0.25 0.635 ;
      RECT  0.15 0.635 0.655 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.39 1.37 0.52 1.75 ;
      RECT  0.0 1.75 2.8 1.85 ;
      RECT  0.955 1.21 1.075 1.75 ;
      RECT  1.485 1.41 1.615 1.75 ;
      RECT  2.025 1.41 2.155 1.75 ;
      RECT  2.57 1.21 2.69 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      RECT  0.925 0.05 1.095 0.31 ;
      RECT  0.365 0.05 0.495 0.39 ;
      RECT  2.025 0.05 2.155 0.39 ;
      RECT  1.49 0.05 1.61 0.59 ;
      RECT  2.57 0.05 2.69 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.745 0.48 2.45 0.6 ;
      RECT  2.35 0.6 2.45 1.11 ;
      RECT  1.18 1.11 2.45 1.29 ;
    END
    ANTENNADIFFAREA 0.548 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.695 0.28 0.805 0.4 ;
      RECT  0.695 0.4 1.36 0.5 ;
      RECT  0.745 0.5 0.85 0.78 ;
      RECT  0.745 0.78 2.245 0.89 ;
      RECT  0.745 0.89 0.84 1.145 ;
      RECT  0.07 1.145 0.84 1.255 ;
  END
END SEN_BUF_S_6
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_S_8
#      Description : "Symmetric rise/fall delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_S_8
  CLASS CORE ;
  FOREIGN SEN_BUF_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 0.655 ;
      RECT  0.15 0.655 0.86 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2619 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      RECT  1.115 1.41 1.245 1.75 ;
      RECT  1.635 1.41 1.765 1.75 ;
      RECT  2.155 1.41 2.285 1.75 ;
      RECT  2.675 1.41 2.805 1.75 ;
      RECT  3.21 1.21 3.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.595 0.05 0.725 0.345 ;
      RECT  1.11 0.05 1.245 0.345 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  1.635 0.05 1.765 0.39 ;
      RECT  2.155 0.05 2.285 0.39 ;
      RECT  2.67 0.05 2.805 0.39 ;
      RECT  3.21 0.05 3.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.865 0.48 3.11 0.595 ;
      RECT  2.68 0.595 2.85 1.11 ;
      RECT  1.35 1.11 3.085 1.29 ;
    END
    ANTENNADIFFAREA 0.732 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.24 0.46 0.435 ;
      RECT  0.34 0.435 1.5 0.545 ;
      RECT  0.86 0.24 0.98 0.435 ;
      RECT  1.38 0.24 1.5 0.435 ;
      RECT  1.125 0.545 1.5 0.555 ;
      RECT  1.125 0.555 1.235 0.775 ;
      RECT  1.125 0.775 2.57 0.89 ;
      RECT  1.125 0.89 1.235 1.21 ;
      RECT  0.315 1.21 1.235 1.32 ;
  END
END SEN_BUF_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_10
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_10
  CLASS CORE ;
  FOREIGN SEN_BUF_10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.84 1.44 0.97 1.75 ;
      RECT  1.365 1.21 1.485 1.75 ;
      RECT  1.88 1.41 2.01 1.75 ;
      RECT  2.4 1.41 2.53 1.75 ;
      RECT  2.92 1.41 3.05 1.75 ;
      RECT  3.44 1.41 3.57 1.75 ;
      RECT  3.98 1.21 4.1 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  1.86 0.05 2.03 0.335 ;
      RECT  2.38 0.05 2.55 0.335 ;
      RECT  2.9 0.05 3.07 0.335 ;
      RECT  3.42 0.05 3.59 0.335 ;
      RECT  0.3 0.05 0.47 0.36 ;
      RECT  0.82 0.05 0.99 0.36 ;
      RECT  1.365 0.05 1.485 0.59 ;
      RECT  3.98 0.05 4.1 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.575 0.435 3.875 0.555 ;
      RECT  1.575 0.555 3.45 0.565 ;
      RECT  3.2 0.565 3.45 1.11 ;
      RECT  1.6 1.11 3.85 1.29 ;
    END
    ANTENNADIFFAREA 1.08 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.35 0.185 0.45 ;
      RECT  0.065 0.45 1.25 0.575 ;
      RECT  1.15 0.575 1.25 0.76 ;
      RECT  1.15 0.76 3.1 0.895 ;
      RECT  1.15 0.895 1.25 1.23 ;
      RECT  0.065 1.23 1.25 1.35 ;
      RECT  0.065 1.35 0.185 1.45 ;
  END
END SEN_BUF_10
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_1P5
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_1P5
  CLASS CORE ;
  FOREIGN SEN_BUF_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.64 0.25 1.175 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.445 0.45 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.945 1.41 1.075 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.32 0.05 0.45 0.365 ;
      RECT  0.945 0.05 1.075 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.85 0.49 ;
      RECT  0.75 0.49 0.85 1.31 ;
      RECT  0.55 1.31 0.85 1.49 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.32 0.185 0.455 ;
      RECT  0.065 0.455 0.445 0.545 ;
      RECT  0.355 0.545 0.445 0.795 ;
      RECT  0.355 0.795 0.66 0.905 ;
      RECT  0.355 0.905 0.46 1.265 ;
      RECT  0.065 1.265 0.46 1.355 ;
      RECT  0.065 1.355 0.185 1.485 ;
  END
END SEN_BUF_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_BUF_20
#      Description : "Non-inverting buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_BUF_20
  CLASS CORE ;
  FOREIGN SEN_BUF_20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.7 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.58 1.42 0.71 1.75 ;
      RECT  1.1 1.42 1.23 1.75 ;
      RECT  1.62 1.42 1.75 1.75 ;
      RECT  2.14 1.42 2.27 1.75 ;
      RECT  2.665 1.21 2.785 1.75 ;
      RECT  3.16 1.455 3.33 1.75 ;
      RECT  3.68 1.455 3.85 1.75 ;
      RECT  4.2 1.455 4.37 1.75 ;
      RECT  4.72 1.455 4.89 1.75 ;
      RECT  5.24 1.455 5.41 1.75 ;
      RECT  5.76 1.455 5.93 1.75 ;
      RECT  6.28 1.455 6.45 1.75 ;
      RECT  6.8 1.455 6.97 1.75 ;
      RECT  7.32 1.455 7.49 1.75 ;
      RECT  7.89 1.21 8.01 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  3.16 0.05 3.33 0.305 ;
      RECT  3.68 0.05 3.85 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.72 0.05 4.89 0.305 ;
      RECT  5.24 0.05 5.41 0.305 ;
      RECT  5.76 0.05 5.93 0.305 ;
      RECT  6.28 0.05 6.45 0.305 ;
      RECT  6.8 0.05 6.97 0.305 ;
      RECT  7.32 0.05 7.49 0.305 ;
      RECT  0.56 0.05 0.73 0.345 ;
      RECT  1.08 0.05 1.25 0.345 ;
      RECT  1.6 0.05 1.77 0.345 ;
      RECT  2.12 0.05 2.29 0.345 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  2.665 0.05 2.785 0.59 ;
      RECT  7.89 0.05 8.01 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.875 0.405 7.75 0.525 ;
      RECT  4.49 0.525 7.75 0.57 ;
      RECT  4.49 0.57 6.05 0.625 ;
      RECT  5.61 0.625 6.05 1.08 ;
      RECT  3.95 1.08 6.05 1.11 ;
      RECT  3.95 1.11 7.75 1.21 ;
      RECT  2.88 1.21 7.75 1.33 ;
    END
    ANTENNADIFFAREA 2.16 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.435 2.56 0.565 ;
      RECT  1.9 0.565 2.56 0.605 ;
      RECT  2.34 0.605 2.56 0.71 ;
      RECT  2.34 0.71 4.45 0.745 ;
      RECT  2.34 0.745 5.48 0.93 ;
      RECT  2.34 0.93 2.56 1.16 ;
      RECT  1.87 1.16 2.56 1.21 ;
      RECT  0.28 1.21 2.56 1.33 ;
      RECT  6.4 0.745 7.56 0.895 ;
      LAYER M2 ;
      RECT  3.74 0.75 7.295 0.85 ;
      LAYER V1 ;
      RECT  3.78 0.75 3.88 0.85 ;
      RECT  4.075 0.75 4.175 0.85 ;
      RECT  4.41 0.75 4.51 0.85 ;
      RECT  4.745 0.75 4.845 0.85 ;
      RECT  5.08 0.75 5.18 0.85 ;
      RECT  6.55 0.75 6.65 0.85 ;
      RECT  6.75 0.75 6.85 0.85 ;
      RECT  6.95 0.75 7.05 0.85 ;
      RECT  7.15 0.75 7.25 0.85 ;
  END
END SEN_BUF_20
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLS_1
#      Description : "Clock Gater, positive clock, synchronous enable, post control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLS_1
  CLASS CORE ;
  FOREIGN SEN_CKGTPLS_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0402 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.31 4.315 0.49 ;
      RECT  4.15 0.49 4.25 1.3 ;
    END
    ANTENNADIFFAREA 0.168 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.65 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  1.13 1.45 1.25 1.75 ;
      RECT  1.89 1.63 2.06 1.75 ;
      RECT  2.645 1.615 2.815 1.75 ;
      RECT  3.775 1.2 3.895 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  2.1 0.05 2.27 0.185 ;
      RECT  1.85 0.05 1.97 0.225 ;
      RECT  3.37 0.05 3.54 0.35 ;
      RECT  1.03 0.05 1.15 0.38 ;
      RECT  0.065 0.05 0.185 0.39 ;
      RECT  3.935 0.05 4.055 0.58 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.36 0.14 3.06 0.23 ;
      RECT  2.36 0.23 2.45 0.32 ;
      RECT  2.97 0.23 3.06 0.62 ;
      RECT  1.595 0.2 1.7 0.32 ;
      RECT  1.595 0.32 2.45 0.41 ;
      RECT  1.595 0.41 1.685 1.07 ;
      RECT  2.97 0.62 3.235 0.71 ;
      RECT  3.135 0.71 3.235 0.95 ;
      RECT  1.595 1.07 1.79 1.18 ;
      RECT  0.5 0.24 0.795 0.36 ;
      RECT  0.705 0.36 0.795 0.5 ;
      RECT  0.705 0.5 1.31 0.59 ;
      RECT  1.21 0.59 1.31 0.91 ;
      RECT  0.705 0.59 0.795 1.2 ;
      RECT  0.55 1.2 0.795 1.32 ;
      RECT  1.26 0.24 1.505 0.36 ;
      RECT  1.4 0.36 1.505 1.09 ;
      RECT  0.98 0.695 1.07 1.09 ;
      RECT  0.98 1.09 1.505 1.18 ;
      RECT  3.15 0.21 3.255 0.44 ;
      RECT  3.15 0.44 3.775 0.53 ;
      RECT  3.655 0.21 3.775 0.44 ;
      RECT  1.97 0.5 2.455 0.62 ;
      RECT  2.365 0.62 2.455 1.185 ;
      RECT  1.955 1.185 2.455 1.27 ;
      RECT  0.905 1.27 2.455 1.305 ;
      RECT  0.905 1.305 2.05 1.36 ;
      RECT  0.905 1.36 0.995 1.455 ;
      RECT  0.34 0.57 0.6 0.68 ;
      RECT  0.34 0.68 0.43 1.455 ;
      RECT  0.34 1.455 0.995 1.545 ;
      RECT  2.545 0.34 2.665 0.98 ;
      RECT  2.545 0.98 2.84 1.15 ;
      RECT  2.545 1.15 2.67 1.41 ;
      RECT  2.375 1.41 2.67 1.45 ;
      RECT  1.435 1.45 2.67 1.5 ;
      RECT  1.435 1.5 2.545 1.54 ;
      RECT  1.435 1.54 1.55 1.66 ;
      RECT  3.955 0.7 4.045 0.98 ;
      RECT  3.555 0.98 4.045 1.07 ;
      RECT  3.555 1.07 3.645 1.38 ;
      RECT  2.775 0.34 2.88 0.8 ;
      RECT  2.775 0.8 3.045 0.89 ;
      RECT  2.94 0.89 3.045 1.38 ;
      RECT  2.94 1.38 3.645 1.47 ;
  END
END SEN_CKGTPLS_1
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLS_12
#      Description : "Clock Gater, positive clock, synchronous enable, post control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLS_12
  CLASS CORE ;
  FOREIGN SEN_CKGTPLS_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 0.71 ;
      RECT  1.75 0.71 2.015 0.9 ;
      RECT  1.75 0.9 1.85 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0372 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0552 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.845 0.435 8.12 0.565 ;
      RECT  7.41 0.565 7.66 1.11 ;
      RECT  5.85 1.11 8.07 1.23 ;
      RECT  5.325 1.23 8.07 1.29 ;
      RECT  5.325 1.29 5.95 1.35 ;
    END
    ANTENNADIFFAREA 1.153 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.51 5.455 0.71 ;
      RECT  4.55 0.71 5.455 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1719 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.18 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  1.025 1.47 1.195 1.75 ;
      RECT  1.795 1.61 1.965 1.75 ;
      RECT  2.64 1.21 2.76 1.75 ;
      RECT  3.24 1.44 3.37 1.75 ;
      RECT  4.565 1.45 4.695 1.75 ;
      RECT  5.09 1.21 5.21 1.75 ;
      RECT  5.605 1.44 5.735 1.75 ;
      RECT  6.125 1.41 6.255 1.75 ;
      RECT  6.645 1.41 6.775 1.75 ;
      RECT  7.165 1.41 7.295 1.75 ;
      RECT  7.685 1.41 7.815 1.75 ;
      RECT  8.21 1.21 8.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  1.815 0.05 1.945 0.235 ;
      RECT  6.105 0.05 6.275 0.325 ;
      RECT  6.625 0.05 6.795 0.325 ;
      RECT  7.145 0.05 7.315 0.325 ;
      RECT  7.665 0.05 7.835 0.325 ;
      RECT  3.865 0.05 3.995 0.35 ;
      RECT  4.385 0.05 4.515 0.35 ;
      RECT  4.905 0.05 5.035 0.35 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  2.315 0.05 2.445 0.415 ;
      RECT  0.98 0.05 1.11 0.495 ;
      RECT  5.59 0.05 5.71 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.335 0.14 1.445 0.22 ;
      RECT  1.335 0.22 1.605 0.31 ;
      RECT  1.515 0.31 1.605 0.325 ;
      RECT  1.515 0.325 2.21 0.415 ;
      RECT  2.105 0.415 2.21 0.835 ;
      RECT  2.105 0.835 2.505 0.925 ;
      RECT  2.415 0.755 2.505 0.835 ;
      RECT  2.105 0.925 2.21 1.25 ;
      RECT  0.705 1.25 2.21 1.34 ;
      RECT  0.705 1.34 0.8 1.56 ;
      RECT  5.14 0.215 5.35 0.335 ;
      RECT  5.14 0.335 5.23 0.44 ;
      RECT  3.04 0.235 3.73 0.35 ;
      RECT  3.61 0.35 3.73 0.44 ;
      RECT  3.61 0.44 5.23 0.56 ;
      RECT  0.515 0.39 0.635 0.585 ;
      RECT  0.515 0.585 1.205 0.675 ;
      RECT  1.115 0.675 1.205 0.935 ;
      RECT  0.515 0.675 0.62 1.22 ;
      RECT  2.595 0.405 2.7 0.835 ;
      RECT  2.595 0.835 3.335 0.945 ;
      RECT  2.595 0.945 2.685 1.02 ;
      RECT  2.32 1.02 2.685 1.11 ;
      RECT  2.32 1.11 2.44 1.43 ;
      RECT  1.295 1.43 2.44 1.52 ;
      RECT  1.295 1.52 1.385 1.66 ;
      RECT  5.545 0.765 7.28 0.875 ;
      RECT  5.545 0.875 5.65 1.0 ;
      RECT  4.05 1.0 5.65 1.12 ;
      RECT  4.05 1.12 4.17 1.24 ;
      RECT  2.79 0.44 3.515 0.56 ;
      RECT  3.425 0.56 3.515 1.24 ;
      RECT  2.935 1.24 4.17 1.35 ;
      RECT  3.75 0.71 4.24 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
      RECT  0.885 0.765 0.975 1.07 ;
      RECT  0.885 1.07 1.425 1.16 ;
      RECT  1.32 0.42 1.425 1.07 ;
      RECT  1.55 0.51 1.66 1.16 ;
      RECT  4.31 1.24 4.975 1.36 ;
      RECT  4.31 1.36 4.43 1.44 ;
      RECT  3.765 1.44 4.43 1.56 ;
      LAYER M2 ;
      RECT  1.51 0.95 3.89 1.05 ;
      LAYER V1 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  3.75 0.95 3.85 1.05 ;
  END
END SEN_CKGTPLS_12
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLS_16
#      Description : "Clock Gater, positive clock, synchronous enable, post control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLS_16
  CLASS CORE ;
  FOREIGN SEN_CKGTPLS_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 0.71 ;
      RECT  1.75 0.71 2.015 0.9 ;
      RECT  1.75 0.9 1.85 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0387 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.84 0.415 9.13 0.535 ;
      RECT  6.385 0.535 9.13 0.585 ;
      RECT  7.93 0.585 9.13 0.69 ;
      RECT  7.93 0.69 8.25 1.11 ;
      RECT  6.35 1.11 9.13 1.23 ;
      RECT  5.32 1.23 9.13 1.35 ;
    END
    ANTENNADIFFAREA 1.555 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.51 5.455 0.71 ;
      RECT  4.55 0.71 5.455 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.18 1.75 ;
      RECT  0.0 1.75 9.2 1.85 ;
      RECT  1.025 1.47 1.195 1.75 ;
      RECT  1.795 1.61 1.965 1.75 ;
      RECT  2.67 1.24 2.79 1.75 ;
      RECT  3.26 1.44 3.39 1.75 ;
      RECT  4.585 1.45 4.715 1.75 ;
      RECT  5.11 1.215 5.23 1.75 ;
      RECT  5.625 1.44 5.755 1.75 ;
      RECT  6.145 1.44 6.275 1.75 ;
      RECT  6.665 1.44 6.795 1.75 ;
      RECT  7.185 1.44 7.315 1.75 ;
      RECT  7.705 1.44 7.835 1.75 ;
      RECT  8.225 1.44 8.355 1.75 ;
      RECT  8.745 1.44 8.875 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.2 0.05 ;
      RECT  1.815 0.05 1.945 0.235 ;
      RECT  6.125 0.05 6.295 0.325 ;
      RECT  6.645 0.05 6.815 0.325 ;
      RECT  7.165 0.05 7.335 0.325 ;
      RECT  7.685 0.05 7.855 0.325 ;
      RECT  8.205 0.05 8.375 0.325 ;
      RECT  8.725 0.05 8.895 0.325 ;
      RECT  3.885 0.05 4.015 0.35 ;
      RECT  4.405 0.05 4.535 0.35 ;
      RECT  4.925 0.05 5.055 0.35 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  0.98 0.05 1.11 0.495 ;
      RECT  2.34 0.05 2.46 0.59 ;
      RECT  5.58 0.05 5.7 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.34 0.14 1.44 0.22 ;
      RECT  1.34 0.22 1.605 0.31 ;
      RECT  1.515 0.31 1.605 0.325 ;
      RECT  1.515 0.325 2.21 0.415 ;
      RECT  2.105 0.415 2.21 0.835 ;
      RECT  2.105 0.835 2.51 0.925 ;
      RECT  2.41 0.755 2.51 0.835 ;
      RECT  2.105 0.925 2.21 1.25 ;
      RECT  0.705 1.25 2.21 1.34 ;
      RECT  0.705 1.34 0.795 1.56 ;
      RECT  5.16 0.215 5.36 0.335 ;
      RECT  5.16 0.335 5.25 0.44 ;
      RECT  3.06 0.24 3.75 0.35 ;
      RECT  3.63 0.35 3.75 0.44 ;
      RECT  3.63 0.44 5.25 0.56 ;
      RECT  0.515 0.375 0.635 0.585 ;
      RECT  0.515 0.585 1.205 0.675 ;
      RECT  1.115 0.675 1.205 0.935 ;
      RECT  0.515 0.675 0.62 1.22 ;
      RECT  2.6 0.475 2.72 0.795 ;
      RECT  2.6 0.795 3.355 0.905 ;
      RECT  2.6 0.905 2.705 1.015 ;
      RECT  2.34 1.015 2.705 1.105 ;
      RECT  2.34 1.105 2.46 1.43 ;
      RECT  1.295 1.43 2.46 1.52 ;
      RECT  1.295 1.52 1.385 1.66 ;
      RECT  5.545 0.72 7.78 0.83 ;
      RECT  5.545 0.83 5.65 1.0 ;
      RECT  4.07 1.0 5.65 1.12 ;
      RECT  4.07 1.12 4.19 1.24 ;
      RECT  2.81 0.44 3.535 0.56 ;
      RECT  3.445 0.56 3.535 1.24 ;
      RECT  2.955 1.24 4.19 1.35 ;
      RECT  3.75 0.71 4.24 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
      RECT  0.885 0.765 0.975 1.07 ;
      RECT  0.885 1.07 1.425 1.16 ;
      RECT  1.32 0.44 1.425 1.07 ;
      RECT  1.55 0.51 1.66 1.16 ;
      RECT  4.33 1.24 5.02 1.36 ;
      RECT  4.33 1.36 4.45 1.44 ;
      RECT  3.76 1.44 4.45 1.56 ;
      LAYER M2 ;
      RECT  1.51 0.95 3.89 1.05 ;
      LAYER V1 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  3.75 0.95 3.85 1.05 ;
  END
END SEN_CKGTPLS_16
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLS_2
#      Description : "Clock Gater, positive clock, synchronous enable, post control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLS_2
  CLASS CORE ;
  FOREIGN SEN_CKGTPLS_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0354 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0432 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.31 4.25 1.3 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.65 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0447 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  1.13 1.45 1.25 1.75 ;
      RECT  1.89 1.63 2.06 1.75 ;
      RECT  2.645 1.615 2.815 1.75 ;
      RECT  3.775 1.2 3.895 1.75 ;
      RECT  4.405 1.21 4.525 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.1 0.05 2.27 0.185 ;
      RECT  1.85 0.05 1.97 0.225 ;
      RECT  3.37 0.05 3.54 0.35 ;
      RECT  1.03 0.05 1.15 0.38 ;
      RECT  0.065 0.05 0.185 0.39 ;
      RECT  3.885 0.05 4.005 0.39 ;
      RECT  4.405 0.05 4.525 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.36 0.14 3.06 0.23 ;
      RECT  2.36 0.23 2.45 0.32 ;
      RECT  2.97 0.23 3.06 0.62 ;
      RECT  1.595 0.2 1.7 0.32 ;
      RECT  1.595 0.32 2.45 0.41 ;
      RECT  1.595 0.41 1.685 1.07 ;
      RECT  2.97 0.62 3.235 0.71 ;
      RECT  3.135 0.71 3.235 0.96 ;
      RECT  1.595 1.07 1.79 1.18 ;
      RECT  0.5 0.24 0.795 0.36 ;
      RECT  0.705 0.36 0.795 0.5 ;
      RECT  0.705 0.5 1.31 0.59 ;
      RECT  1.21 0.59 1.31 0.915 ;
      RECT  0.705 0.59 0.795 1.2 ;
      RECT  0.55 1.2 0.795 1.32 ;
      RECT  1.26 0.24 1.505 0.36 ;
      RECT  1.4 0.36 1.505 1.09 ;
      RECT  0.98 0.695 1.07 1.09 ;
      RECT  0.98 1.09 1.505 1.18 ;
      RECT  3.15 0.225 3.255 0.44 ;
      RECT  3.15 0.44 3.775 0.53 ;
      RECT  3.655 0.225 3.775 0.44 ;
      RECT  1.97 0.5 2.455 0.62 ;
      RECT  2.365 0.62 2.455 1.185 ;
      RECT  1.955 1.185 2.455 1.27 ;
      RECT  0.905 1.27 2.455 1.305 ;
      RECT  0.905 1.305 2.05 1.36 ;
      RECT  0.905 1.36 0.995 1.455 ;
      RECT  0.34 0.57 0.6 0.68 ;
      RECT  0.34 0.68 0.43 1.455 ;
      RECT  0.34 1.455 0.995 1.545 ;
      RECT  2.545 0.34 2.665 0.98 ;
      RECT  2.545 0.98 2.84 1.15 ;
      RECT  2.545 1.15 2.67 1.41 ;
      RECT  2.375 1.41 2.67 1.45 ;
      RECT  1.46 1.45 2.67 1.5 ;
      RECT  1.46 1.5 2.545 1.54 ;
      RECT  1.46 1.54 1.57 1.66 ;
      RECT  3.955 0.685 4.045 0.98 ;
      RECT  3.555 0.98 4.045 1.07 ;
      RECT  3.555 1.07 3.645 1.38 ;
      RECT  2.775 0.34 2.88 0.8 ;
      RECT  2.775 0.8 3.045 0.89 ;
      RECT  2.94 0.89 3.045 1.38 ;
      RECT  2.94 1.38 3.645 1.47 ;
  END
END SEN_CKGTPLS_2
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLS_3
#      Description : "Clock Gater, positive clock, synchronous enable, post control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLS_3
  CLASS CORE ;
  FOREIGN SEN_CKGTPLS_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0459 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.31 4.28 0.51 ;
      RECT  4.15 0.51 4.45 0.6 ;
      RECT  4.35 0.6 4.45 1.11 ;
      RECT  3.92 1.11 4.535 1.29 ;
    END
    ANTENNADIFFAREA 0.293 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.65 0.89 ;
      RECT  3.55 0.89 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  1.085 1.45 1.205 1.75 ;
      RECT  1.845 1.62 2.015 1.75 ;
      RECT  2.725 1.45 2.845 1.75 ;
      RECT  3.61 1.45 3.73 1.75 ;
      RECT  4.165 1.415 4.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.2 0.05 2.37 0.175 ;
      RECT  1.78 0.05 1.95 0.185 ;
      RECT  3.905 0.05 4.025 0.37 ;
      RECT  1.02 0.05 1.15 0.385 ;
      RECT  4.425 0.05 4.545 0.385 ;
      RECT  0.065 0.05 0.185 0.39 ;
      RECT  3.41 0.05 3.58 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.495 0.145 3.08 0.235 ;
      RECT  2.495 0.235 2.585 0.295 ;
      RECT  2.99 0.235 3.08 0.71 ;
      RECT  1.545 0.295 2.585 0.385 ;
      RECT  1.545 0.385 1.65 0.915 ;
      RECT  2.99 0.71 3.245 0.8 ;
      RECT  3.135 0.8 3.245 1.0 ;
      RECT  1.55 0.915 1.65 1.065 ;
      RECT  1.55 1.065 1.76 1.17 ;
      RECT  1.26 0.24 1.455 0.36 ;
      RECT  1.355 0.36 1.455 0.99 ;
      RECT  1.355 0.99 1.46 1.07 ;
      RECT  0.925 0.815 1.035 1.07 ;
      RECT  0.925 1.07 1.46 1.16 ;
      RECT  0.47 0.265 0.78 0.385 ;
      RECT  0.69 0.385 0.78 0.51 ;
      RECT  0.69 0.51 1.26 0.6 ;
      RECT  1.14 0.6 1.26 0.75 ;
      RECT  0.69 0.6 0.78 1.19 ;
      RECT  0.54 1.19 0.78 1.36 ;
      RECT  3.17 0.38 3.28 0.51 ;
      RECT  3.17 0.51 3.815 0.6 ;
      RECT  3.695 0.415 3.815 0.51 ;
      RECT  1.91 0.515 2.435 0.62 ;
      RECT  2.34 0.62 2.435 1.26 ;
      RECT  0.87 1.26 2.435 1.35 ;
      RECT  0.87 1.35 0.96 1.46 ;
      RECT  0.36 0.59 0.595 0.7 ;
      RECT  0.36 0.7 0.45 1.46 ;
      RECT  0.36 1.46 0.96 1.55 ;
      RECT  2.525 0.52 2.63 0.8 ;
      RECT  2.525 0.8 2.72 0.97 ;
      RECT  2.525 0.97 2.635 1.44 ;
      RECT  1.375 1.44 2.635 1.53 ;
      RECT  3.74 0.78 4.26 0.895 ;
      RECT  3.74 0.895 3.83 1.24 ;
      RECT  2.69 0.325 2.9 0.43 ;
      RECT  2.81 0.43 2.9 1.24 ;
      RECT  2.81 1.24 3.83 1.36 ;
  END
END SEN_CKGTPLS_3
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLS_4
#      Description : "Clock Gater, positive clock, synchronous enable, post control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLS_4
  CLASS CORE ;
  FOREIGN SEN_CKGTPLS_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0387 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0477 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.6 0.36 4.72 0.51 ;
      RECT  3.95 0.51 4.72 0.69 ;
      RECT  4.35 0.69 4.45 1.11 ;
      RECT  3.82 1.11 4.45 1.295 ;
    END
    ANTENNADIFFAREA 0.394 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.45 0.755 ;
      RECT  3.35 0.755 3.515 0.925 ;
      RECT  3.35 0.925 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  1.13 1.44 1.25 1.75 ;
      RECT  1.895 1.63 2.065 1.75 ;
      RECT  2.735 1.415 2.85 1.75 ;
      RECT  3.55 1.415 3.67 1.75 ;
      RECT  4.08 1.415 4.2 1.75 ;
      RECT  4.6 1.215 4.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  2.255 0.05 2.425 0.2 ;
      RECT  3.3 0.05 3.47 0.2 ;
      RECT  1.905 0.05 2.035 0.28 ;
      RECT  4.34 0.05 4.48 0.37 ;
      RECT  1.085 0.05 1.205 0.385 ;
      RECT  0.065 0.05 0.185 0.39 ;
      RECT  3.82 0.05 3.94 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.53 0.24 0.805 0.36 ;
      RECT  0.715 0.36 0.805 0.51 ;
      RECT  0.715 0.51 1.31 0.6 ;
      RECT  1.21 0.6 1.31 0.775 ;
      RECT  0.715 0.6 0.805 1.18 ;
      RECT  0.56 1.18 0.805 1.3 ;
      RECT  1.37 0.215 1.49 0.385 ;
      RECT  1.4 0.385 1.49 0.99 ;
      RECT  1.4 0.99 1.505 1.07 ;
      RECT  0.96 0.815 1.07 1.07 ;
      RECT  0.96 1.07 1.505 1.16 ;
      RECT  3.02 0.29 3.715 0.41 ;
      RECT  3.595 0.41 3.715 0.67 ;
      RECT  1.99 0.5 2.45 0.62 ;
      RECT  2.355 0.62 2.45 1.26 ;
      RECT  0.91 1.26 2.45 1.35 ;
      RECT  0.91 1.35 1.0 1.46 ;
      RECT  0.36 0.605 0.6 0.715 ;
      RECT  0.36 0.715 0.45 1.46 ;
      RECT  0.36 1.46 1.0 1.55 ;
      RECT  2.555 0.5 2.685 0.77 ;
      RECT  2.555 0.77 2.75 0.94 ;
      RECT  2.555 0.94 2.645 1.44 ;
      RECT  1.545 1.44 2.645 1.53 ;
      RECT  2.315 1.53 2.485 1.655 ;
      RECT  1.545 1.53 1.655 1.66 ;
      RECT  3.605 0.785 4.26 0.895 ;
      RECT  3.605 0.895 3.695 1.205 ;
      RECT  2.795 0.42 2.93 0.615 ;
      RECT  2.84 0.615 2.93 1.205 ;
      RECT  2.84 1.205 3.695 1.325 ;
      RECT  1.6 0.24 1.72 1.065 ;
      RECT  1.6 1.065 1.81 1.17 ;
      RECT  3.14 0.51 3.25 1.09 ;
      LAYER M2 ;
      RECT  1.58 0.55 3.28 0.65 ;
      LAYER V1 ;
      RECT  1.62 0.55 1.72 0.65 ;
      RECT  3.14 0.55 3.24 0.65 ;
  END
END SEN_CKGTPLS_4
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLS_6
#      Description : "Clock Gater, positive clock, synchronous enable, post control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLS_6
  CLASS CORE ;
  FOREIGN SEN_CKGTPLS_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0399 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.91 0.45 1.09 ;
      RECT  0.35 1.09 0.45 1.5 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0501 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.19 0.48 5.87 0.6 ;
      RECT  5.75 0.6 5.87 1.11 ;
      RECT  5.15 1.11 5.87 1.19 ;
      RECT  4.7 1.19 5.87 1.29 ;
    END
    ANTENNADIFFAREA 0.552 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 4.85 0.7 ;
      RECT  4.15 0.7 4.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0768 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  1.245 1.21 1.375 1.75 ;
      RECT  2.025 1.38 2.145 1.75 ;
      RECT  2.88 1.36 3.01 1.75 ;
      RECT  3.405 1.44 3.52 1.75 ;
      RECT  4.465 1.215 4.585 1.75 ;
      RECT  4.98 1.4 5.11 1.75 ;
      RECT  5.5 1.4 5.63 1.75 ;
      RECT  6.02 1.41 6.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  3.65 0.05 3.82 0.21 ;
      RECT  1.175 0.05 1.28 0.37 ;
      RECT  4.24 0.05 4.37 0.385 ;
      RECT  5.5 0.05 5.63 0.39 ;
      RECT  6.02 0.05 6.145 0.39 ;
      RECT  2.625 0.05 2.745 0.42 ;
      RECT  2.14 0.05 2.255 0.435 ;
      RECT  0.065 0.05 0.185 0.545 ;
      RECT  4.96 0.05 5.08 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.37 0.15 2.05 0.24 ;
      RECT  1.37 0.24 1.46 0.46 ;
      RECT  1.96 0.24 2.05 0.53 ;
      RECT  0.34 0.14 0.905 0.23 ;
      RECT  0.815 0.23 0.905 0.46 ;
      RECT  0.815 0.46 1.46 0.55 ;
      RECT  1.96 0.53 2.485 0.62 ;
      RECT  2.365 0.29 2.485 0.53 ;
      RECT  2.375 0.62 2.485 1.44 ;
      RECT  2.27 1.44 2.485 1.56 ;
      RECT  3.365 0.3 4.065 0.42 ;
      RECT  3.945 0.42 4.065 0.5 ;
      RECT  3.945 0.5 4.66 0.59 ;
      RECT  4.545 0.26 4.66 0.5 ;
      RECT  0.555 0.5 0.675 0.66 ;
      RECT  0.555 0.66 1.46 0.75 ;
      RECT  1.35 0.75 1.46 0.86 ;
      RECT  0.555 0.75 0.675 1.35 ;
      RECT  2.885 0.27 3.005 0.88 ;
      RECT  2.885 0.88 3.065 0.92 ;
      RECT  2.625 0.92 3.065 1.05 ;
      RECT  2.625 1.05 2.745 1.49 ;
      RECT  4.96 0.785 5.66 0.895 ;
      RECT  4.96 0.895 5.05 1.01 ;
      RECT  4.21 1.01 5.05 1.1 ;
      RECT  4.21 1.1 4.3 1.23 ;
      RECT  3.155 0.19 3.265 1.23 ;
      RECT  3.155 1.23 4.3 1.35 ;
      RECT  3.155 1.35 3.265 1.53 ;
      RECT  1.55 0.33 1.655 0.95 ;
      RECT  1.095 0.95 1.655 1.04 ;
      RECT  1.535 1.04 1.655 1.42 ;
      RECT  3.36 0.51 3.46 0.95 ;
      RECT  3.36 0.95 3.83 1.05 ;
      RECT  1.765 0.33 1.87 1.42 ;
      RECT  3.61 1.465 4.355 1.585 ;
      RECT  0.895 0.865 1.005 1.66 ;
      LAYER M2 ;
      RECT  1.73 0.55 3.5 0.65 ;
      RECT  0.865 1.35 2.78 1.45 ;
      LAYER V1 ;
      RECT  1.77 0.55 1.87 0.65 ;
      RECT  3.36 0.55 3.46 0.65 ;
      RECT  0.905 1.35 1.005 1.45 ;
      RECT  2.64 1.35 2.74 1.45 ;
  END
END SEN_CKGTPLS_6
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLS_8
#      Description : "Clock Gater, positive clock, synchronous enable, post control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN):Q=CK&(iq|SE)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLS_8
  CLASS CORE ;
  FOREIGN SEN_CKGTPLS_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  2.15 0.71 2.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0537 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.97 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.31 6.85 0.45 ;
      RECT  5.0 0.45 6.85 0.58 ;
      RECT  6.68 0.58 6.85 1.11 ;
      RECT  5.15 1.11 6.88 1.29 ;
    END
    ANTENNADIFFAREA 0.765 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.45 0.71 ;
      RECT  4.35 0.71 4.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1032 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.18 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  1.485 1.255 1.605 1.75 ;
      RECT  2.19 1.41 2.32 1.75 ;
      RECT  2.965 1.215 3.085 1.75 ;
      RECT  3.48 1.44 3.61 1.75 ;
      RECT  4.415 1.41 4.545 1.75 ;
      RECT  4.94 1.21 5.06 1.75 ;
      RECT  5.455 1.415 5.585 1.75 ;
      RECT  5.975 1.415 6.105 1.75 ;
      RECT  6.495 1.415 6.625 1.75 ;
      RECT  7.015 1.41 7.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  1.26 0.05 1.43 0.185 ;
      RECT  2.12 0.05 2.29 0.185 ;
      RECT  3.82 0.05 3.99 0.185 ;
      RECT  4.425 0.05 4.595 0.185 ;
      RECT  5.315 0.05 5.445 0.36 ;
      RECT  5.885 0.05 6.015 0.36 ;
      RECT  6.455 0.05 6.585 0.36 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  2.575 0.05 2.745 0.39 ;
      RECT  7.0 0.05 7.12 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.055 0.18 3.175 0.275 ;
      RECT  3.055 0.275 4.92 0.39 ;
      RECT  0.43 0.275 2.45 0.385 ;
      RECT  2.34 0.385 2.45 0.485 ;
      RECT  0.43 0.385 0.53 0.97 ;
      RECT  2.34 0.485 2.63 0.605 ;
      RECT  2.54 0.605 2.63 0.715 ;
      RECT  2.54 0.715 2.875 0.815 ;
      RECT  2.54 0.815 2.63 1.17 ;
      RECT  2.4 1.17 2.63 1.29 ;
      RECT  0.62 0.495 1.45 0.585 ;
      RECT  1.36 0.585 1.45 0.865 ;
      RECT  0.62 0.585 0.735 1.17 ;
      RECT  1.36 0.865 1.655 0.975 ;
      RECT  1.84 0.475 2.05 0.595 ;
      RECT  1.945 0.595 2.05 1.63 ;
      RECT  2.82 0.485 3.095 0.595 ;
      RECT  2.985 0.595 3.095 0.745 ;
      RECT  2.985 0.745 3.455 0.855 ;
      RECT  2.985 0.855 3.095 0.95 ;
      RECT  2.72 0.95 3.095 1.05 ;
      RECT  2.72 1.05 2.825 1.34 ;
      RECT  1.54 0.485 1.735 0.605 ;
      RECT  1.625 0.605 1.735 0.685 ;
      RECT  1.625 0.685 1.855 0.775 ;
      RECT  1.745 0.775 1.855 1.07 ;
      RECT  1.175 0.88 1.27 1.07 ;
      RECT  1.175 1.07 1.855 1.16 ;
      RECT  1.745 1.16 1.855 1.39 ;
      RECT  4.78 0.715 6.57 0.825 ;
      RECT  4.78 0.825 4.87 0.98 ;
      RECT  3.26 0.48 4.12 0.59 ;
      RECT  4.03 0.59 4.12 0.98 ;
      RECT  4.03 0.98 4.87 1.07 ;
      RECT  4.03 1.07 4.12 1.23 ;
      RECT  3.185 1.23 4.12 1.35 ;
      RECT  0.83 0.71 1.085 0.89 ;
      RECT  0.975 0.89 1.085 1.17 ;
      RECT  3.825 0.685 3.92 0.895 ;
      RECT  3.575 0.895 3.92 1.095 ;
      RECT  0.33 1.07 0.435 1.26 ;
      RECT  0.33 1.26 1.16 1.38 ;
      RECT  4.21 1.16 4.84 1.28 ;
      RECT  4.21 1.28 4.3 1.55 ;
      RECT  3.715 1.44 3.835 1.55 ;
      RECT  3.715 1.55 4.3 1.64 ;
      RECT  0.45 1.47 1.375 1.585 ;
      LAYER M2 ;
      RECT  0.945 0.95 2.9 1.05 ;
      RECT  3.07 0.95 3.915 1.05 ;
      RECT  3.07 1.05 3.17 1.15 ;
      RECT  1.91 1.15 3.17 1.25 ;
      LAYER V1 ;
      RECT  0.985 0.95 1.085 1.05 ;
      RECT  2.76 0.95 2.86 1.05 ;
      RECT  3.575 0.95 3.675 1.05 ;
      RECT  3.775 0.95 3.875 1.05 ;
      RECT  1.95 1.15 2.05 1.25 ;
  END
END SEN_CKGTPLS_8
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLT_1
#      Description : "Clock Gater, positive clock, synchronous enable, pre control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLT_1
  CLASS CORE ;
  FOREIGN SEN_CKGTPLT_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  2.15 0.71 2.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.27 4.135 0.44 ;
      RECT  3.95 0.44 4.05 1.29 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.0 ;
      RECT  0.15 1.0 0.45 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0402 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  1.365 1.245 1.495 1.75 ;
      RECT  2.15 1.52 2.32 1.75 ;
      RECT  2.965 1.41 3.095 1.75 ;
      RECT  3.525 1.55 3.675 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  2.15 0.05 2.32 0.175 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  2.965 0.05 3.095 0.39 ;
      RECT  3.735 0.05 3.86 0.39 ;
      RECT  1.345 0.05 1.515 0.495 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.74 0.14 1.85 0.265 ;
      RECT  1.74 0.265 2.58 0.355 ;
      RECT  2.46 0.355 2.58 0.53 ;
      RECT  2.46 0.53 2.63 0.62 ;
      RECT  2.54 0.62 2.63 0.845 ;
      RECT  2.54 0.845 2.96 0.955 ;
      RECT  2.54 0.955 2.63 1.195 ;
      RECT  2.46 1.195 2.63 1.34 ;
      RECT  1.775 1.34 2.63 1.43 ;
      RECT  1.775 1.43 1.885 1.63 ;
      RECT  0.065 0.26 0.185 0.49 ;
      RECT  0.065 0.49 0.705 0.58 ;
      RECT  0.585 0.21 0.705 0.49 ;
      RECT  3.49 0.22 3.61 0.5 ;
      RECT  3.49 0.5 3.855 0.59 ;
      RECT  3.745 0.59 3.855 1.34 ;
      RECT  3.205 1.34 3.855 1.46 ;
      RECT  1.86 0.445 2.035 0.565 ;
      RECT  1.86 0.565 1.965 1.13 ;
      RECT  1.86 1.13 2.37 1.25 ;
      RECT  0.845 0.41 0.975 0.585 ;
      RECT  0.845 0.585 1.55 0.675 ;
      RECT  1.44 0.675 1.55 0.92 ;
      RECT  0.845 0.675 0.955 1.5 ;
      RECT  2.72 0.21 2.83 0.6 ;
      RECT  2.72 0.6 3.16 0.69 ;
      RECT  3.06 0.69 3.16 1.08 ;
      RECT  2.72 1.08 3.16 1.17 ;
      RECT  2.72 1.17 2.83 1.545 ;
      RECT  2.48 1.545 2.83 1.655 ;
      RECT  1.21 0.765 1.32 1.055 ;
      RECT  1.21 1.055 1.76 1.145 ;
      RECT  1.64 0.46 1.76 1.055 ;
      RECT  3.34 0.715 3.45 1.15 ;
      RECT  3.25 1.15 3.45 1.25 ;
      LAYER M2 ;
      RECT  2.19 1.15 3.43 1.25 ;
      LAYER V1 ;
      RECT  2.23 1.15 2.33 1.25 ;
      RECT  3.29 1.15 3.39 1.25 ;
  END
END SEN_CKGTPLT_1
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLT_12
#      Description : "Clock Gater, positive clock, synchronous enable, pre control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLT_12
  CLASS CORE ;
  FOREIGN SEN_CKGTPLT_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.73 ;
      RECT  2.15 0.73 2.345 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0372 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0597 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.23 0.46 7.535 0.585 ;
      RECT  5.23 0.585 7.05 0.59 ;
      RECT  6.8 0.59 7.05 1.11 ;
      RECT  4.74 1.11 7.65 1.29 ;
    END
    ANTENNADIFFAREA 1.158 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0597 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.195 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  1.34 1.495 1.51 1.75 ;
      RECT  2.125 1.615 2.295 1.75 ;
      RECT  2.93 1.21 3.05 1.75 ;
      RECT  3.445 1.45 3.575 1.75 ;
      RECT  3.98 1.45 4.11 1.75 ;
      RECT  4.5 1.45 4.63 1.75 ;
      RECT  5.02 1.41 5.15 1.75 ;
      RECT  5.54 1.41 5.67 1.75 ;
      RECT  6.06 1.41 6.19 1.75 ;
      RECT  6.58 1.41 6.71 1.75 ;
      RECT  7.1 1.41 7.23 1.75 ;
      RECT  7.62 1.41 7.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  2.11 0.05 2.28 0.22 ;
      RECT  5.52 0.05 5.69 0.325 ;
      RECT  6.04 0.05 6.21 0.325 ;
      RECT  6.56 0.05 6.73 0.325 ;
      RECT  7.08 0.05 7.25 0.325 ;
      RECT  0.325 0.05 0.455 0.35 ;
      RECT  3.445 0.05 3.575 0.35 ;
      RECT  2.925 0.05 3.055 0.36 ;
      RECT  1.315 0.05 1.445 0.46 ;
      RECT  5.0 0.05 5.12 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.705 0.14 1.92 0.31 ;
      RECT  1.83 0.31 2.525 0.4 ;
      RECT  2.435 0.4 2.525 0.835 ;
      RECT  2.435 0.835 2.88 0.925 ;
      RECT  2.79 0.755 2.88 0.835 ;
      RECT  2.435 0.925 2.525 1.255 ;
      RECT  1.36 1.255 2.525 1.3 ;
      RECT  0.98 1.3 2.525 1.345 ;
      RECT  0.98 1.345 1.45 1.39 ;
      RECT  0.98 1.39 1.07 1.605 ;
      RECT  3.71 0.24 4.415 0.36 ;
      RECT  3.71 0.36 3.83 0.44 ;
      RECT  3.15 0.44 3.83 0.56 ;
      RECT  0.07 0.34 0.19 0.44 ;
      RECT  0.07 0.44 0.76 0.56 ;
      RECT  0.85 0.36 0.97 0.55 ;
      RECT  0.85 0.55 1.54 0.675 ;
      RECT  1.45 0.675 1.54 0.825 ;
      RECT  0.85 0.675 0.96 1.09 ;
      RECT  0.755 1.09 0.96 1.21 ;
      RECT  3.93 0.45 4.625 0.57 ;
      RECT  4.505 0.57 4.625 0.745 ;
      RECT  4.505 0.745 6.68 0.88 ;
      RECT  4.505 0.88 4.625 1.24 ;
      RECT  3.14 1.24 4.625 1.36 ;
      RECT  2.62 0.455 3.06 0.575 ;
      RECT  2.97 0.575 3.06 0.74 ;
      RECT  2.97 0.74 3.625 0.85 ;
      RECT  2.97 0.85 3.06 1.015 ;
      RECT  2.67 1.015 3.06 1.105 ;
      RECT  2.67 1.105 2.79 1.435 ;
      RECT  1.61 1.435 2.79 1.525 ;
      RECT  1.61 1.525 1.7 1.66 ;
      RECT  1.215 0.765 1.31 0.915 ;
      RECT  1.215 0.915 1.74 1.005 ;
      RECT  1.63 0.435 1.74 0.915 ;
      RECT  1.635 1.005 1.74 1.16 ;
      RECT  3.83 0.83 4.365 0.935 ;
      RECT  3.83 0.935 3.94 0.95 ;
      RECT  3.29 0.95 3.94 1.05 ;
      RECT  1.865 0.52 1.985 1.16 ;
      LAYER M2 ;
      RECT  1.83 0.95 3.47 1.05 ;
      LAYER V1 ;
      RECT  1.87 0.95 1.97 1.05 ;
      RECT  3.33 0.95 3.43 1.05 ;
  END
END SEN_CKGTPLT_12
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLT_16
#      Description : "Clock Gater, positive clock, synchronous enable, pre control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLT_16
  CLASS CORE ;
  FOREIGN SEN_CKGTPLT_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.75 ;
      RECT  2.15 0.75 2.345 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0387 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.235 0.415 8.525 0.535 ;
      RECT  5.78 0.535 8.525 0.585 ;
      RECT  7.33 0.585 8.525 0.69 ;
      RECT  7.33 0.69 7.65 1.11 ;
      RECT  5.745 1.11 8.525 1.23 ;
      RECT  4.715 1.23 8.525 1.35 ;
    END
    ANTENNADIFFAREA 1.555 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.195 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  1.34 1.495 1.51 1.75 ;
      RECT  2.125 1.615 2.295 1.75 ;
      RECT  2.93 1.21 3.05 1.75 ;
      RECT  3.445 1.45 3.575 1.75 ;
      RECT  3.98 1.45 4.11 1.75 ;
      RECT  4.5 1.45 4.63 1.75 ;
      RECT  5.02 1.44 5.15 1.75 ;
      RECT  5.54 1.44 5.67 1.75 ;
      RECT  6.06 1.44 6.19 1.75 ;
      RECT  6.58 1.44 6.71 1.75 ;
      RECT  7.1 1.44 7.23 1.75 ;
      RECT  7.62 1.44 7.75 1.75 ;
      RECT  8.14 1.44 8.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  2.11 0.05 2.28 0.22 ;
      RECT  5.52 0.05 5.69 0.325 ;
      RECT  6.04 0.05 6.21 0.325 ;
      RECT  6.56 0.05 6.73 0.325 ;
      RECT  7.08 0.05 7.25 0.325 ;
      RECT  7.6 0.05 7.77 0.325 ;
      RECT  8.12 0.05 8.29 0.325 ;
      RECT  0.325 0.05 0.455 0.35 ;
      RECT  3.445 0.05 3.575 0.35 ;
      RECT  2.925 0.05 3.055 0.415 ;
      RECT  1.315 0.05 1.445 0.46 ;
      RECT  5.0 0.05 5.12 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.705 0.14 1.91 0.31 ;
      RECT  1.82 0.31 2.525 0.4 ;
      RECT  2.435 0.4 2.525 0.835 ;
      RECT  2.435 0.835 2.88 0.925 ;
      RECT  2.78 0.735 2.88 0.835 ;
      RECT  2.435 0.925 2.54 1.255 ;
      RECT  1.36 1.255 2.54 1.3 ;
      RECT  0.98 1.3 2.54 1.345 ;
      RECT  0.98 1.345 1.45 1.39 ;
      RECT  0.98 1.39 1.07 1.605 ;
      RECT  3.71 0.24 4.415 0.36 ;
      RECT  3.71 0.36 3.83 0.44 ;
      RECT  3.15 0.44 3.83 0.56 ;
      RECT  0.07 0.34 0.19 0.44 ;
      RECT  0.07 0.44 0.76 0.56 ;
      RECT  0.85 0.375 0.97 0.55 ;
      RECT  0.85 0.55 1.54 0.675 ;
      RECT  1.45 0.675 1.54 0.825 ;
      RECT  0.85 0.675 0.96 1.09 ;
      RECT  0.765 1.09 0.96 1.21 ;
      RECT  3.935 0.45 4.625 0.57 ;
      RECT  4.505 0.57 4.625 0.725 ;
      RECT  4.505 0.725 7.22 0.84 ;
      RECT  4.505 0.84 4.625 1.24 ;
      RECT  3.165 1.24 4.625 1.36 ;
      RECT  2.625 0.505 3.06 0.625 ;
      RECT  2.97 0.625 3.06 0.74 ;
      RECT  2.97 0.74 3.635 0.85 ;
      RECT  2.97 0.85 3.06 1.015 ;
      RECT  2.67 1.015 3.06 1.105 ;
      RECT  2.67 1.105 2.79 1.435 ;
      RECT  1.61 1.435 2.79 1.525 ;
      RECT  1.61 1.525 1.7 1.66 ;
      RECT  3.83 0.785 4.365 0.89 ;
      RECT  3.83 0.89 3.925 0.95 ;
      RECT  3.29 0.95 3.925 1.05 ;
      RECT  1.215 0.765 1.31 0.915 ;
      RECT  1.215 0.915 1.74 1.005 ;
      RECT  1.63 0.445 1.74 0.915 ;
      RECT  1.635 1.005 1.74 1.16 ;
      RECT  1.865 0.52 1.985 1.16 ;
      LAYER M2 ;
      RECT  1.83 0.95 3.47 1.05 ;
      LAYER V1 ;
      RECT  1.87 0.95 1.97 1.05 ;
      RECT  3.33 0.95 3.43 1.05 ;
  END
END SEN_CKGTPLT_16
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLT_2
#      Description : "Clock Gater, positive clock, synchronous enable, pre control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLT_2
  CLASS CORE ;
  FOREIGN SEN_CKGTPLT_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.91 2.45 1.095 ;
      RECT  2.15 1.095 2.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0354 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0354 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.22 4.25 1.11 ;
      RECT  3.805 1.11 4.545 1.32 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0432 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  1.37 1.395 1.5 1.75 ;
      RECT  2.215 1.57 2.345 1.75 ;
      RECT  2.975 1.41 3.105 1.75 ;
      RECT  3.525 1.41 3.655 1.75 ;
      RECT  4.11 1.41 4.24 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.215 0.05 2.345 0.215 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  3.875 0.05 4.005 0.39 ;
      RECT  4.395 0.05 4.525 0.39 ;
      RECT  3.195 0.05 3.325 0.395 ;
      RECT  1.36 0.05 1.49 0.46 ;
      RECT  2.72 0.05 2.83 0.48 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.755 0.14 1.855 0.305 ;
      RECT  1.755 0.305 2.63 0.42 ;
      RECT  2.54 0.42 2.63 0.765 ;
      RECT  2.54 0.765 2.915 0.875 ;
      RECT  2.81 0.64 2.915 0.765 ;
      RECT  2.54 0.875 2.63 1.26 ;
      RECT  2.49 1.26 2.63 1.38 ;
      RECT  1.755 1.38 2.63 1.47 ;
      RECT  1.755 1.47 1.865 1.66 ;
      RECT  2.97 0.285 3.095 0.46 ;
      RECT  3.005 0.46 3.095 0.83 ;
      RECT  3.005 0.83 3.255 0.94 ;
      RECT  3.005 0.94 3.095 1.0 ;
      RECT  2.72 1.0 3.095 1.09 ;
      RECT  2.72 1.09 2.84 1.51 ;
      RECT  0.065 0.28 0.185 0.48 ;
      RECT  0.065 0.48 0.705 0.57 ;
      RECT  0.585 0.24 0.705 0.48 ;
      RECT  1.945 0.545 2.45 0.655 ;
      RECT  1.945 0.655 2.06 1.275 ;
      RECT  3.185 0.51 3.535 0.69 ;
      RECT  3.43 0.69 3.535 1.035 ;
      RECT  0.79 0.6 1.625 0.72 ;
      RECT  1.525 0.72 1.625 1.03 ;
      RECT  0.79 0.72 0.88 1.44 ;
      RECT  0.79 1.44 1.01 1.56 ;
      RECT  3.625 0.32 3.77 0.745 ;
      RECT  3.625 0.745 4.06 0.855 ;
      RECT  3.625 0.855 3.715 1.19 ;
      RECT  3.18 1.19 3.715 1.31 ;
      RECT  1.215 0.89 1.435 1.0 ;
      RECT  1.345 1.0 1.435 1.17 ;
      RECT  1.345 1.17 1.82 1.29 ;
      RECT  1.715 0.53 1.82 1.17 ;
      RECT  0.97 0.88 1.075 1.18 ;
      RECT  0.97 1.18 1.25 1.27 ;
      RECT  1.15 1.27 1.25 1.51 ;
      LAYER M2 ;
      RECT  2.27 0.55 3.325 0.65 ;
      RECT  1.11 1.35 2.86 1.45 ;
      LAYER V1 ;
      RECT  2.31 0.55 2.41 0.65 ;
      RECT  3.185 0.55 3.285 0.65 ;
      RECT  1.15 1.35 1.25 1.45 ;
      RECT  2.72 1.35 2.82 1.45 ;
  END
END SEN_CKGTPLT_2
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLT_3
#      Description : "Clock Gater, positive clock, synchronous enable, pre control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLT_3
  CLASS CORE ;
  FOREIGN SEN_CKGTPLT_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.76 ;
      RECT  2.15 0.76 2.33 0.94 ;
      RECT  2.15 0.94 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.31 4.05 1.11 ;
      RECT  3.55 1.11 4.33 1.29 ;
    END
    ANTENNADIFFAREA 0.298 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.11 ;
      RECT  0.15 1.11 0.255 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0459 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  1.35 1.205 1.475 1.75 ;
      RECT  2.105 1.56 2.235 1.75 ;
      RECT  2.84 1.215 2.955 1.75 ;
      RECT  3.385 1.41 3.515 1.75 ;
      RECT  3.935 1.41 4.065 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  2.085 0.05 2.255 0.19 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  1.345 0.05 1.475 0.565 ;
      RECT  2.905 0.05 3.025 0.59 ;
      RECT  3.675 0.05 3.8 0.59 ;
      RECT  4.21 0.05 4.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.75 0.14 1.86 0.28 ;
      RECT  1.75 0.28 2.56 0.39 ;
      RECT  2.46 0.39 2.56 1.11 ;
      RECT  2.355 1.11 2.56 1.23 ;
      RECT  2.355 1.23 2.445 1.38 ;
      RECT  1.865 1.38 2.445 1.47 ;
      RECT  1.865 1.47 1.955 1.55 ;
      RECT  1.67 1.55 1.955 1.66 ;
      RECT  0.065 0.3 0.185 0.485 ;
      RECT  0.065 0.485 0.705 0.575 ;
      RECT  0.585 0.24 0.705 0.485 ;
      RECT  3.115 0.44 3.585 0.56 ;
      RECT  3.495 0.56 3.585 0.735 ;
      RECT  3.115 0.56 3.21 1.285 ;
      RECT  3.495 0.735 3.84 0.845 ;
      RECT  1.585 0.48 1.755 0.59 ;
      RECT  1.665 0.59 1.755 1.025 ;
      RECT  1.2 0.845 1.31 1.025 ;
      RECT  1.2 1.025 1.755 1.115 ;
      RECT  1.61 1.115 1.755 1.34 ;
      RECT  0.855 0.41 0.98 0.665 ;
      RECT  0.75 0.665 1.535 0.755 ;
      RECT  1.435 0.755 1.535 0.925 ;
      RECT  0.75 0.755 0.84 1.415 ;
      RECT  0.75 1.415 1.02 1.535 ;
      RECT  2.65 0.24 2.755 0.76 ;
      RECT  2.65 0.76 2.995 0.87 ;
      RECT  2.65 0.87 2.75 1.44 ;
      RECT  2.54 1.44 2.75 1.56 ;
      RECT  0.945 0.845 1.045 1.235 ;
      RECT  0.945 1.235 1.25 1.325 ;
      RECT  1.15 1.325 1.25 1.51 ;
      RECT  1.845 0.48 1.96 1.29 ;
      RECT  3.3 0.73 3.405 1.29 ;
      LAYER M2 ;
      RECT  1.82 1.15 3.44 1.25 ;
      RECT  1.11 1.35 2.79 1.45 ;
      LAYER V1 ;
      RECT  1.86 1.15 1.96 1.25 ;
      RECT  3.3 1.15 3.4 1.25 ;
      RECT  1.15 1.35 1.25 1.45 ;
      RECT  2.65 1.35 2.75 1.45 ;
  END
END SEN_CKGTPLT_3
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLT_4
#      Description : "Clock Gater, positive clock, synchronous enable, pre control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLT_4
  CLASS CORE ;
  FOREIGN SEN_CKGTPLT_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.75 ;
      RECT  2.15 0.75 2.34 0.93 ;
      RECT  2.15 0.93 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0387 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0387 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.89 0.31 4.05 0.485 ;
      RECT  3.89 0.485 4.53 0.575 ;
      RECT  4.41 0.31 4.53 0.485 ;
      RECT  4.15 0.575 4.26 1.11 ;
      RECT  3.55 1.11 4.26 1.29 ;
    END
    ANTENNADIFFAREA 0.363 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.11 ;
      RECT  0.15 1.11 0.255 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0477 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  1.35 1.245 1.47 1.75 ;
      RECT  2.105 1.565 2.235 1.75 ;
      RECT  2.84 1.21 2.955 1.75 ;
      RECT  3.36 1.41 3.49 1.75 ;
      RECT  3.885 1.41 4.015 1.75 ;
      RECT  4.41 1.21 4.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.085 0.05 2.255 0.2 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  3.625 0.05 3.755 0.385 ;
      RECT  4.145 0.05 4.275 0.385 ;
      RECT  1.345 0.05 1.475 0.59 ;
      RECT  2.905 0.05 3.025 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.69 0.14 1.8 0.29 ;
      RECT  1.69 0.29 2.56 0.39 ;
      RECT  2.46 0.39 2.56 1.155 ;
      RECT  2.345 1.155 2.56 1.275 ;
      RECT  2.345 1.275 2.435 1.38 ;
      RECT  1.865 1.38 2.435 1.47 ;
      RECT  1.865 1.47 1.955 1.57 ;
      RECT  1.67 1.57 1.955 1.66 ;
      RECT  0.065 0.31 0.185 0.485 ;
      RECT  0.065 0.485 0.705 0.575 ;
      RECT  0.585 0.26 0.705 0.485 ;
      RECT  1.585 0.48 1.755 0.6 ;
      RECT  1.665 0.6 1.755 1.065 ;
      RECT  1.2 0.87 1.31 1.065 ;
      RECT  1.2 1.065 1.755 1.155 ;
      RECT  1.61 1.155 1.755 1.39 ;
      RECT  3.115 0.485 3.7 0.605 ;
      RECT  3.61 0.605 3.7 0.72 ;
      RECT  3.115 0.605 3.21 1.21 ;
      RECT  3.61 0.72 4.05 0.83 ;
      RECT  0.86 0.41 0.98 0.69 ;
      RECT  0.75 0.69 1.565 0.78 ;
      RECT  1.465 0.78 1.565 0.945 ;
      RECT  0.75 0.78 0.84 1.445 ;
      RECT  0.75 1.445 1.02 1.565 ;
      RECT  2.65 0.26 2.755 0.815 ;
      RECT  2.65 0.815 3.025 0.915 ;
      RECT  2.65 0.915 2.75 1.44 ;
      RECT  2.54 1.44 2.75 1.56 ;
      RECT  0.97 0.87 1.08 1.255 ;
      RECT  0.97 1.255 1.25 1.345 ;
      RECT  1.15 1.345 1.25 1.51 ;
      RECT  1.845 0.48 1.96 1.29 ;
      RECT  3.3 0.725 3.405 1.29 ;
      LAYER M2 ;
      RECT  1.82 1.15 3.44 1.25 ;
      RECT  1.11 1.35 2.79 1.45 ;
      LAYER V1 ;
      RECT  1.86 1.15 1.96 1.25 ;
      RECT  3.3 1.15 3.4 1.25 ;
      RECT  1.15 1.35 1.25 1.45 ;
      RECT  2.65 1.35 2.75 1.45 ;
  END
END SEN_CKGTPLT_4
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLT_6
#      Description : "Clock Gater, positive clock, synchronous enable, pre control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLT_6
  CLASS CORE ;
  FOREIGN SEN_CKGTPLT_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  2.15 0.71 2.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0399 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.91 ;
      RECT  0.55 0.91 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0399 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.7 0.445 5.45 0.565 ;
      RECT  5.32 0.565 5.45 1.11 ;
      RECT  4.15 1.11 5.45 1.29 ;
    END
    ANTENNADIFFAREA 0.512 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0501 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  1.34 1.24 1.47 1.75 ;
      RECT  2.1 1.56 2.23 1.75 ;
      RECT  2.9 1.2 3.005 1.75 ;
      RECT  3.39 1.59 3.56 1.75 ;
      RECT  3.945 1.215 4.06 1.75 ;
      RECT  4.46 1.41 4.59 1.75 ;
      RECT  5.0 1.41 5.13 1.75 ;
      RECT  5.56 1.21 5.68 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  2.1 0.05 2.23 0.225 ;
      RECT  5.0 0.05 5.13 0.355 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  2.6 0.05 2.73 0.39 ;
      RECT  3.405 0.05 3.535 0.39 ;
      RECT  1.34 0.05 1.47 0.575 ;
      RECT  4.465 0.05 4.585 0.59 ;
      RECT  5.58 0.05 5.7 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.685 0.14 4.325 0.23 ;
      RECT  4.205 0.23 4.325 0.43 ;
      RECT  3.685 0.23 3.805 0.5 ;
      RECT  3.135 0.26 3.255 0.5 ;
      RECT  3.135 0.5 3.805 0.59 ;
      RECT  1.66 0.15 1.96 0.25 ;
      RECT  1.87 0.25 1.96 0.315 ;
      RECT  1.87 0.315 2.455 0.405 ;
      RECT  2.335 0.19 2.455 0.315 ;
      RECT  2.34 0.405 2.455 0.51 ;
      RECT  2.34 0.51 2.63 0.6 ;
      RECT  2.54 0.6 2.63 0.78 ;
      RECT  2.54 0.78 2.865 0.89 ;
      RECT  2.54 0.89 2.63 1.095 ;
      RECT  2.21 1.095 2.63 1.215 ;
      RECT  2.21 1.215 2.3 1.38 ;
      RECT  1.835 1.38 2.3 1.47 ;
      RECT  1.835 1.47 1.925 1.545 ;
      RECT  1.665 1.545 1.925 1.66 ;
      RECT  2.85 0.24 3.045 0.36 ;
      RECT  2.955 0.36 3.045 0.785 ;
      RECT  2.955 0.785 3.31 0.895 ;
      RECT  2.955 0.895 3.045 1.02 ;
      RECT  2.72 1.02 3.045 1.11 ;
      RECT  2.72 1.11 2.81 1.34 ;
      RECT  2.39 1.34 2.81 1.46 ;
      RECT  0.065 0.33 0.185 0.485 ;
      RECT  0.065 0.485 0.705 0.575 ;
      RECT  0.585 0.26 0.705 0.485 ;
      RECT  0.855 0.37 0.975 0.665 ;
      RECT  0.78 0.665 1.53 0.755 ;
      RECT  1.43 0.755 1.53 0.97 ;
      RECT  0.78 0.755 0.87 1.44 ;
      RECT  0.78 1.44 1.02 1.56 ;
      RECT  3.945 0.32 4.065 0.755 ;
      RECT  3.945 0.755 5.21 0.865 ;
      RECT  3.945 0.865 4.06 1.02 ;
      RECT  3.685 1.02 4.06 1.11 ;
      RECT  3.685 1.11 3.805 1.38 ;
      RECT  3.12 1.38 3.805 1.5 ;
      RECT  3.4 0.81 3.84 0.915 ;
      RECT  3.4 0.915 3.5 1.29 ;
      RECT  1.2 0.845 1.3 1.06 ;
      RECT  1.2 1.06 1.725 1.15 ;
      RECT  1.62 0.41 1.725 1.06 ;
      RECT  1.605 1.15 1.725 1.39 ;
      RECT  0.965 0.845 1.075 1.25 ;
      RECT  0.965 1.25 1.25 1.34 ;
      RECT  1.15 1.34 1.25 1.51 ;
      RECT  1.835 0.5 1.955 1.29 ;
      LAYER M2 ;
      RECT  1.815 1.15 3.54 1.25 ;
      RECT  1.11 1.35 2.57 1.45 ;
      LAYER V1 ;
      RECT  1.855 1.15 1.955 1.25 ;
      RECT  3.4 1.15 3.5 1.25 ;
      RECT  1.15 1.35 1.25 1.45 ;
      RECT  2.43 1.35 2.53 1.45 ;
  END
END SEN_CKGTPLT_6
#-----------------------------------------------------------------------
#      Cell        : SEN_CKGTPLT_8
#      Description : "Clock Gater, positive clock, synchronous enable, pre control"
#      Equation    : iq,iqn=latch(enable=!CK,data_in=EN|SE):Q=CK&iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CKGTPLT_8
  CLASS CORE ;
  FOREIGN SEN_CKGTPLT_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  2.15 0.71 2.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0537 ;
  END CK
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0537 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.74 0.29 4.85 0.425 ;
      RECT  4.74 0.425 5.91 0.545 ;
      RECT  5.48 0.545 5.65 1.11 ;
      RECT  4.15 1.11 6.05 1.29 ;
    END
    ANTENNADIFFAREA 0.684 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  1.345 1.24 1.465 1.75 ;
      RECT  2.1 1.56 2.23 1.75 ;
      RECT  2.9 1.2 3.005 1.75 ;
      RECT  3.39 1.59 3.56 1.75 ;
      RECT  3.945 1.235 4.06 1.75 ;
      RECT  4.46 1.41 4.59 1.75 ;
      RECT  4.98 1.41 5.11 1.75 ;
      RECT  5.5 1.41 5.63 1.75 ;
      RECT  6.02 1.41 6.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  2.1 0.05 2.23 0.225 ;
      RECT  4.96 0.05 5.13 0.335 ;
      RECT  5.48 0.05 5.65 0.335 ;
      RECT  3.405 0.05 3.535 0.385 ;
      RECT  2.6 0.05 2.73 0.39 ;
      RECT  4.46 0.05 4.59 0.39 ;
      RECT  6.02 0.05 6.145 0.39 ;
      RECT  0.32 0.05 0.45 0.41 ;
      RECT  1.34 0.05 1.47 0.57 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.65 0.145 1.96 0.255 ;
      RECT  1.87 0.255 1.96 0.315 ;
      RECT  1.87 0.315 2.455 0.41 ;
      RECT  2.34 0.41 2.455 0.51 ;
      RECT  2.34 0.51 2.63 0.6 ;
      RECT  2.54 0.6 2.63 0.78 ;
      RECT  2.54 0.78 2.865 0.89 ;
      RECT  2.54 0.89 2.63 1.04 ;
      RECT  2.21 1.04 2.63 1.16 ;
      RECT  2.21 1.16 2.3 1.38 ;
      RECT  1.835 1.38 2.3 1.47 ;
      RECT  1.835 1.47 1.925 1.545 ;
      RECT  1.65 1.545 1.925 1.655 ;
      RECT  3.685 0.215 4.37 0.335 ;
      RECT  3.685 0.335 3.805 0.475 ;
      RECT  3.135 0.34 3.255 0.475 ;
      RECT  3.135 0.475 3.805 0.565 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.59 ;
      RECT  0.585 0.37 0.705 0.5 ;
      RECT  2.82 0.44 3.045 0.56 ;
      RECT  2.955 0.56 3.045 0.655 ;
      RECT  2.955 0.655 3.4 0.76 ;
      RECT  2.955 0.76 3.045 1.02 ;
      RECT  2.72 1.02 3.045 1.11 ;
      RECT  2.72 1.11 2.81 1.34 ;
      RECT  2.39 1.34 2.81 1.46 ;
      RECT  0.845 0.41 0.965 0.66 ;
      RECT  0.78 0.66 1.53 0.75 ;
      RECT  1.43 0.75 1.53 0.97 ;
      RECT  0.78 0.75 0.87 1.44 ;
      RECT  0.78 1.44 1.02 1.56 ;
      RECT  3.945 0.425 4.065 0.73 ;
      RECT  3.945 0.73 5.375 0.84 ;
      RECT  3.945 0.84 4.06 1.055 ;
      RECT  3.685 1.055 4.06 1.145 ;
      RECT  3.685 1.145 3.805 1.38 ;
      RECT  3.12 1.38 3.805 1.5 ;
      RECT  3.4 0.86 3.83 0.965 ;
      RECT  3.4 0.965 3.5 1.29 ;
      RECT  1.2 0.845 1.3 1.06 ;
      RECT  1.2 1.06 1.725 1.15 ;
      RECT  1.62 0.42 1.725 1.06 ;
      RECT  1.605 1.15 1.725 1.39 ;
      RECT  0.96 0.845 1.065 1.24 ;
      RECT  0.96 1.24 1.25 1.33 ;
      RECT  1.15 1.33 1.25 1.51 ;
      RECT  1.835 0.51 1.955 1.29 ;
      LAYER M2 ;
      RECT  1.815 1.15 3.54 1.25 ;
      RECT  1.11 1.35 2.57 1.45 ;
      LAYER V1 ;
      RECT  1.855 1.15 1.955 1.25 ;
      RECT  3.4 1.15 3.5 1.25 ;
      RECT  1.15 1.35 1.25 1.45 ;
      RECT  2.43 1.35 2.53 1.45 ;
  END
END SEN_CKGTPLT_8
#-----------------------------------------------------------------------
#      Cell        : SEN_DEL_L4_1
#      Description : "Delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DEL_L4_1
  CLASS CORE ;
  FOREIGN SEN_DEL_L4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.295 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.19 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.235 1.175 1.355 1.75 ;
      RECT  2.14 1.0 2.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.235 0.05 1.355 0.6 ;
      RECT  0.065 0.05 0.19 0.62 ;
      RECT  2.14 0.05 2.26 0.68 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.225 2.545 0.395 ;
      RECT  2.35 0.395 2.45 1.015 ;
      RECT  2.35 1.015 2.545 1.19 ;
    END
    ANTENNADIFFAREA 0.141 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.5 0.215 1.08 0.335 ;
      RECT  0.99 0.335 1.08 0.785 ;
      RECT  0.99 0.785 1.81 0.895 ;
      RECT  0.99 0.895 1.08 1.42 ;
      RECT  0.42 1.42 1.08 1.54 ;
      RECT  0.335 0.465 0.455 0.675 ;
      RECT  0.365 0.675 0.455 0.785 ;
      RECT  0.365 0.785 0.9 0.895 ;
      RECT  0.365 0.895 0.455 1.0 ;
      RECT  0.34 1.0 0.455 1.225 ;
      RECT  1.92 0.2 2.04 0.78 ;
      RECT  1.92 0.78 2.24 0.89 ;
      RECT  1.92 0.89 2.04 1.59 ;
  END
END SEN_DEL_L4_1
#-----------------------------------------------------------------------
#      Cell        : SEN_DEL_L4_2
#      Description : "Delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DEL_L4_2
  CLASS CORE ;
  FOREIGN SEN_DEL_L4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 2.8 1.85 ;
      RECT  1.17 1.2 1.29 1.75 ;
      RECT  2.105 1.2 2.225 1.75 ;
      RECT  2.62 1.4 2.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      RECT  2.62 0.05 2.745 0.4 ;
      RECT  0.065 0.05 0.19 0.6 ;
      RECT  1.17 0.05 1.29 0.6 ;
      RECT  2.105 0.05 2.225 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.31 2.485 0.485 ;
      RECT  2.35 0.485 2.45 1.315 ;
      RECT  2.35 1.315 2.485 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.41 0.215 1.05 0.335 ;
      RECT  0.96 0.335 1.05 0.73 ;
      RECT  0.96 0.73 1.7 0.9 ;
      RECT  0.96 0.9 1.05 1.285 ;
      RECT  0.485 1.285 1.05 1.375 ;
      RECT  0.485 1.375 0.605 1.63 ;
      RECT  1.855 0.23 1.975 0.73 ;
      RECT  1.855 0.73 2.26 0.9 ;
      RECT  1.855 0.9 1.975 1.555 ;
      RECT  0.34 0.5 0.455 0.785 ;
      RECT  0.34 0.785 0.87 0.895 ;
      RECT  0.34 0.895 0.455 1.2 ;
  END
END SEN_DEL_L4_2
#-----------------------------------------------------------------------
#      Cell        : SEN_DEL_L4_4
#      Description : "Delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DEL_L4_4
  CLASS CORE ;
  FOREIGN SEN_DEL_L4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  1.195 1.21 1.315 1.75 ;
      RECT  2.13 1.21 2.25 1.75 ;
      RECT  2.645 1.41 2.775 1.75 ;
      RECT  3.18 1.21 3.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  2.645 0.05 2.775 0.39 ;
      RECT  3.18 0.05 3.3 0.59 ;
      RECT  1.195 0.05 1.315 0.6 ;
      RECT  2.13 0.05 2.25 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 3.05 0.69 ;
      RECT  2.95 0.69 3.05 1.11 ;
      RECT  2.35 1.11 3.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.46 0.215 1.08 0.335 ;
      RECT  0.99 0.335 1.08 0.78 ;
      RECT  0.99 0.78 1.78 0.9 ;
      RECT  0.99 0.9 1.08 1.465 ;
      RECT  0.46 1.465 1.08 1.585 ;
      RECT  0.34 0.49 0.455 0.78 ;
      RECT  0.34 0.78 0.9 0.9 ;
      RECT  0.34 0.9 0.455 1.305 ;
      RECT  1.88 0.32 2.0 0.78 ;
      RECT  1.88 0.78 2.84 0.9 ;
      RECT  1.88 0.9 2.0 1.4 ;
  END
END SEN_DEL_L4_4
#-----------------------------------------------------------------------
#      Cell        : SEN_DEL_L4_8
#      Description : "Delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DEL_L4_8
  CLASS CORE ;
  FOREIGN SEN_DEL_L4_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.455 1.21 1.575 1.75 ;
      RECT  2.32 1.41 2.45 1.75 ;
      RECT  2.84 1.41 2.97 1.75 ;
      RECT  3.36 1.41 3.49 1.75 ;
      RECT  3.88 1.41 4.01 1.75 ;
      RECT  4.41 1.21 4.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.84 0.05 2.97 0.38 ;
      RECT  3.36 0.05 3.49 0.38 ;
      RECT  3.88 0.05 4.01 0.38 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.535 0.05 0.655 0.51 ;
      RECT  4.41 0.05 4.53 0.59 ;
      RECT  1.455 0.05 1.575 0.6 ;
      RECT  2.34 0.05 2.445 0.68 ;
      RECT  0.535 0.51 0.76 0.63 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 4.25 0.69 ;
      RECT  4.15 0.69 4.25 1.11 ;
      RECT  2.55 1.11 4.25 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.745 0.235 1.33 0.355 ;
      RECT  1.24 0.355 1.33 0.785 ;
      RECT  1.24 0.785 2.015 0.895 ;
      RECT  1.24 0.895 1.33 1.04 ;
      RECT  0.72 1.04 1.33 1.16 ;
      RECT  0.34 0.315 0.445 0.785 ;
      RECT  0.34 0.785 1.135 0.895 ;
      RECT  0.34 0.895 0.445 1.285 ;
      RECT  2.14 0.18 2.25 0.785 ;
      RECT  2.14 0.785 3.765 0.895 ;
      RECT  2.14 0.895 2.26 1.23 ;
  END
END SEN_DEL_L4_8
#-----------------------------------------------------------------------
#      Cell        : SEN_DEL_L6_1
#      Description : "Delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DEL_L6_1
  CLASS CORE ;
  FOREIGN SEN_DEL_L6_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  1.235 1.175 1.355 1.75 ;
      RECT  2.85 1.175 2.97 1.75 ;
      RECT  3.765 1.0 3.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  3.73 0.05 3.855 0.41 ;
      RECT  1.235 0.05 1.355 0.6 ;
      RECT  2.85 0.05 2.97 0.6 ;
      RECT  0.065 0.05 0.19 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.31 4.135 0.49 ;
      RECT  3.95 0.49 4.05 1.115 ;
      RECT  3.95 1.115 4.135 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.55 0.2 0.67 0.335 ;
      RECT  0.55 0.335 1.14 0.425 ;
      RECT  1.05 0.425 1.14 0.76 ;
      RECT  1.05 0.76 1.81 0.87 ;
      RECT  1.05 0.87 1.14 1.37 ;
      RECT  0.495 1.37 1.14 1.49 ;
      RECT  2.115 0.24 2.64 0.36 ;
      RECT  2.55 0.36 2.64 0.785 ;
      RECT  2.55 0.785 3.425 0.895 ;
      RECT  2.55 0.895 2.64 1.055 ;
      RECT  2.13 1.055 2.64 1.175 ;
      RECT  1.92 0.425 2.04 0.78 ;
      RECT  1.92 0.78 2.45 0.89 ;
      RECT  1.92 0.89 2.04 1.585 ;
      RECT  0.34 0.425 0.455 0.785 ;
      RECT  0.34 0.785 0.96 0.895 ;
      RECT  0.34 0.895 0.455 1.23 ;
      RECT  3.535 0.475 3.655 0.79 ;
      RECT  3.535 0.79 3.84 0.9 ;
      RECT  3.535 0.9 3.655 1.59 ;
  END
END SEN_DEL_L6_1
#-----------------------------------------------------------------------
#      Cell        : SEN_DEL_L6_2
#      Description : "Delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DEL_L6_2
  CLASS CORE ;
  FOREIGN SEN_DEL_L6_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  1.205 1.175 1.325 1.75 ;
      RECT  2.73 1.37 2.86 1.75 ;
      RECT  3.695 1.21 3.815 1.75 ;
      RECT  4.215 1.21 4.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  2.73 0.05 2.86 0.4 ;
      RECT  3.695 0.05 3.815 0.59 ;
      RECT  4.215 0.05 4.335 0.59 ;
      RECT  0.06 0.05 0.19 0.6 ;
      RECT  1.205 0.05 1.325 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.31 4.075 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.415 0.215 1.04 0.335 ;
      RECT  0.95 0.335 1.04 0.785 ;
      RECT  0.95 0.785 1.75 0.895 ;
      RECT  0.95 0.895 1.04 1.31 ;
      RECT  0.47 1.31 1.04 1.43 ;
      RECT  1.845 0.215 2.065 0.335 ;
      RECT  1.845 0.335 1.935 0.795 ;
      RECT  1.845 0.795 2.61 0.905 ;
      RECT  1.845 0.905 1.935 1.455 ;
      RECT  1.845 1.455 2.06 1.575 ;
      RECT  2.025 0.545 2.81 0.665 ;
      RECT  2.72 0.665 2.81 0.76 ;
      RECT  2.72 0.76 3.31 0.87 ;
      RECT  2.72 0.87 2.81 1.015 ;
      RECT  2.025 1.015 2.81 1.135 ;
      RECT  0.34 0.485 0.445 0.785 ;
      RECT  0.34 0.785 0.855 0.895 ;
      RECT  0.34 0.895 0.445 1.195 ;
      RECT  3.42 0.23 3.54 0.785 ;
      RECT  3.42 0.785 3.86 0.895 ;
      RECT  3.42 0.895 3.54 1.53 ;
  END
END SEN_DEL_L6_2
#-----------------------------------------------------------------------
#      Cell        : SEN_DEL_L6_4
#      Description : "Delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DEL_L6_4
  CLASS CORE ;
  FOREIGN SEN_DEL_L6_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.195 1.19 1.315 1.75 ;
      RECT  2.75 1.175 2.87 1.75 ;
      RECT  3.735 1.18 3.855 1.75 ;
      RECT  4.265 1.4 4.395 1.75 ;
      RECT  4.79 1.21 4.91 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  4.265 0.05 4.395 0.38 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  3.75 0.05 3.87 0.59 ;
      RECT  4.79 0.05 4.91 0.59 ;
      RECT  1.195 0.05 1.315 0.6 ;
      RECT  2.75 0.05 2.87 0.615 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.01 0.51 4.65 0.69 ;
      RECT  4.55 0.69 4.65 1.11 ;
      RECT  3.95 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.46 0.215 1.09 0.335 ;
      RECT  1.0 0.335 1.09 0.785 ;
      RECT  1.0 0.785 1.77 0.895 ;
      RECT  1.0 0.895 1.09 1.465 ;
      RECT  0.46 1.465 1.09 1.585 ;
      RECT  2.015 0.215 2.66 0.335 ;
      RECT  2.57 0.335 2.66 0.785 ;
      RECT  2.57 0.785 3.33 0.895 ;
      RECT  2.57 0.895 2.66 1.18 ;
      RECT  2.04 1.18 2.66 1.3 ;
      RECT  0.34 0.46 0.445 0.785 ;
      RECT  0.34 0.785 0.91 0.895 ;
      RECT  0.34 0.895 0.455 1.19 ;
      RECT  1.86 0.495 2.0 0.785 ;
      RECT  1.86 0.785 2.48 0.895 ;
      RECT  1.86 0.895 1.95 1.44 ;
      RECT  1.86 1.44 2.0 1.61 ;
      RECT  3.435 0.32 3.555 0.785 ;
      RECT  3.435 0.785 4.44 0.895 ;
      RECT  3.435 0.895 3.555 1.42 ;
  END
END SEN_DEL_L6_4
#-----------------------------------------------------------------------
#      Cell        : SEN_DEL_L6_8
#      Description : "Delay buffer"
#      Equation    : X=A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DEL_L6_8
  CLASS CORE ;
  FOREIGN SEN_DEL_L6_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.455 1.19 1.575 1.75 ;
      RECT  3.01 1.19 3.13 1.75 ;
      RECT  3.945 1.2 4.06 1.75 ;
      RECT  4.46 1.41 4.59 1.75 ;
      RECT  4.98 1.41 5.11 1.75 ;
      RECT  5.5 1.41 5.63 1.75 ;
      RECT  6.02 1.41 6.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  0.58 0.05 0.71 0.375 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  4.46 0.05 4.59 0.39 ;
      RECT  4.98 0.05 5.11 0.39 ;
      RECT  5.5 0.05 5.63 0.39 ;
      RECT  6.02 0.05 6.145 0.39 ;
      RECT  3.945 0.05 4.06 0.605 ;
      RECT  1.455 0.05 1.575 0.61 ;
      RECT  3.01 0.05 3.13 0.64 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.51 5.885 0.69 ;
      RECT  5.715 0.69 5.885 1.11 ;
      RECT  4.15 1.11 5.885 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.09 0.21 2.26 0.38 ;
      RECT  2.09 0.38 2.19 0.785 ;
      RECT  2.09 0.785 2.74 0.895 ;
      RECT  2.09 0.895 2.19 1.465 ;
      RECT  2.09 1.465 2.31 1.585 ;
      RECT  0.72 0.515 1.365 0.635 ;
      RECT  1.275 0.635 1.365 0.785 ;
      RECT  1.275 0.785 1.985 0.895 ;
      RECT  1.275 0.895 1.365 1.04 ;
      RECT  0.72 1.04 1.365 1.16 ;
      RECT  2.285 0.515 2.92 0.635 ;
      RECT  2.83 0.635 2.92 0.785 ;
      RECT  2.83 0.785 3.58 0.895 ;
      RECT  2.83 0.895 2.92 1.04 ;
      RECT  2.3 1.04 2.92 1.16 ;
      RECT  0.34 0.45 0.445 0.785 ;
      RECT  0.34 0.785 1.185 0.895 ;
      RECT  0.34 0.895 0.445 1.23 ;
      RECT  3.695 0.42 3.815 0.785 ;
      RECT  3.695 0.785 5.6 0.895 ;
      RECT  3.695 0.895 3.815 1.26 ;
  END
END SEN_DEL_L6_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_0P5
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_0P5
  CLASS CORE ;
  FOREIGN SEN_EN2_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.2 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.815 ;
      RECT  1.35 0.815 1.515 0.985 ;
      RECT  1.35 0.985 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.34 0.175 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.215 1.615 1.385 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.235 0.05 1.405 0.42 ;
      RECT  0.055 0.05 0.175 0.49 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.335 0.685 1.455 ;
    END
    ANTENNADIFFAREA 0.102 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.39 0.14 0.87 0.23 ;
      RECT  0.775 0.23 0.87 1.435 ;
      RECT  0.775 1.435 1.725 1.525 ;
      RECT  1.605 0.26 1.725 1.435 ;
      RECT  0.775 1.525 0.87 1.57 ;
      RECT  0.65 1.57 0.87 1.66 ;
      RECT  0.315 0.335 0.44 0.505 ;
      RECT  0.34 0.505 0.44 1.285 ;
      RECT  0.315 1.285 0.44 1.455 ;
      RECT  1.16 0.57 1.26 1.29 ;
      RECT  0.96 0.31 1.07 1.345 ;
      LAYER M2 ;
      RECT  0.3 1.15 1.3 1.25 ;
      LAYER V1 ;
      RECT  0.34 1.15 0.44 1.25 ;
      RECT  1.16 1.15 1.26 1.25 ;
  END
END SEN_EN2_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_1
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_1
  CLASS CORE ;
  FOREIGN SEN_EN2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.71 0.45 0.97 ;
      RECT  0.35 0.97 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 1.29 ;
      RECT  0.95 0.7 1.05 1.29 ;
      LAYER M2 ;
      RECT  0.91 1.15 2.09 1.25 ;
      LAYER V1 ;
      RECT  1.95 1.15 2.05 1.25 ;
      RECT  0.95 1.15 1.05 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.435 0.445 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  2.015 1.41 2.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.325 0.05 0.445 0.385 ;
      RECT  2.01 0.05 2.13 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.14 0.48 1.26 1.31 ;
      RECT  1.14 1.31 1.45 1.49 ;
    END
    ANTENNADIFFAREA 0.226 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.54 0.2 1.52 0.29 ;
      RECT  0.54 0.29 0.64 0.5 ;
      RECT  1.4 0.29 1.52 0.73 ;
      RECT  0.065 0.5 0.64 0.59 ;
      RECT  0.54 0.59 0.64 0.96 ;
      RECT  0.065 0.59 0.185 1.22 ;
      RECT  1.4 0.73 1.66 0.84 ;
      RECT  1.54 0.84 1.66 1.225 ;
      RECT  0.73 0.425 1.0 0.545 ;
      RECT  0.73 0.545 0.845 1.22 ;
      RECT  1.755 0.23 1.855 1.425 ;
      RECT  1.755 1.425 1.875 1.595 ;
  END
END SEN_EN2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_2
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_2
  CLASS CORE ;
  FOREIGN SEN_EN2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.97 0.87 3.585 0.96 ;
      RECT  3.35 0.96 3.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1824 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.175 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.575 1.41 0.695 1.75 ;
      RECT  1.035 1.625 1.205 1.75 ;
      RECT  3.44 1.41 3.56 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  1.035 0.05 1.205 0.175 ;
      RECT  0.055 0.05 0.175 0.39 ;
      RECT  0.575 0.05 0.695 0.39 ;
      RECT  3.365 0.05 3.485 0.58 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.14 0.2 2.805 0.315 ;
      RECT  2.14 0.315 2.26 0.405 ;
      RECT  1.595 0.405 2.26 0.445 ;
      RECT  1.15 0.445 2.26 0.535 ;
      RECT  1.15 0.535 1.25 1.24 ;
      RECT  1.15 1.24 2.26 1.355 ;
      RECT  1.595 1.355 2.26 1.36 ;
      RECT  2.14 1.36 2.26 1.48 ;
      RECT  2.14 1.48 2.805 1.6 ;
    END
    ANTENNADIFFAREA 0.408 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.335 0.205 2.025 0.265 ;
      RECT  0.875 0.265 2.025 0.315 ;
      RECT  0.875 0.315 1.45 0.355 ;
      RECT  0.875 0.355 0.995 0.51 ;
      RECT  0.76 0.51 0.995 0.68 ;
      RECT  0.875 0.68 0.995 1.035 ;
      RECT  0.76 1.035 0.995 1.205 ;
      RECT  0.875 1.205 0.995 1.445 ;
      RECT  0.875 1.445 1.505 1.485 ;
      RECT  0.875 1.485 2.025 1.535 ;
      RECT  1.335 1.535 2.025 1.6 ;
      RECT  2.92 0.16 3.03 0.405 ;
      RECT  2.375 0.405 3.03 0.52 ;
      RECT  2.375 0.52 2.465 0.68 ;
      RECT  1.34 0.68 2.465 0.77 ;
      RECT  1.34 0.77 1.43 1.04 ;
      RECT  1.34 1.04 2.485 1.13 ;
      RECT  2.375 1.13 2.485 1.24 ;
      RECT  2.375 1.24 3.04 1.36 ;
      RECT  2.92 1.36 3.04 1.61 ;
      RECT  0.315 0.37 0.435 0.5 ;
      RECT  0.315 0.5 0.64 0.59 ;
      RECT  0.55 0.59 0.64 0.775 ;
      RECT  0.55 0.775 0.785 0.945 ;
      RECT  0.55 0.945 0.64 1.01 ;
      RECT  0.34 1.01 0.64 1.1 ;
      RECT  0.34 1.1 0.43 1.21 ;
      RECT  0.31 1.21 0.43 1.43 ;
      RECT  3.12 0.49 3.225 0.625 ;
      RECT  2.675 0.625 3.225 0.67 ;
      RECT  2.675 0.67 3.745 0.725 ;
      RECT  3.625 0.49 3.745 0.67 ;
      RECT  3.12 0.725 3.745 0.76 ;
      RECT  2.675 0.725 2.78 0.86 ;
      RECT  1.63 0.86 2.78 0.95 ;
      RECT  2.675 0.95 2.78 1.055 ;
      RECT  2.675 1.055 3.25 1.145 ;
      RECT  3.14 1.145 3.25 1.33 ;
  END
END SEN_EN2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_3
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_3
  CLASS CORE ;
  FOREIGN SEN_EN2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.515 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.5 4.25 0.71 ;
      RECT  3.95 0.71 4.25 0.89 ;
      RECT  2.35 0.49 2.45 0.71 ;
      RECT  1.93 0.71 2.45 0.89 ;
      LAYER M2 ;
      RECT  2.31 0.55 4.295 0.65 ;
      LAYER V1 ;
      RECT  4.15 0.55 4.25 0.65 ;
      RECT  2.35 0.55 2.45 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2736 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.39 0.445 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.845 1.2 0.965 1.75 ;
      RECT  1.365 1.415 1.485 1.75 ;
      RECT  3.955 1.415 4.075 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  1.365 0.05 1.485 0.375 ;
      RECT  0.325 0.05 0.445 0.385 ;
      RECT  3.685 0.05 3.795 0.39 ;
      RECT  4.195 0.05 4.315 0.39 ;
      RECT  0.845 0.05 0.965 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.86 0.215 3.595 0.33 ;
      RECT  3.505 0.33 3.595 0.7 ;
      RECT  3.35 0.7 3.595 0.89 ;
      RECT  3.35 0.89 3.45 1.11 ;
      RECT  2.75 1.11 3.45 1.29 ;
      RECT  2.75 1.29 2.85 1.33 ;
      RECT  2.11 1.33 2.85 1.45 ;
    END
    ANTENNADIFFAREA 0.686 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.37 1.225 0.47 ;
      RECT  1.105 0.47 2.26 0.59 ;
      RECT  2.145 0.42 2.26 0.47 ;
      RECT  1.265 0.59 1.365 1.21 ;
      RECT  1.105 1.21 1.745 1.3 ;
      RECT  1.105 1.3 1.225 1.43 ;
      RECT  1.625 1.3 1.745 1.55 ;
      RECT  1.625 1.55 3.585 1.64 ;
      RECT  2.945 1.435 3.065 1.55 ;
      RECT  3.465 1.42 3.585 1.55 ;
      RECT  3.305 0.42 3.415 0.47 ;
      RECT  2.57 0.47 3.415 0.59 ;
      RECT  2.57 0.59 2.66 1.12 ;
      RECT  1.455 0.795 1.645 0.885 ;
      RECT  1.555 0.885 1.645 1.01 ;
      RECT  1.555 1.01 1.995 1.1 ;
      RECT  1.875 1.1 1.995 1.12 ;
      RECT  1.875 1.12 2.66 1.235 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.59 ;
      RECT  0.585 0.37 0.705 0.5 ;
      RECT  0.605 0.59 0.705 0.79 ;
      RECT  0.605 0.79 1.175 0.89 ;
      RECT  0.605 0.89 0.705 1.21 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.585 1.3 0.705 1.43 ;
      RECT  3.935 0.36 4.055 0.5 ;
      RECT  3.695 0.5 4.055 0.59 ;
      RECT  3.695 0.59 3.795 1.03 ;
      RECT  3.59 1.03 3.795 1.14 ;
      RECT  3.695 1.14 3.795 1.21 ;
      RECT  3.695 1.21 4.335 1.3 ;
      RECT  3.695 1.3 3.815 1.43 ;
      RECT  4.215 1.3 4.335 1.46 ;
  END
END SEN_EN2_3
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_4
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_4
  CLASS CORE ;
  FOREIGN SEN_EN2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.715 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.45 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
      RECT  2.95 0.8 3.14 1.09 ;
      LAYER M2 ;
      RECT  2.94 0.95 5.29 1.05 ;
      LAYER V1 ;
      RECT  5.15 0.95 5.25 1.05 ;
      RECT  2.995 0.95 3.095 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3645 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  1.105 1.2 1.225 1.75 ;
      RECT  1.625 1.2 1.745 1.75 ;
      RECT  2.12 1.465 2.29 1.75 ;
      RECT  4.815 1.41 4.935 1.75 ;
      RECT  5.335 1.41 5.455 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  0.585 0.05 0.705 0.385 ;
      RECT  5.075 0.05 5.195 0.385 ;
      RECT  5.6 0.05 5.72 0.39 ;
      RECT  1.625 0.05 1.745 0.42 ;
      RECT  2.145 0.05 2.265 0.42 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.105 0.05 1.225 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.2 4.65 0.31 ;
      RECT  2.41 0.31 2.53 0.42 ;
      RECT  4.49 0.31 4.65 0.6 ;
      RECT  3.95 0.6 4.65 0.69 ;
      RECT  3.95 0.69 4.05 1.11 ;
      RECT  3.505 1.11 4.665 1.3 ;
      RECT  3.505 1.3 3.625 1.36 ;
      RECT  2.32 1.08 2.65 1.18 ;
      RECT  2.56 1.18 2.65 1.36 ;
      RECT  2.56 1.36 3.625 1.46 ;
    END
    ANTENNADIFFAREA 0.931 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.815 0.32 4.935 0.495 ;
      RECT  4.815 0.495 5.46 0.585 ;
      RECT  5.34 0.32 5.46 0.495 ;
      RECT  4.815 0.585 4.935 0.815 ;
      RECT  4.15 0.815 4.935 0.925 ;
      RECT  4.815 0.925 4.935 1.21 ;
      RECT  4.815 1.21 5.195 1.31 ;
      RECT  5.075 1.31 5.195 1.43 ;
      RECT  0.325 0.37 0.445 0.5 ;
      RECT  0.325 0.5 0.965 0.59 ;
      RECT  0.845 0.59 0.965 0.79 ;
      RECT  0.845 0.79 1.635 0.89 ;
      RECT  0.845 0.89 0.965 1.21 ;
      RECT  0.325 1.21 0.965 1.3 ;
      RECT  0.325 1.3 0.445 1.43 ;
      RECT  3.71 0.4 4.375 0.505 ;
      RECT  3.71 0.505 3.83 0.77 ;
      RECT  3.245 0.77 3.83 0.88 ;
      RECT  3.245 0.88 3.365 1.18 ;
      RECT  1.94 0.79 2.845 0.885 ;
      RECT  2.74 0.885 2.845 1.18 ;
      RECT  2.74 1.18 3.365 1.27 ;
      RECT  1.365 0.46 1.485 0.56 ;
      RECT  1.365 0.56 3.36 0.68 ;
      RECT  1.735 0.68 1.835 1.01 ;
      RECT  1.36 1.01 2.005 1.1 ;
      RECT  1.36 1.1 1.49 1.23 ;
      RECT  1.885 1.1 2.005 1.27 ;
      RECT  1.885 1.27 2.47 1.36 ;
      RECT  2.38 1.36 2.47 1.55 ;
      RECT  2.38 1.55 4.405 1.64 ;
      RECT  3.765 1.435 3.885 1.55 ;
      RECT  4.285 1.435 4.405 1.55 ;
  END
END SEN_EN2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_5
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_5
  CLASS CORE ;
  FOREIGN SEN_EN2_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.955 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.71 6.05 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
      RECT  3.075 0.71 3.65 0.915 ;
      RECT  3.55 0.915 3.65 0.95 ;
      RECT  3.55 0.95 3.73 1.05 ;
      LAYER M2 ;
      RECT  3.55 0.95 5.69 1.05 ;
      LAYER V1 ;
      RECT  5.55 0.95 5.65 1.05 ;
      RECT  3.59 0.95 3.69 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4125 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.415 0.44 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.83 1.415 0.96 1.75 ;
      RECT  1.355 1.21 1.475 1.75 ;
      RECT  1.87 1.435 2.0 1.75 ;
      RECT  2.39 1.435 2.52 1.75 ;
      RECT  5.435 1.44 5.565 1.75 ;
      RECT  6.04 1.21 6.16 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  0.31 0.05 0.44 0.385 ;
      RECT  0.83 0.05 0.96 0.385 ;
      RECT  1.87 0.05 2.0 0.385 ;
      RECT  2.39 0.05 2.52 0.385 ;
      RECT  5.695 0.05 5.825 0.395 ;
      RECT  6.215 0.05 6.34 0.44 ;
      RECT  1.355 0.05 1.475 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.435 0.5 5.25 0.69 ;
      RECT  4.545 0.69 4.655 1.11 ;
      RECT  4.015 1.11 5.14 1.29 ;
      RECT  4.015 1.29 4.125 1.345 ;
      RECT  2.865 1.345 4.125 1.46 ;
      RECT  2.865 0.46 4.1 0.58 ;
      RECT  3.75 0.58 4.1 0.69 ;
      LAYER M2 ;
      RECT  3.71 0.55 4.58 0.65 ;
      LAYER V1 ;
      RECT  4.44 0.55 4.54 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  3.95 0.55 4.05 0.65 ;
    END
    ANTENNADIFFAREA 0.978 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.23 0.215 5.425 0.335 ;
      RECT  4.23 0.335 4.34 0.91 ;
      RECT  3.82 0.91 4.34 1.02 ;
      RECT  3.82 1.02 3.925 1.14 ;
      RECT  2.2 0.785 2.985 0.895 ;
      RECT  2.875 0.895 2.985 1.14 ;
      RECT  2.875 1.14 3.925 1.255 ;
      RECT  0.055 0.19 0.175 0.485 ;
      RECT  0.055 0.485 1.215 0.605 ;
      RECT  1.095 0.605 1.215 0.785 ;
      RECT  1.095 0.785 1.93 0.895 ;
      RECT  1.095 0.895 1.215 1.195 ;
      RECT  0.055 1.195 1.215 1.315 ;
      RECT  0.055 1.315 0.175 1.61 ;
      RECT  5.355 0.485 6.13 0.6 ;
      RECT  5.355 0.6 5.45 0.81 ;
      RECT  4.745 0.81 5.45 0.92 ;
      RECT  5.35 0.92 5.45 1.23 ;
      RECT  5.35 1.23 5.88 1.35 ;
      RECT  4.215 1.415 4.905 1.535 ;
      RECT  4.215 1.535 4.335 1.55 ;
      RECT  2.655 0.24 3.865 0.36 ;
      RECT  2.655 0.36 2.775 0.485 ;
      RECT  1.565 0.485 2.775 0.605 ;
      RECT  2.02 0.605 2.11 1.225 ;
      RECT  1.565 1.225 2.775 1.345 ;
      RECT  2.655 1.345 2.775 1.55 ;
      RECT  2.655 1.55 4.335 1.66 ;
      LAYER M2 ;
      RECT  1.065 0.95 3.02 1.05 ;
      LAYER V1 ;
      RECT  1.105 0.95 1.205 1.05 ;
      RECT  2.88 0.95 2.98 1.05 ;
  END
END SEN_EN2_5
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_6
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_6
  CLASS CORE ;
  FOREIGN SEN_EN2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.25 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.65 0.905 ;
      RECT  7.15 0.905 7.25 1.09 ;
      RECT  3.84 0.71 4.45 0.925 ;
      RECT  4.35 0.925 4.45 0.95 ;
      RECT  4.35 0.95 4.63 1.05 ;
      LAYER M2 ;
      RECT  4.45 0.95 7.29 1.05 ;
      LAYER V1 ;
      RECT  7.15 0.95 7.25 1.05 ;
      RECT  4.49 0.95 4.59 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5004 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.59 1.255 0.71 1.75 ;
      RECT  1.11 1.255 1.23 1.75 ;
      RECT  1.63 1.21 1.75 1.75 ;
      RECT  2.15 1.255 2.27 1.75 ;
      RECT  2.67 1.255 2.79 1.75 ;
      RECT  3.19 1.255 3.31 1.75 ;
      RECT  7.025 1.45 7.155 1.75 ;
      RECT  7.57 1.21 7.69 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  0.585 0.05 0.715 0.345 ;
      RECT  1.105 0.05 1.235 0.345 ;
      RECT  7.285 0.05 7.415 0.355 ;
      RECT  6.77 0.05 6.895 0.36 ;
      RECT  2.145 0.05 2.275 0.365 ;
      RECT  2.665 0.05 2.795 0.365 ;
      RECT  3.185 0.05 3.305 0.365 ;
      RECT  1.63 0.05 1.75 0.585 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.395 0.22 6.68 0.35 ;
      RECT  6.55 0.35 6.68 0.65 ;
      RECT  5.52 0.65 6.68 0.74 ;
      RECT  5.52 0.74 5.65 1.11 ;
      RECT  4.95 1.11 6.25 1.29 ;
      RECT  4.95 1.29 5.05 1.35 ;
      RECT  3.885 1.35 5.05 1.46 ;
    END
    ANTENNADIFFAREA 1.141 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.96 0.44 6.455 0.56 ;
      RECT  4.96 0.56 5.08 0.675 ;
      RECT  4.72 0.675 5.08 0.795 ;
      RECT  4.72 0.795 4.84 1.14 ;
      RECT  3.62 0.91 3.72 1.14 ;
      RECT  3.62 1.14 4.84 1.26 ;
      RECT  0.285 0.435 1.515 0.565 ;
      RECT  1.385 0.565 1.515 0.77 ;
      RECT  1.385 0.77 2.845 0.9 ;
      RECT  1.385 0.9 1.515 1.035 ;
      RECT  0.34 1.035 1.515 1.165 ;
      RECT  0.34 1.165 0.45 1.26 ;
      RECT  6.785 0.45 7.72 0.57 ;
      RECT  6.785 0.57 6.875 0.83 ;
      RECT  5.74 0.83 6.875 0.94 ;
      RECT  6.77 0.94 6.875 1.24 ;
      RECT  6.77 1.24 7.46 1.36 ;
      RECT  1.84 0.455 4.865 0.585 ;
      RECT  3.4 0.585 3.53 1.035 ;
      RECT  1.84 1.035 3.53 1.165 ;
      RECT  3.4 1.165 3.53 1.55 ;
      RECT  3.4 1.55 6.45 1.56 ;
      RECT  5.2 1.44 6.45 1.55 ;
      RECT  3.4 1.56 5.31 1.66 ;
      LAYER M2 ;
      RECT  1.375 0.55 5.11 0.65 ;
      RECT  1.375 0.95 3.76 1.05 ;
      LAYER V1 ;
      RECT  1.415 0.55 1.515 0.65 ;
      RECT  4.97 0.55 5.07 0.65 ;
      RECT  1.415 0.95 1.515 1.05 ;
      RECT  3.62 0.95 3.72 1.05 ;
  END
END SEN_EN2_6
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_8
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_8
  CLASS CORE ;
  FOREIGN SEN_EN2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.95 0.71 9.25 0.89 ;
      RECT  8.95 0.89 9.05 1.09 ;
      RECT  4.88 0.855 5.89 0.95 ;
      RECT  4.88 0.95 5.975 0.955 ;
      RECT  5.79 0.955 5.975 1.05 ;
      LAYER M2 ;
      RECT  5.795 0.95 9.09 1.05 ;
      LAYER V1 ;
      RECT  8.95 0.95 9.05 1.05 ;
      RECT  5.835 0.95 5.935 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.666 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.215 0.19 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.59 1.255 0.71 1.75 ;
      RECT  1.11 1.255 1.23 1.75 ;
      RECT  1.63 1.255 1.75 1.75 ;
      RECT  2.15 1.215 2.27 1.75 ;
      RECT  2.67 1.255 2.79 1.75 ;
      RECT  3.19 1.255 3.31 1.75 ;
      RECT  3.71 1.255 3.83 1.75 ;
      RECT  4.26 1.56 4.43 1.75 ;
      RECT  8.38 1.215 8.495 1.75 ;
      RECT  8.895 1.45 9.015 1.75 ;
      RECT  9.415 1.215 9.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  0.59 0.05 0.71 0.345 ;
      RECT  1.11 0.05 1.23 0.345 ;
      RECT  1.63 0.05 1.75 0.345 ;
      RECT  8.38 0.05 8.495 0.36 ;
      RECT  8.895 0.05 9.015 0.36 ;
      RECT  2.67 0.05 2.79 0.365 ;
      RECT  3.19 0.05 3.31 0.365 ;
      RECT  3.71 0.05 3.83 0.365 ;
      RECT  4.23 0.05 4.35 0.56 ;
      RECT  9.415 0.05 9.535 0.56 ;
      RECT  0.07 0.05 0.19 0.585 ;
      RECT  2.15 0.05 2.27 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.82 0.51 8.09 0.69 ;
      RECT  6.92 0.69 7.09 1.11 ;
      RECT  4.75 0.51 6.475 0.69 ;
      RECT  6.31 0.69 6.475 1.11 ;
      RECT  6.31 1.11 8.09 1.29 ;
      RECT  6.31 1.29 6.44 1.34 ;
      RECT  4.74 1.34 6.44 1.46 ;
    END
    ANTENNADIFFAREA 1.466 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.585 0.24 8.29 0.36 ;
      RECT  6.585 0.36 6.7 0.505 ;
      RECT  4.48 0.235 6.21 0.365 ;
      RECT  4.48 0.365 4.64 0.67 ;
      RECT  2.385 0.455 4.115 0.585 ;
      RECT  3.94 0.585 4.115 0.67 ;
      RECT  3.94 0.67 4.64 0.82 ;
      RECT  3.94 0.82 4.115 1.035 ;
      RECT  2.385 1.035 4.115 1.165 ;
      RECT  3.99 1.165 4.115 1.34 ;
      RECT  3.99 1.34 4.635 1.45 ;
      RECT  4.525 1.45 4.635 1.55 ;
      RECT  4.525 1.55 8.29 1.56 ;
      RECT  6.545 1.44 8.29 1.55 ;
      RECT  4.525 1.56 6.655 1.66 ;
      RECT  1.88 0.31 2.05 0.435 ;
      RECT  0.305 0.435 2.05 0.565 ;
      RECT  1.88 0.565 2.05 0.75 ;
      RECT  1.88 0.75 3.715 0.92 ;
      RECT  1.88 0.92 2.05 1.035 ;
      RECT  0.34 1.035 2.05 1.165 ;
      RECT  0.34 1.165 0.45 1.285 ;
      RECT  8.635 0.45 9.3 0.57 ;
      RECT  8.635 0.57 8.755 0.86 ;
      RECT  7.18 0.86 8.755 0.97 ;
      RECT  8.635 0.97 8.755 1.24 ;
      RECT  8.635 1.24 9.3 1.36 ;
      RECT  4.505 0.91 4.625 1.14 ;
      RECT  4.505 1.14 6.21 1.25 ;
      LAYER M2 ;
      RECT  1.91 0.35 6.725 0.45 ;
      RECT  1.91 0.95 4.65 1.05 ;
      LAYER V1 ;
      RECT  1.95 0.35 2.05 0.45 ;
      RECT  6.585 0.35 6.685 0.45 ;
      RECT  1.95 0.95 2.05 1.05 ;
      RECT  4.51 0.95 4.61 1.05 ;
  END
END SEN_EN2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_DG_1
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_DG_1
  CLASS CORE ;
  FOREIGN SEN_EN2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.625 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.445 1.45 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.735 1.44 1.865 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.32 0.05 0.45 0.345 ;
      RECT  1.74 0.05 1.86 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.445 2.155 0.555 ;
      RECT  1.95 0.555 2.05 1.045 ;
      RECT  1.95 1.045 2.155 1.155 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.755 0.16 1.645 0.33 ;
      RECT  1.545 0.33 1.645 1.05 ;
      RECT  1.345 1.05 1.645 1.16 ;
      RECT  0.065 0.2 0.185 0.435 ;
      RECT  0.065 0.435 0.505 0.535 ;
      RECT  0.4 0.535 0.505 1.235 ;
      RECT  0.07 1.235 0.505 1.325 ;
      RECT  0.07 1.325 0.18 1.58 ;
      RECT  1.75 0.73 1.85 1.25 ;
      RECT  1.455 1.25 1.85 1.35 ;
      RECT  1.455 1.35 1.555 1.45 ;
      RECT  0.855 0.42 0.975 1.45 ;
      RECT  0.855 1.45 1.555 1.55 ;
      RECT  1.12 0.42 1.235 1.335 ;
      RECT  0.595 0.41 0.71 1.58 ;
      LAYER M2 ;
      RECT  0.36 1.15 1.26 1.25 ;
      LAYER V1 ;
      RECT  0.4 1.15 0.5 1.25 ;
      RECT  1.12 1.15 1.22 1.25 ;
  END
END SEN_EN2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_DG_16
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_DG_16
  CLASS CORE ;
  FOREIGN SEN_EN2_DG_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.72 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.87 0.71 4.65 0.89 ;
      RECT  4.55 0.89 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.105 1.21 1.225 1.75 ;
      RECT  1.62 1.44 1.75 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  4.71 1.48 4.88 1.75 ;
      RECT  5.23 1.48 5.4 1.75 ;
      RECT  5.77 1.41 5.9 1.75 ;
      RECT  6.29 1.41 6.42 1.75 ;
      RECT  6.81 1.41 6.94 1.75 ;
      RECT  7.33 1.41 7.46 1.75 ;
      RECT  7.85 1.41 7.98 1.75 ;
      RECT  8.37 1.41 8.5 1.75 ;
      RECT  8.89 1.41 9.02 1.75 ;
      RECT  9.415 1.21 9.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  0.58 0.05 0.71 0.35 ;
      RECT  5.77 0.05 5.9 0.35 ;
      RECT  6.29 0.05 6.42 0.35 ;
      RECT  6.81 0.05 6.94 0.35 ;
      RECT  7.33 0.05 7.46 0.35 ;
      RECT  7.85 0.05 7.98 0.35 ;
      RECT  8.37 0.05 8.5 0.35 ;
      RECT  8.89 0.05 9.02 0.35 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.14 0.05 2.265 0.36 ;
      RECT  4.73 0.05 4.86 0.37 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.105 0.05 1.225 0.59 ;
      RECT  5.255 0.05 5.375 0.59 ;
      RECT  9.415 0.05 9.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.345 0.44 8.845 0.49 ;
      RECT  5.515 0.49 8.845 0.51 ;
      RECT  5.515 0.51 9.275 0.69 ;
      RECT  8.53 0.69 8.85 1.04 ;
      RECT  7.615 1.04 8.85 1.11 ;
      RECT  5.515 1.11 9.275 1.29 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 0.44 0.99 0.56 ;
      RECT  0.89 0.56 0.99 0.785 ;
      RECT  0.89 0.785 1.975 0.895 ;
      RECT  0.89 0.895 0.99 1.24 ;
      RECT  0.275 1.24 0.99 1.35 ;
      RECT  1.315 0.45 3.33 0.56 ;
      RECT  2.335 0.56 2.425 1.24 ;
      RECT  1.315 1.24 4.395 1.35 ;
      RECT  3.61 0.44 4.395 0.56 ;
      RECT  3.61 0.56 3.71 1.04 ;
      RECT  2.64 0.91 2.74 1.04 ;
      RECT  2.64 1.04 3.71 1.15 ;
      RECT  3.42 0.51 3.52 0.785 ;
      RECT  2.88 0.785 3.52 0.895 ;
      RECT  5.255 0.8 8.385 0.91 ;
      RECT  5.255 0.91 7.51 0.97 ;
      RECT  5.255 0.97 5.425 1.22 ;
      RECT  2.355 0.24 4.605 0.35 ;
      RECT  4.485 0.35 4.605 0.48 ;
      RECT  4.485 0.48 4.88 0.595 ;
      RECT  4.76 0.595 4.88 1.22 ;
      RECT  4.76 1.22 5.425 1.27 ;
      RECT  4.485 1.27 5.425 1.39 ;
      RECT  4.485 1.39 4.605 1.44 ;
      RECT  2.38 1.44 4.605 1.56 ;
      RECT  4.97 0.415 5.115 1.03 ;
      RECT  4.97 1.03 5.14 1.12 ;
      LAYER M2 ;
      RECT  3.38 0.55 5.14 0.65 ;
      RECT  0.85 0.95 2.78 1.05 ;
      LAYER V1 ;
      RECT  3.42 0.55 3.52 0.65 ;
      RECT  5.0 0.55 5.1 0.65 ;
      RECT  0.89 0.95 0.99 1.05 ;
      RECT  2.64 0.95 2.74 1.05 ;
  END
END SEN_EN2_DG_16
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_DG_2
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_DG_2
  CLASS CORE ;
  FOREIGN SEN_EN2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.64 0.25 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.535 0.46 1.65 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.435 0.45 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.66 1.44 1.79 1.75 ;
      RECT  2.215 1.21 2.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  1.67 0.05 1.8 0.37 ;
      RECT  2.215 0.05 2.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.415 2.075 0.645 ;
      RECT  1.95 0.645 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.234 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.765 0.19 1.485 0.36 ;
      RECT  1.355 0.36 1.445 1.05 ;
      RECT  1.355 1.05 1.57 1.16 ;
      RECT  0.07 0.22 0.18 0.45 ;
      RECT  0.07 0.45 0.51 0.55 ;
      RECT  0.41 0.55 0.51 1.245 ;
      RECT  0.065 1.245 0.51 1.345 ;
      RECT  0.065 1.345 0.185 1.51 ;
      RECT  1.765 0.725 1.86 1.25 ;
      RECT  1.46 1.25 1.86 1.35 ;
      RECT  1.46 1.35 1.57 1.41 ;
      RECT  0.855 0.45 0.975 1.41 ;
      RECT  0.855 1.41 1.57 1.53 ;
      RECT  1.12 0.45 1.22 1.29 ;
      RECT  0.6 0.45 0.71 1.52 ;
      LAYER M2 ;
      RECT  0.37 1.15 1.26 1.25 ;
      LAYER V1 ;
      RECT  0.41 1.15 0.51 1.25 ;
      RECT  1.12 1.15 1.22 1.25 ;
  END
END SEN_EN2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_DG_4
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_DG_4
  CLASS CORE ;
  FOREIGN SEN_EN2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.65 0.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.645 1.28 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.45 0.45 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.855 1.465 2.025 1.75 ;
      RECT  2.395 1.41 2.525 1.75 ;
      RECT  2.96 1.21 3.08 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.32 0.05 0.45 0.345 ;
      RECT  2.425 0.05 2.555 0.39 ;
      RECT  1.88 0.05 2.0 0.59 ;
      RECT  2.96 0.05 3.08 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.85 0.69 ;
      RECT  2.75 0.69 2.85 1.11 ;
      RECT  2.14 1.11 2.85 1.29 ;
    END
    ANTENNADIFFAREA 0.474 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.34 0.185 0.44 ;
      RECT  0.065 0.44 0.51 0.56 ;
      RECT  0.41 0.56 0.51 1.24 ;
      RECT  0.065 1.24 0.51 1.36 ;
      RECT  0.065 1.36 0.185 1.48 ;
      RECT  0.97 0.445 1.24 0.555 ;
      RECT  0.97 0.555 1.06 1.06 ;
      RECT  0.835 1.06 1.06 1.15 ;
      RECT  0.835 1.15 0.955 1.29 ;
      RECT  1.96 0.79 2.64 0.89 ;
      RECT  1.96 0.89 2.05 1.255 ;
      RECT  0.795 0.23 1.475 0.34 ;
      RECT  1.37 0.34 1.475 1.255 ;
      RECT  1.05 1.255 2.05 1.365 ;
      RECT  0.78 0.45 0.88 0.97 ;
      RECT  1.605 0.21 1.725 1.16 ;
      RECT  0.6 0.445 0.69 1.46 ;
      RECT  0.6 1.46 1.525 1.57 ;
      LAYER M2 ;
      RECT  0.74 0.55 1.765 0.65 ;
      RECT  0.37 1.15 0.995 1.25 ;
      LAYER V1 ;
      RECT  0.78 0.55 0.88 0.65 ;
      RECT  1.625 0.55 1.725 0.65 ;
      RECT  0.41 1.15 0.51 1.25 ;
      RECT  0.855 1.15 0.955 1.25 ;
  END
END SEN_EN2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_DG_8
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_DG_8
  CLASS CORE ;
  FOREIGN SEN_EN2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.645 0.45 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.91 ;
      RECT  2.15 0.91 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  2.93 1.44 3.06 1.75 ;
      RECT  3.45 1.41 3.58 1.75 ;
      RECT  3.97 1.41 4.1 1.75 ;
      RECT  4.49 1.41 4.62 1.75 ;
      RECT  5.015 1.21 5.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.91 0.05 3.08 0.305 ;
      RECT  0.58 0.05 0.71 0.355 ;
      RECT  1.115 0.05 1.24 0.36 ;
      RECT  3.45 0.05 3.58 0.39 ;
      RECT  3.97 0.05 4.1 0.39 ;
      RECT  4.49 0.05 4.62 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.015 0.05 5.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 4.88 0.69 ;
      RECT  4.28 0.69 4.45 1.11 ;
      RECT  3.15 1.11 4.865 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.345 0.245 2.82 0.355 ;
      RECT  2.73 0.355 2.82 0.395 ;
      RECT  2.73 0.395 3.05 0.485 ;
      RECT  2.95 0.485 3.05 0.785 ;
      RECT  2.95 0.785 4.19 0.895 ;
      RECT  2.95 0.895 3.05 1.25 ;
      RECT  2.505 1.25 3.05 1.35 ;
      RECT  2.505 1.35 2.6 1.445 ;
      RECT  1.32 1.445 2.6 1.555 ;
      RECT  0.275 0.445 0.73 0.555 ;
      RECT  0.63 0.555 0.73 0.785 ;
      RECT  0.63 0.785 0.98 0.895 ;
      RECT  0.63 0.895 0.73 1.24 ;
      RECT  0.275 1.24 0.73 1.35 ;
      RECT  0.82 0.45 1.8 0.555 ;
      RECT  1.3 0.555 1.8 0.565 ;
      RECT  1.3 0.565 1.39 1.245 ;
      RECT  0.82 1.245 2.325 1.35 ;
      RECT  1.96 0.445 2.26 0.555 ;
      RECT  2.15 0.555 2.26 0.615 ;
      RECT  1.96 0.555 2.06 1.045 ;
      RECT  1.52 1.045 2.06 1.155 ;
      RECT  2.625 0.575 2.82 0.68 ;
      RECT  2.72 0.68 2.82 1.015 ;
      RECT  2.625 1.015 2.82 1.135 ;
      RECT  1.53 0.69 1.87 0.91 ;
      LAYER M2 ;
      RECT  0.59 0.55 2.13 0.65 ;
      RECT  1.47 0.75 2.86 0.85 ;
      LAYER V1 ;
      RECT  0.63 0.55 0.73 0.65 ;
      RECT  1.96 0.55 2.06 0.65 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  2.72 0.75 2.82 0.85 ;
  END
END SEN_EN2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_S_0P5
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_S_0P5
  CLASS CORE ;
  FOREIGN SEN_EN2_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.71 0.45 0.935 ;
      RECT  0.35 0.935 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 1.11 0.65 1.57 ;
      RECT  0.55 1.57 1.85 1.66 ;
      RECT  1.75 1.31 1.85 1.57 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0492 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.34 0.46 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  2.01 0.99 2.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.33 0.05 0.455 0.38 ;
      RECT  2.01 0.05 2.14 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.32 1.165 0.44 ;
      RECT  0.95 0.44 1.05 0.91 ;
      RECT  0.95 0.91 1.385 1.09 ;
      RECT  1.265 1.09 1.385 1.46 ;
    END
    ANTENNADIFFAREA 0.1 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.545 0.14 1.385 0.23 ;
      RECT  0.545 0.23 0.635 0.5 ;
      RECT  1.265 0.23 1.385 0.65 ;
      RECT  0.065 0.24 0.185 0.5 ;
      RECT  0.065 0.5 0.635 0.59 ;
      RECT  0.545 0.59 0.635 0.925 ;
      RECT  0.065 0.59 0.17 1.55 ;
      RECT  1.265 0.65 1.645 0.74 ;
      RECT  1.525 0.74 1.645 1.46 ;
      RECT  1.495 0.215 1.875 0.325 ;
      RECT  1.755 0.325 1.875 1.19 ;
      RECT  0.74 0.32 0.845 1.355 ;
      RECT  0.74 1.355 1.175 1.475 ;
  END
END SEN_EN2_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_S_1
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_S_1
  CLASS CORE ;
  FOREIGN SEN_EN2_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.71 0.45 0.925 ;
      RECT  0.35 0.925 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0633 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 1.11 0.65 1.53 ;
      RECT  0.55 1.53 1.85 1.62 ;
      RECT  1.75 1.31 1.85 1.53 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0927 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.39 0.46 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  2.01 1.02 2.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.33 0.05 0.455 0.39 ;
      RECT  2.01 0.05 2.14 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.44 1.165 0.56 ;
      RECT  0.95 0.56 1.05 0.91 ;
      RECT  0.95 0.91 1.385 1.09 ;
      RECT  1.265 1.09 1.385 1.29 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.545 0.18 1.385 0.27 ;
      RECT  0.545 0.27 0.635 0.5 ;
      RECT  1.265 0.27 1.385 0.65 ;
      RECT  0.065 0.5 0.635 0.59 ;
      RECT  0.545 0.59 0.635 0.925 ;
      RECT  0.065 0.59 0.17 1.3 ;
      RECT  1.265 0.65 1.645 0.74 ;
      RECT  1.525 0.74 1.645 1.34 ;
      RECT  1.495 0.255 1.875 0.345 ;
      RECT  1.755 0.345 1.875 1.19 ;
      RECT  0.74 0.415 0.845 1.255 ;
      RECT  0.74 1.255 1.15 1.375 ;
  END
END SEN_EN2_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_S_2
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_S_2
  CLASS CORE ;
  FOREIGN SEN_EN2_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1266 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 1.09 ;
      RECT  1.95 0.51 2.05 0.64 ;
      RECT  1.55 0.64 2.05 0.73 ;
      RECT  1.55 0.73 1.65 0.95 ;
      LAYER M2 ;
      RECT  1.91 0.55 3.29 0.65 ;
      LAYER V1 ;
      RECT  3.15 0.55 3.25 0.65 ;
      RECT  1.95 0.55 2.05 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1851 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.6 1.21 0.72 1.75 ;
      RECT  1.125 1.44 1.255 1.75 ;
      RECT  3.19 1.21 3.31 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  1.125 0.05 1.245 0.36 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  2.645 0.05 2.775 0.39 ;
      RECT  3.185 0.05 3.315 0.39 ;
      RECT  0.595 0.05 0.715 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.335 0.2 2.545 0.32 ;
      RECT  2.35 0.32 2.45 1.11 ;
      RECT  2.13 1.11 2.775 1.29 ;
      RECT  2.13 1.29 2.25 1.325 ;
      RECT  1.565 1.325 2.25 1.445 ;
    END
    ANTENNADIFFAREA 0.497 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.335 0.41 1.79 0.475 ;
      RECT  0.885 0.475 1.79 0.53 ;
      RECT  0.885 0.53 1.425 0.565 ;
      RECT  0.885 0.565 0.99 1.26 ;
      RECT  0.885 1.26 1.445 1.35 ;
      RECT  1.355 1.35 1.445 1.555 ;
      RECT  1.355 1.555 2.51 1.645 ;
      RECT  2.39 1.38 2.51 1.555 ;
      RECT  0.34 0.445 0.445 0.755 ;
      RECT  0.34 0.755 0.795 0.845 ;
      RECT  0.695 0.845 0.795 1.11 ;
      RECT  0.34 0.845 0.445 1.255 ;
      RECT  2.155 0.46 2.245 0.845 ;
      RECT  1.935 0.845 2.245 0.935 ;
      RECT  1.935 0.935 2.025 1.055 ;
      RECT  1.115 0.91 1.215 1.055 ;
      RECT  1.115 1.055 2.025 1.17 ;
      RECT  2.91 0.29 3.03 0.85 ;
      RECT  2.54 0.85 3.03 0.94 ;
      RECT  2.91 0.94 3.03 1.395 ;
      LAYER M2 ;
      RECT  0.62 0.95 1.29 1.05 ;
      LAYER V1 ;
      RECT  0.695 0.95 0.795 1.05 ;
      RECT  1.115 0.95 1.215 1.05 ;
  END
END SEN_EN2_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_S_3
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_S_3
  CLASS CORE ;
  FOREIGN SEN_EN2_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.495 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1899 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.51 4.25 1.09 ;
      RECT  2.45 0.51 2.55 0.71 ;
      RECT  1.95 0.71 2.55 0.8 ;
      RECT  1.95 0.8 2.385 0.94 ;
      LAYER M2 ;
      RECT  2.41 0.55 4.29 0.65 ;
      LAYER V1 ;
      RECT  4.15 0.55 4.25 0.65 ;
      RECT  2.45 0.55 2.55 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2778 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.435 0.45 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.845 1.21 0.965 1.75 ;
      RECT  1.36 1.435 1.49 1.75 ;
      RECT  3.695 1.21 3.815 1.75 ;
      RECT  4.215 1.21 4.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  1.36 0.05 1.49 0.365 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  4.21 0.05 4.34 0.39 ;
      RECT  0.845 0.05 0.965 0.59 ;
      RECT  3.695 0.05 3.815 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.83 0.215 3.555 0.32 ;
      RECT  3.435 0.32 3.555 0.635 ;
      RECT  2.95 0.635 3.555 0.725 ;
      RECT  2.95 0.725 3.05 1.11 ;
      RECT  2.67 1.11 3.45 1.29 ;
      RECT  2.67 1.29 2.8 1.335 ;
      RECT  2.11 1.335 2.8 1.455 ;
    END
    ANTENNADIFFAREA 0.646 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.315 0.185 0.47 ;
      RECT  0.065 0.47 0.705 0.56 ;
      RECT  0.585 0.56 0.705 0.785 ;
      RECT  0.585 0.785 1.51 0.895 ;
      RECT  0.585 0.895 0.7 1.255 ;
      RECT  0.065 1.255 0.7 1.345 ;
      RECT  0.065 1.345 0.185 1.485 ;
      RECT  2.65 0.425 3.34 0.545 ;
      RECT  2.65 0.545 2.775 0.89 ;
      RECT  2.49 0.89 2.775 0.98 ;
      RECT  2.49 0.98 2.58 1.11 ;
      RECT  1.87 1.11 2.58 1.22 ;
      RECT  1.87 1.22 1.995 1.365 ;
      RECT  3.955 0.445 4.06 0.815 ;
      RECT  3.14 0.815 4.06 0.925 ;
      RECT  3.955 0.925 4.06 1.485 ;
      RECT  2.89 1.425 3.605 1.545 ;
      RECT  2.89 1.545 2.98 1.57 ;
      RECT  1.055 0.455 2.315 0.575 ;
      RECT  1.625 0.575 1.745 1.225 ;
      RECT  1.055 1.225 1.745 1.345 ;
      RECT  1.625 1.345 1.745 1.57 ;
      RECT  1.625 1.57 2.98 1.66 ;
      LAYER M2 ;
      RECT  0.56 1.15 2.02 1.25 ;
      LAYER V1 ;
      RECT  0.6 1.15 0.7 1.25 ;
      RECT  1.88 1.15 1.98 1.25 ;
  END
END SEN_EN2_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_S_4
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_S_4
  CLASS CORE ;
  FOREIGN SEN_EN2_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.775 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2532 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.45 0.89 ;
      RECT  5.35 0.89 5.45 1.09 ;
      RECT  2.55 0.71 3.05 0.94 ;
      RECT  2.95 0.94 3.05 1.09 ;
      LAYER M2 ;
      RECT  2.91 0.95 5.49 1.05 ;
      LAYER V1 ;
      RECT  5.35 0.95 5.45 1.05 ;
      RECT  2.95 0.95 3.05 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3708 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.59 1.25 0.71 1.75 ;
      RECT  1.11 1.21 1.23 1.75 ;
      RECT  1.63 1.25 1.75 1.75 ;
      RECT  2.15 1.21 2.265 1.75 ;
      RECT  4.81 1.21 4.93 1.75 ;
      RECT  5.35 1.21 5.47 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.585 0.05 0.715 0.35 ;
      RECT  4.9 0.05 5.03 0.35 ;
      RECT  1.625 0.05 1.755 0.36 ;
      RECT  2.145 0.05 2.265 0.36 ;
      RECT  5.42 0.05 5.545 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  1.11 0.05 1.23 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.46 0.17 4.565 0.24 ;
      RECT  2.355 0.24 4.565 0.35 ;
      RECT  4.46 0.35 4.565 0.65 ;
      RECT  3.95 0.65 4.565 0.74 ;
      RECT  3.95 0.74 4.05 1.11 ;
      RECT  3.535 1.11 4.68 1.245 ;
      RECT  4.55 1.245 4.68 1.335 ;
      RECT  3.535 1.245 3.65 1.445 ;
      RECT  2.355 1.445 3.65 1.56 ;
    END
    ANTENNADIFFAREA 0.91 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.285 0.44 1.0 0.56 ;
      RECT  0.91 0.56 1.0 0.8 ;
      RECT  0.91 0.8 1.8 0.89 ;
      RECT  0.91 0.89 1.01 1.04 ;
      RECT  0.34 1.04 1.01 1.16 ;
      RECT  0.34 1.16 0.45 1.285 ;
      RECT  3.645 0.44 4.365 0.56 ;
      RECT  3.645 0.56 3.735 0.855 ;
      RECT  3.355 0.855 3.735 0.945 ;
      RECT  3.355 0.945 3.445 1.24 ;
      RECT  2.36 0.91 2.46 1.24 ;
      RECT  2.36 1.24 3.445 1.355 ;
      RECT  4.655 0.44 5.34 0.56 ;
      RECT  4.655 0.56 4.765 0.85 ;
      RECT  4.15 0.85 4.86 0.94 ;
      RECT  4.77 0.94 4.86 0.98 ;
      RECT  4.77 0.98 5.19 1.07 ;
      RECT  5.07 1.07 5.19 1.35 ;
      RECT  1.32 0.45 3.335 0.57 ;
      RECT  1.89 0.57 2.01 1.055 ;
      RECT  1.345 1.055 2.01 1.16 ;
      RECT  1.89 1.16 2.01 1.49 ;
      RECT  3.75 1.34 4.46 1.46 ;
      LAYER M2 ;
      RECT  0.87 0.95 2.5 1.05 ;
      RECT  1.855 1.35 3.93 1.45 ;
      LAYER V1 ;
      RECT  0.91 0.95 1.01 1.05 ;
      RECT  2.36 0.95 2.46 1.05 ;
      RECT  1.895 1.35 1.995 1.45 ;
      RECT  3.79 1.35 3.89 1.45 ;
  END
END SEN_EN2_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_S_6
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_S_6
  CLASS CORE ;
  FOREIGN SEN_EN2_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.25 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3798 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.65 0.91 ;
      RECT  7.15 0.91 7.25 1.09 ;
      RECT  3.84 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 0.95 ;
      RECT  4.35 0.95 4.63 1.05 ;
      LAYER M2 ;
      RECT  4.45 0.95 7.29 1.05 ;
      LAYER V1 ;
      RECT  7.15 0.95 7.25 1.05 ;
      RECT  4.49 0.95 4.59 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5553 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 8.0 1.85 ;
      RECT  0.59 1.255 0.71 1.75 ;
      RECT  1.11 1.255 1.23 1.75 ;
      RECT  1.63 1.21 1.75 1.75 ;
      RECT  2.15 1.255 2.27 1.75 ;
      RECT  2.67 1.255 2.79 1.75 ;
      RECT  3.19 1.255 3.31 1.75 ;
      RECT  7.025 1.45 7.155 1.75 ;
      RECT  7.64 1.21 7.76 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      RECT  0.585 0.05 0.715 0.345 ;
      RECT  1.105 0.05 1.235 0.345 ;
      RECT  7.285 0.05 7.415 0.355 ;
      RECT  6.77 0.05 6.895 0.36 ;
      RECT  2.145 0.05 2.275 0.365 ;
      RECT  2.665 0.05 2.795 0.365 ;
      RECT  3.185 0.05 3.305 0.365 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  1.63 0.05 1.75 0.59 ;
      RECT  7.81 0.05 7.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.395 0.21 6.68 0.34 ;
      RECT  6.55 0.34 6.68 0.62 ;
      RECT  5.35 0.62 6.68 0.75 ;
      RECT  5.35 0.75 5.48 1.11 ;
      RECT  4.95 1.11 6.25 1.29 ;
      RECT  4.95 1.29 5.05 1.345 ;
      RECT  3.89 1.345 5.05 1.46 ;
    END
    ANTENNADIFFAREA 1.221 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.96 0.43 6.425 0.53 ;
      RECT  4.96 0.53 5.08 0.675 ;
      RECT  4.72 0.675 5.08 0.795 ;
      RECT  4.72 0.795 4.84 1.14 ;
      RECT  3.62 0.91 3.72 1.14 ;
      RECT  3.62 1.14 4.84 1.255 ;
      RECT  6.785 0.45 7.715 0.56 ;
      RECT  6.785 0.56 6.875 0.84 ;
      RECT  5.625 0.84 6.875 0.94 ;
      RECT  6.77 0.94 6.875 1.24 ;
      RECT  6.77 1.24 7.46 1.36 ;
      RECT  0.28 0.435 1.515 0.565 ;
      RECT  1.385 0.565 1.515 0.77 ;
      RECT  1.385 0.77 2.845 0.9 ;
      RECT  1.385 0.9 1.515 1.035 ;
      RECT  0.34 1.035 1.515 1.165 ;
      RECT  0.34 1.165 0.45 1.285 ;
      RECT  1.84 0.455 4.865 0.585 ;
      RECT  3.4 0.585 3.53 1.035 ;
      RECT  1.84 1.035 3.53 1.165 ;
      RECT  3.4 1.165 3.53 1.55 ;
      RECT  3.4 1.55 6.45 1.56 ;
      RECT  5.2 1.44 6.45 1.55 ;
      RECT  3.4 1.56 5.31 1.66 ;
      LAYER M2 ;
      RECT  1.375 0.55 5.11 0.65 ;
      RECT  1.375 0.95 3.76 1.05 ;
      LAYER V1 ;
      RECT  1.415 0.55 1.515 0.65 ;
      RECT  4.97 0.55 5.07 0.65 ;
      RECT  1.415 0.95 1.515 1.05 ;
      RECT  3.62 0.95 3.72 1.05 ;
  END
END SEN_EN2_S_6
#-----------------------------------------------------------------------
#      Cell        : SEN_EN2_S_8
#      Description : "2-Input exclusive NOR"
#      Equation    : X=!(A1^A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN2_S_8
  CLASS CORE ;
  FOREIGN SEN_EN2_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5064 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.15 0.71 9.905 0.93 ;
      RECT  9.15 0.93 9.25 1.09 ;
      RECT  5.15 0.71 6.05 0.905 ;
      RECT  5.95 0.905 6.05 0.95 ;
      RECT  5.95 0.95 6.19 1.05 ;
      LAYER M2 ;
      RECT  6.01 0.95 9.29 1.05 ;
      LAYER V1 ;
      RECT  9.15 0.95 9.25 1.05 ;
      RECT  6.05 0.95 6.15 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.741 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 10.4 1.85 ;
      RECT  0.59 1.255 0.71 1.75 ;
      RECT  1.11 1.255 1.23 1.75 ;
      RECT  1.63 1.255 1.75 1.75 ;
      RECT  2.15 1.21 2.27 1.75 ;
      RECT  2.67 1.255 2.79 1.75 ;
      RECT  3.19 1.255 3.31 1.75 ;
      RECT  3.71 1.255 3.83 1.75 ;
      RECT  4.23 1.255 4.35 1.75 ;
      RECT  8.595 1.21 8.71 1.75 ;
      RECT  9.105 1.45 9.235 1.75 ;
      RECT  9.66 1.21 9.78 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.4 0.05 ;
      RECT  0.585 0.05 0.715 0.345 ;
      RECT  1.105 0.05 1.235 0.345 ;
      RECT  1.625 0.05 1.755 0.345 ;
      RECT  8.85 0.05 8.975 0.36 ;
      RECT  9.365 0.05 9.495 0.36 ;
      RECT  9.885 0.05 10.015 0.36 ;
      RECT  2.665 0.05 2.795 0.365 ;
      RECT  3.185 0.05 3.315 0.365 ;
      RECT  3.705 0.05 3.835 0.365 ;
      RECT  4.225 0.05 4.345 0.365 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  2.15 0.05 2.27 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.435 0.22 8.76 0.35 ;
      RECT  8.63 0.35 8.76 0.65 ;
      RECT  7.28 0.65 8.76 0.78 ;
      RECT  7.28 0.78 7.45 1.11 ;
      RECT  6.51 1.11 8.33 1.29 ;
      RECT  6.51 1.29 6.61 1.34 ;
      RECT  4.925 1.34 6.61 1.46 ;
    END
    ANTENNADIFFAREA 1.611 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.54 0.44 8.53 0.56 ;
      RECT  6.54 0.56 6.66 0.675 ;
      RECT  6.28 0.675 6.66 0.795 ;
      RECT  6.28 0.795 6.4 1.14 ;
      RECT  4.695 0.91 4.795 1.14 ;
      RECT  4.695 1.14 6.4 1.25 ;
      RECT  0.28 0.435 2.05 0.565 ;
      RECT  1.88 0.565 2.05 0.75 ;
      RECT  1.88 0.75 3.715 0.92 ;
      RECT  1.88 0.92 2.05 1.035 ;
      RECT  0.34 1.035 2.05 1.165 ;
      RECT  0.34 1.165 0.45 1.255 ;
      RECT  8.865 0.45 10.32 0.57 ;
      RECT  8.865 0.57 8.97 0.87 ;
      RECT  7.54 0.87 8.97 0.97 ;
      RECT  8.85 0.97 8.97 1.24 ;
      RECT  8.85 1.24 9.54 1.36 ;
      RECT  2.36 0.455 6.425 0.585 ;
      RECT  3.93 0.585 4.57 0.625 ;
      RECT  4.4 0.625 4.57 0.995 ;
      RECT  3.93 0.995 4.57 1.035 ;
      RECT  2.36 1.035 4.57 1.165 ;
      RECT  4.44 1.165 4.57 1.55 ;
      RECT  4.44 1.55 8.505 1.56 ;
      RECT  6.75 1.44 8.505 1.55 ;
      RECT  4.44 1.56 6.86 1.66 ;
      LAYER M2 ;
      RECT  1.91 0.55 6.69 0.65 ;
      RECT  1.91 0.95 4.835 1.05 ;
      LAYER V1 ;
      RECT  1.95 0.55 2.05 0.65 ;
      RECT  6.55 0.55 6.65 0.65 ;
      RECT  1.95 0.95 2.05 1.05 ;
      RECT  4.695 0.95 4.795 1.05 ;
  END
END SEN_EN2_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_0P5
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_0P5
  CLASS CORE ;
  FOREIGN SEN_EN3_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0744 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.28 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.59 0.485 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  2.66 1.36 2.79 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  2.67 0.05 2.8 0.225 ;
      RECT  0.335 0.05 0.465 0.24 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.515 0.4 3.65 1.475 ;
    END
    ANTENNADIFFAREA 0.11 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.89 0.2 3.915 0.29 ;
      RECT  2.89 0.29 2.99 0.315 ;
      RECT  3.795 0.29 3.915 1.45 ;
      RECT  1.72 0.315 2.99 0.405 ;
      RECT  1.72 0.405 1.825 0.96 ;
      RECT  1.72 0.96 2.085 1.05 ;
      RECT  1.965 1.05 2.085 1.27 ;
      RECT  0.43 0.33 1.225 0.42 ;
      RECT  1.135 0.42 1.225 0.43 ;
      RECT  0.43 0.42 0.52 0.525 ;
      RECT  1.135 0.43 1.63 0.55 ;
      RECT  0.07 0.4 0.19 0.525 ;
      RECT  0.07 0.525 0.52 0.615 ;
      RECT  1.54 0.55 1.63 1.14 ;
      RECT  0.43 0.615 0.52 1.38 ;
      RECT  1.54 1.14 1.85 1.185 ;
      RECT  1.385 1.185 1.85 1.29 ;
      RECT  0.07 1.38 0.52 1.5 ;
      RECT  0.07 1.5 0.19 1.6 ;
      RECT  3.15 0.425 3.375 0.545 ;
      RECT  3.27 0.545 3.375 1.46 ;
      RECT  2.175 0.52 2.525 0.635 ;
      RECT  2.42 0.635 2.525 1.57 ;
      RECT  2.945 0.495 3.06 0.71 ;
      RECT  2.945 0.71 3.16 0.88 ;
      RECT  2.945 0.88 3.065 1.565 ;
      RECT  2.945 1.565 3.88 1.66 ;
      RECT  1.965 0.495 2.085 0.78 ;
      RECT  1.965 0.78 2.33 0.87 ;
      RECT  2.225 0.87 2.33 1.45 ;
      RECT  0.61 0.51 0.73 1.445 ;
      RECT  0.61 1.445 1.01 1.45 ;
      RECT  0.89 1.205 1.01 1.445 ;
      RECT  0.61 1.45 2.33 1.54 ;
      RECT  0.89 0.51 1.01 1.025 ;
      RECT  0.89 1.025 1.2 1.115 ;
      RECT  1.1 1.115 1.2 1.145 ;
      RECT  1.1 1.145 1.27 1.315 ;
      LAYER M2 ;
      RECT  1.06 1.15 3.415 1.25 ;
      LAYER V1 ;
      RECT  1.1 1.15 1.2 1.25 ;
      RECT  3.275 1.15 3.375 1.25 ;
  END
END SEN_EN3_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_1P5
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_1P5
  CLASS CORE ;
  FOREIGN SEN_EN3_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.65 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.73 0.71 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
      RECT  2.05 0.75 2.245 0.85 ;
      RECT  2.05 0.85 2.145 1.04 ;
      RECT  1.95 1.04 2.145 1.15 ;
      LAYER M2 ;
      RECT  2.065 0.75 3.87 0.85 ;
      LAYER V1 ;
      RECT  3.73 0.75 3.83 0.85 ;
      RECT  2.105 0.75 2.205 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2052 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.91 ;
      RECT  0.15 0.91 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.39 0.18 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.58 1.375 0.71 1.75 ;
      RECT  1.12 1.28 1.25 1.75 ;
      RECT  4.015 1.53 4.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.58 0.05 0.71 0.24 ;
      RECT  1.13 0.05 1.26 0.24 ;
      RECT  0.055 0.05 0.175 0.395 ;
      RECT  3.78 0.05 3.91 0.44 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.385 0.14 5.545 0.23 ;
      RECT  4.385 0.23 4.505 0.38 ;
      RECT  4.905 0.23 5.05 1.355 ;
      RECT  5.425 0.23 5.545 1.365 ;
    END
    ANTENNADIFFAREA 0.319 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.37 0.14 3.625 0.24 ;
      RECT  3.52 0.24 3.625 0.755 ;
      RECT  3.46 0.755 3.625 0.925 ;
      RECT  3.52 0.925 3.625 1.045 ;
      RECT  3.52 1.045 3.86 1.165 ;
      RECT  0.265 0.33 2.055 0.42 ;
      RECT  0.265 0.42 0.765 0.45 ;
      RECT  1.935 0.42 2.055 0.57 ;
      RECT  0.655 0.45 0.765 1.185 ;
      RECT  1.935 0.57 2.56 0.66 ;
      RECT  2.44 0.52 2.56 0.57 ;
      RECT  2.44 0.66 2.56 1.045 ;
      RECT  2.44 1.045 3.175 1.16 ;
      RECT  0.265 1.185 0.765 1.285 ;
      RECT  2.17 0.34 2.855 0.43 ;
      RECT  2.17 0.43 2.34 0.465 ;
      RECT  2.735 0.43 2.855 0.795 ;
      RECT  2.735 0.795 3.37 0.885 ;
      RECT  3.265 0.41 3.37 0.795 ;
      RECT  3.265 0.885 3.37 1.17 ;
      RECT  4.055 0.21 4.175 0.47 ;
      RECT  4.055 0.47 4.555 0.56 ;
      RECT  4.455 0.56 4.555 1.12 ;
      RECT  4.335 1.12 4.555 1.24 ;
      RECT  1.135 0.56 1.78 0.65 ;
      RECT  1.135 0.65 1.255 0.765 ;
      RECT  1.65 0.65 1.78 1.26 ;
      RECT  1.65 1.26 4.245 1.335 ;
      RECT  1.65 1.335 4.765 1.365 ;
      RECT  4.645 0.325 4.765 1.335 ;
      RECT  4.135 1.365 4.765 1.44 ;
      RECT  2.955 0.33 3.125 0.705 ;
      RECT  0.855 0.51 0.975 1.1 ;
      RECT  0.855 1.1 1.535 1.19 ;
      RECT  1.415 0.74 1.535 1.1 ;
      RECT  0.855 1.19 0.975 1.45 ;
      RECT  1.415 1.19 1.535 1.455 ;
      RECT  1.415 1.455 3.7 1.565 ;
      RECT  5.165 0.34 5.285 1.385 ;
      RECT  4.23 1.56 5.34 1.66 ;
      LAYER M2 ;
      RECT  0.825 0.55 3.095 0.65 ;
      RECT  3.225 0.55 5.305 0.65 ;
      LAYER V1 ;
      RECT  0.865 0.55 0.965 0.65 ;
      RECT  2.955 0.55 3.055 0.65 ;
      RECT  3.265 0.55 3.365 0.65 ;
      RECT  5.165 0.55 5.265 0.65 ;
  END
END SEN_EN3_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_3
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_3
  CLASS CORE ;
  FOREIGN SEN_EN3_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.65 0.89 ;
      RECT  7.15 0.89 7.25 0.945 ;
      RECT  7.55 0.89 7.65 1.09 ;
      RECT  6.75 0.945 7.25 1.045 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2061 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.665 2.25 0.91 ;
      RECT  2.15 0.91 2.45 0.945 ;
      RECT  2.15 0.945 3.09 1.09 ;
      RECT  4.26 0.715 4.835 0.85 ;
      LAYER M2 ;
      RECT  4.26 0.75 4.545 0.85 ;
      RECT  4.26 0.85 4.36 0.95 ;
      RECT  2.8 0.95 4.36 1.05 ;
      LAYER V1 ;
      RECT  2.84 0.95 2.94 1.05 ;
      RECT  4.405 0.75 4.505 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.393 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.405 0.45 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.845 1.21 0.965 1.75 ;
      RECT  1.365 1.25 1.485 1.75 ;
      RECT  5.245 1.415 5.37 1.75 ;
      RECT  5.765 1.21 5.885 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  1.36 0.05 1.49 0.35 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  5.225 0.05 5.355 0.445 ;
      RECT  0.845 0.05 0.965 0.59 ;
      RECT  5.765 0.05 5.885 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.545 0.39 6.665 0.44 ;
      RECT  6.545 0.44 7.85 0.56 ;
      RECT  7.75 0.56 7.85 1.315 ;
      RECT  6.47 1.315 7.85 1.405 ;
    END
    ANTENNADIFFAREA 0.55 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.665 0.17 3.295 0.26 ;
      RECT  2.665 0.26 2.785 0.35 ;
      RECT  3.185 0.26 3.295 1.14 ;
      RECT  3.185 1.14 3.4 1.18 ;
      RECT  2.75 1.18 3.4 1.285 ;
      RECT  3.295 1.285 3.4 1.31 ;
      RECT  6.3 0.175 6.925 0.265 ;
      RECT  6.805 0.265 6.925 0.35 ;
      RECT  6.3 0.265 6.45 0.37 ;
      RECT  6.35 0.37 6.45 1.035 ;
      RECT  6.265 1.035 6.45 1.125 ;
      RECT  6.265 1.125 6.375 1.495 ;
      RECT  6.265 1.495 6.95 1.6 ;
      RECT  3.385 0.23 4.06 0.35 ;
      RECT  3.385 0.35 3.49 0.83 ;
      RECT  3.385 0.83 3.6 0.945 ;
      RECT  3.49 0.945 3.6 1.45 ;
      RECT  3.49 1.45 4.17 1.56 ;
      RECT  3.49 1.56 3.6 1.57 ;
      RECT  1.625 0.23 2.32 0.35 ;
      RECT  1.625 0.35 1.745 0.44 ;
      RECT  1.06 0.44 1.745 0.56 ;
      RECT  1.625 0.56 1.745 1.04 ;
      RECT  1.05 1.04 1.745 1.16 ;
      RECT  1.625 1.16 1.745 1.465 ;
      RECT  1.625 1.465 2.29 1.555 ;
      RECT  2.12 1.555 2.29 1.57 ;
      RECT  2.12 1.57 3.6 1.66 ;
      RECT  4.36 0.23 5.05 0.35 ;
      RECT  4.93 0.35 5.05 0.945 ;
      RECT  4.93 0.945 5.155 1.065 ;
      RECT  5.04 1.065 5.155 1.45 ;
      RECT  4.495 1.45 5.155 1.57 ;
      RECT  7.315 0.23 8.05 0.35 ;
      RECT  7.94 0.35 8.05 1.495 ;
      RECT  7.375 1.495 8.05 1.6 ;
      RECT  2.915 0.35 3.095 0.44 ;
      RECT  1.885 0.44 3.095 0.56 ;
      RECT  1.885 0.56 2.005 1.255 ;
      RECT  1.885 1.255 2.59 1.375 ;
      RECT  2.47 1.375 3.21 1.48 ;
      RECT  0.065 0.31 0.185 0.45 ;
      RECT  0.065 0.45 0.705 0.54 ;
      RECT  0.585 0.54 0.705 0.785 ;
      RECT  0.585 0.785 1.505 0.895 ;
      RECT  0.585 0.895 0.705 1.225 ;
      RECT  0.065 1.225 0.705 1.315 ;
      RECT  0.065 1.315 0.185 1.45 ;
      RECT  3.605 0.44 4.84 0.56 ;
      RECT  3.74 0.56 3.86 1.24 ;
      RECT  3.74 1.24 4.925 1.36 ;
      RECT  4.285 1.36 4.385 1.49 ;
      RECT  6.055 0.19 6.175 0.565 ;
      RECT  6.055 0.565 6.26 0.735 ;
      RECT  6.055 0.735 6.175 1.13 ;
      RECT  6.025 1.13 6.175 1.315 ;
      RECT  6.54 0.705 6.985 0.815 ;
      RECT  6.54 0.815 6.63 1.135 ;
      RECT  6.54 1.135 7.46 1.225 ;
      RECT  7.36 0.99 7.46 1.135 ;
      RECT  2.525 0.705 3.095 0.85 ;
      RECT  3.97 0.675 4.08 0.945 ;
      RECT  3.97 0.945 4.84 1.055 ;
      RECT  5.505 0.31 5.625 1.325 ;
      LAYER M2 ;
      RECT  2.915 0.35 6.49 0.45 ;
      RECT  0.565 0.55 5.07 0.65 ;
      RECT  2.91 0.75 4.115 0.85 ;
      RECT  4.66 0.95 5.645 1.05 ;
      RECT  4.245 1.35 8.085 1.45 ;
      LAYER V1 ;
      RECT  2.955 0.35 3.055 0.45 ;
      RECT  6.35 0.35 6.45 0.45 ;
      RECT  0.605 0.55 0.705 0.65 ;
      RECT  3.195 0.55 3.295 0.65 ;
      RECT  4.93 0.55 5.03 0.65 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  3.975 0.75 4.075 0.85 ;
      RECT  4.7 0.95 4.8 1.05 ;
      RECT  5.505 0.95 5.605 1.05 ;
      RECT  4.285 1.35 4.385 1.45 ;
      RECT  7.945 1.35 8.045 1.45 ;
  END
END SEN_EN3_3
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_6
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_6
  CLASS CORE ;
  FOREIGN SEN_EN3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.95 0.51 12.05 0.71 ;
      RECT  10.515 0.71 12.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3834 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 0.71 9.12 0.935 ;
      RECT  8.55 0.935 8.65 1.09 ;
      RECT  4.915 0.755 5.26 0.795 ;
      RECT  4.175 0.795 5.26 0.89 ;
      RECT  5.16 0.89 5.26 1.105 ;
      LAYER M2 ;
      RECT  5.12 0.95 8.69 1.05 ;
      LAYER V1 ;
      RECT  8.55 0.95 8.65 1.05 ;
      RECT  5.16 0.95 5.26 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7311 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.25 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 13.6 1.85 ;
      RECT  0.58 1.415 0.71 1.75 ;
      RECT  1.1 1.415 1.23 1.75 ;
      RECT  1.62 1.415 1.75 1.75 ;
      RECT  2.14 1.415 2.27 1.75 ;
      RECT  2.66 1.415 2.79 1.75 ;
      RECT  3.185 1.21 3.305 1.75 ;
      RECT  3.7 1.4 3.83 1.75 ;
      RECT  9.795 1.515 9.925 1.75 ;
      RECT  10.425 1.515 10.55 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 13.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
      RECT  11.85 1.75 11.95 1.85 ;
      RECT  12.45 1.75 12.55 1.85 ;
      RECT  13.05 1.75 13.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 13.6 0.05 ;
      RECT  9.885 0.05 10.015 0.29 ;
      RECT  10.425 0.05 10.555 0.29 ;
      RECT  3.7 0.05 3.83 0.35 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.1 0.05 1.23 0.385 ;
      RECT  1.62 0.05 1.75 0.385 ;
      RECT  2.14 0.05 2.27 0.385 ;
      RECT  2.66 0.05 2.79 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.185 0.05 3.305 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 13.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
      RECT  11.85 -0.05 11.95 0.05 ;
      RECT  12.45 -0.05 12.55 0.05 ;
      RECT  13.05 -0.05 13.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.87 0.23 12.26 0.35 ;
      RECT  12.14 0.35 12.26 0.54 ;
      RECT  12.14 0.54 13.3 0.655 ;
      RECT  13.15 0.655 13.3 1.34 ;
      RECT  10.885 1.34 13.3 1.455 ;
    END
    ANTENNADIFFAREA 1.027 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.42 0.24 6.705 0.36 ;
      RECT  4.42 0.36 4.6 0.45 ;
      RECT  12.35 0.33 13.535 0.45 ;
      RECT  13.415 0.45 13.535 1.545 ;
      RECT  10.615 1.35 10.795 1.45 ;
      RECT  10.69 1.45 10.795 1.545 ;
      RECT  10.69 1.545 13.535 1.66 ;
      RECT  6.795 0.35 9.305 0.47 ;
      RECT  6.795 0.47 6.91 0.5 ;
      RECT  9.2 0.47 9.305 0.56 ;
      RECT  5.73 0.5 6.91 0.62 ;
      RECT  9.2 0.56 9.85 0.665 ;
      RECT  6.795 0.62 6.91 1.215 ;
      RECT  4.665 1.215 8.25 1.335 ;
      RECT  4.195 0.44 4.315 0.55 ;
      RECT  4.195 0.55 5.45 0.595 ;
      RECT  4.69 0.475 5.45 0.55 ;
      RECT  4.195 0.595 4.79 0.65 ;
      RECT  5.35 0.595 5.45 1.0 ;
      RECT  5.35 1.0 6.45 1.12 ;
      RECT  3.42 0.44 4.085 0.56 ;
      RECT  3.965 0.56 4.085 1.14 ;
      RECT  3.395 1.14 4.085 1.26 ;
      RECT  0.275 0.475 1.75 0.595 ;
      RECT  1.65 0.595 1.75 0.78 ;
      RECT  1.65 0.78 2.855 0.9 ;
      RECT  1.65 0.9 1.75 1.195 ;
      RECT  0.275 1.195 1.75 1.315 ;
      RECT  1.845 0.475 3.095 0.595 ;
      RECT  2.995 0.595 3.095 1.195 ;
      RECT  1.845 1.195 3.095 1.315 ;
      RECT  7.0 0.56 8.45 0.68 ;
      RECT  7.0 0.68 7.115 0.9 ;
      RECT  8.35 0.68 8.45 1.215 ;
      RECT  8.35 1.215 9.355 1.335 ;
      RECT  5.54 0.51 5.64 0.77 ;
      RECT  5.54 0.77 6.695 0.88 ;
      RECT  12.25 0.775 13.04 0.895 ;
      RECT  12.25 0.895 12.35 0.98 ;
      RECT  10.135 0.575 10.305 0.665 ;
      RECT  10.135 0.665 10.235 0.98 ;
      RECT  10.135 0.98 12.35 1.07 ;
      RECT  10.135 1.07 10.28 1.245 ;
      RECT  10.405 1.16 12.97 1.25 ;
      RECT  10.405 1.25 10.495 1.335 ;
      RECT  7.245 0.14 9.565 0.26 ;
      RECT  9.445 0.26 9.565 0.38 ;
      RECT  9.445 0.38 10.555 0.44 ;
      RECT  9.445 0.44 11.86 0.47 ;
      RECT  10.455 0.47 11.86 0.56 ;
      RECT  9.94 0.47 10.045 1.26 ;
      RECT  9.445 1.26 10.045 1.335 ;
      RECT  9.445 1.335 10.495 1.425 ;
      RECT  9.445 1.425 9.565 1.44 ;
      RECT  7.25 1.44 9.565 1.56 ;
      RECT  4.415 1.29 4.525 1.425 ;
      RECT  4.415 1.425 6.71 1.545 ;
      LAYER M2 ;
      RECT  4.42 0.35 12.53 0.45 ;
      RECT  3.935 0.55 5.68 0.65 ;
      RECT  2.955 0.75 7.145 0.85 ;
      RECT  1.61 1.15 6.935 1.25 ;
      RECT  4.38 1.35 10.795 1.45 ;
      LAYER V1 ;
      RECT  4.46 0.35 4.56 0.45 ;
      RECT  12.39 0.35 12.49 0.45 ;
      RECT  3.975 0.55 4.075 0.65 ;
      RECT  5.54 0.55 5.64 0.65 ;
      RECT  2.995 0.75 3.095 0.85 ;
      RECT  5.35 0.75 5.45 0.85 ;
      RECT  7.005 0.75 7.105 0.85 ;
      RECT  1.65 1.15 1.75 1.25 ;
      RECT  6.795 1.15 6.895 1.25 ;
      RECT  4.42 1.35 4.52 1.45 ;
      RECT  10.655 1.35 10.755 1.45 ;
  END
END SEN_EN3_6
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_1
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_1
  CLASS CORE ;
  FOREIGN SEN_EN3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.555 0.54 1.655 0.96 ;
      RECT  0.995 0.54 1.095 0.985 ;
      LAYER M2 ;
      RECT  0.91 0.75 1.73 0.85 ;
      LAYER V1 ;
      RECT  1.555 0.75 1.655 0.85 ;
      RECT  0.995 0.75 1.095 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0927 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.29 1.59 0.5 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  2.215 1.59 2.425 1.75 ;
      RECT  3.51 1.215 3.66 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.305 0.05 0.515 0.21 ;
      RECT  2.18 0.05 2.39 0.4 ;
      RECT  3.515 0.05 3.66 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.15 3.93 0.6 ;
      RECT  3.75 0.6 3.85 1.2 ;
      RECT  3.75 1.2 3.93 1.65 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.605 0.14 1.835 0.23 ;
      RECT  1.635 0.23 1.835 0.4 ;
      RECT  0.605 0.23 0.725 0.45 ;
      RECT  1.745 0.4 1.835 1.07 ;
      RECT  0.635 0.45 0.725 1.3 ;
      RECT  1.71 1.07 1.835 1.32 ;
      RECT  0.58 1.3 0.725 1.53 ;
      RECT  0.045 0.16 0.215 0.3 ;
      RECT  0.045 0.3 0.49 0.39 ;
      RECT  0.39 0.39 0.49 0.59 ;
      RECT  0.39 0.59 0.535 1.05 ;
      RECT  0.39 1.05 0.49 1.27 ;
      RECT  0.34 1.27 0.49 1.41 ;
      RECT  0.045 1.41 0.49 1.5 ;
      RECT  0.045 1.5 0.19 1.62 ;
      RECT  1.925 0.17 2.09 0.4 ;
      RECT  1.925 0.4 2.015 1.2 ;
      RECT  1.925 1.2 2.17 1.3 ;
      RECT  2.48 0.18 2.68 0.4 ;
      RECT  2.585 0.4 2.68 0.74 ;
      RECT  2.585 0.74 2.76 0.97 ;
      RECT  2.585 0.97 2.68 1.06 ;
      RECT  2.54 1.06 2.68 1.3 ;
      RECT  1.115 0.32 1.285 0.43 ;
      RECT  1.195 0.43 1.285 1.2 ;
      RECT  1.105 1.2 1.285 1.235 ;
      RECT  1.105 1.235 1.32 1.48 ;
      RECT  1.375 0.32 1.545 0.43 ;
      RECT  1.375 0.43 1.465 1.07 ;
      RECT  1.375 1.07 1.62 1.16 ;
      RECT  1.41 1.16 1.62 1.45 ;
      RECT  3.255 0.315 3.425 0.545 ;
      RECT  3.335 0.545 3.425 0.675 ;
      RECT  3.335 0.675 3.66 0.765 ;
      RECT  3.57 0.765 3.66 1.035 ;
      RECT  3.29 1.035 3.66 1.125 ;
      RECT  3.29 1.125 3.39 1.27 ;
      RECT  3.22 1.27 3.39 1.6 ;
      RECT  3.03 0.36 3.165 0.59 ;
      RECT  3.03 0.59 3.13 0.855 ;
      RECT  3.03 0.855 3.46 0.945 ;
      RECT  3.03 0.945 3.13 1.62 ;
      RECT  2.77 0.37 2.94 0.61 ;
      RECT  2.85 0.61 2.94 1.29 ;
      RECT  2.77 1.29 2.94 1.41 ;
      RECT  1.71 1.41 2.94 1.5 ;
      RECT  1.71 1.5 1.8 1.57 ;
      RECT  0.815 0.32 1.025 0.43 ;
      RECT  0.815 0.43 0.905 1.24 ;
      RECT  0.815 1.24 1.015 1.47 ;
      RECT  0.925 1.47 1.015 1.57 ;
      RECT  0.925 1.57 1.8 1.66 ;
      LAYER M2 ;
      RECT  0.31 1.35 1.3 1.45 ;
      RECT  1.42 1.35 3.39 1.45 ;
      LAYER V1 ;
      RECT  0.39 1.35 0.49 1.45 ;
      RECT  1.145 1.35 1.245 1.45 ;
      RECT  1.48 1.35 1.58 1.45 ;
      RECT  3.22 1.35 3.32 1.45 ;
  END
END SEN_EN3_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_2
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_2
  CLASS CORE ;
  FOREIGN SEN_EN3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.84 0.75 4.25 0.97 ;
      RECT  2.76 0.68 3.075 0.89 ;
      RECT  2.93 0.89 3.075 1.13 ;
      LAYER M2 ;
      RECT  2.68 0.75 4.08 0.85 ;
      LAYER V1 ;
      RECT  3.88 0.75 3.98 0.85 ;
      RECT  2.77 0.75 2.87 0.85 ;
      RECT  2.97 0.75 3.07 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0882 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.875 0.52 2.07 0.68 ;
      RECT  1.575 0.68 2.07 0.89 ;
      RECT  1.76 0.89 2.07 0.9 ;
      RECT  1.76 0.9 2.05 1.04 ;
      RECT  1.155 0.675 1.295 1.09 ;
      RECT  0.785 0.37 0.885 0.98 ;
      LAYER M2 ;
      RECT  0.67 0.75 1.96 0.85 ;
      LAYER V1 ;
      RECT  1.575 0.75 1.675 0.85 ;
      RECT  1.775 0.75 1.875 0.85 ;
      RECT  1.17 0.75 1.27 0.85 ;
      RECT  0.785 0.75 0.885 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1854 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.2 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.49 0.47 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  2.91 1.44 3.09 1.75 ;
      RECT  4.17 1.495 4.38 1.75 ;
      RECT  4.79 1.21 4.945 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  4.25 0.05 4.455 0.37 ;
      RECT  0.3 0.05 0.47 0.39 ;
      RECT  2.76 0.05 2.93 0.4 ;
      RECT  4.79 0.05 4.945 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.15 4.68 0.59 ;
      RECT  4.55 0.59 4.65 1.21 ;
      RECT  4.55 1.21 4.68 1.65 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.605 0.16 2.475 0.25 ;
      RECT  2.35 0.25 2.475 0.39 ;
      RECT  0.605 0.25 0.695 1.215 ;
      RECT  2.35 0.39 2.44 1.01 ;
      RECT  2.35 1.01 2.46 1.22 ;
      RECT  0.56 1.215 0.695 1.64 ;
      RECT  3.255 0.16 3.95 0.25 ;
      RECT  3.775 0.25 3.95 0.4 ;
      RECT  3.255 0.25 3.39 0.41 ;
      RECT  3.775 0.4 3.865 0.57 ;
      RECT  3.66 0.57 3.865 0.66 ;
      RECT  3.66 0.66 3.75 1.08 ;
      RECT  3.66 1.08 4.26 1.2 ;
      RECT  3.66 1.2 3.785 1.31 ;
      RECT  1.58 0.34 2.26 0.43 ;
      RECT  1.58 0.43 1.77 0.59 ;
      RECT  2.16 0.43 2.26 1.13 ;
      RECT  1.58 1.0 1.67 1.13 ;
      RECT  1.58 1.13 2.26 1.22 ;
      RECT  2.075 1.22 2.26 1.37 ;
      RECT  0.055 0.175 0.21 0.48 ;
      RECT  0.055 0.48 0.515 0.59 ;
      RECT  0.34 0.59 0.515 0.985 ;
      RECT  0.34 0.985 0.44 1.31 ;
      RECT  0.055 1.31 0.44 1.4 ;
      RECT  0.055 1.4 0.21 1.625 ;
      RECT  3.48 0.34 3.685 0.48 ;
      RECT  3.48 0.48 3.57 1.26 ;
      RECT  2.73 1.26 3.57 1.35 ;
      RECT  3.29 1.35 3.57 1.54 ;
      RECT  2.73 1.35 2.82 1.55 ;
      RECT  0.975 0.35 1.245 0.565 ;
      RECT  0.975 0.565 1.065 1.09 ;
      RECT  0.82 1.09 1.065 1.18 ;
      RECT  0.82 1.18 1.0 1.55 ;
      RECT  0.82 1.55 2.82 1.64 ;
      RECT  3.02 0.16 3.16 0.5 ;
      RECT  3.02 0.5 3.26 0.59 ;
      RECT  3.165 0.59 3.26 0.695 ;
      RECT  3.165 0.695 3.39 0.935 ;
      RECT  3.165 0.935 3.36 1.17 ;
      RECT  4.02 0.465 4.19 0.51 ;
      RECT  4.02 0.51 4.44 0.66 ;
      RECT  4.35 0.66 4.44 1.31 ;
      RECT  3.875 1.31 4.44 1.4 ;
      RECT  3.875 1.4 4.08 1.54 ;
      RECT  1.335 0.35 1.485 0.565 ;
      RECT  1.385 0.565 1.485 1.27 ;
      RECT  1.09 1.27 1.485 1.31 ;
      RECT  1.09 1.31 1.985 1.4 ;
      RECT  1.09 1.4 1.265 1.46 ;
      RECT  1.79 1.4 1.985 1.46 ;
      RECT  2.53 0.465 2.67 0.665 ;
      RECT  2.55 0.665 2.67 0.98 ;
      RECT  2.55 0.98 2.78 1.17 ;
      RECT  2.55 1.17 2.64 1.36 ;
      RECT  2.425 1.36 2.64 1.46 ;
      LAYER M2 ;
      RECT  0.32 0.55 1.58 0.65 ;
      RECT  2.02 0.55 4.28 0.65 ;
      LAYER V1 ;
      RECT  0.415 0.55 0.515 0.65 ;
      RECT  1.385 0.55 1.485 0.65 ;
      RECT  2.16 0.55 2.26 0.65 ;
      RECT  4.08 0.55 4.18 0.65 ;
  END
END SEN_EN3_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_4
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_4
  CLASS CORE ;
  FOREIGN SEN_EN3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.675 0.58 6.855 0.975 ;
      RECT  5.225 0.51 5.525 0.89 ;
      LAYER M2 ;
      RECT  5.14 0.75 7.0 0.85 ;
      LAYER V1 ;
      RECT  6.715 0.75 6.815 0.85 ;
      RECT  5.225 0.75 5.325 0.85 ;
      RECT  5.425 0.75 5.525 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1512 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.315 0.71 4.17 0.86 ;
      RECT  3.315 0.86 3.455 1.0 ;
      RECT  1.34 0.71 1.78 0.91 ;
      LAYER M2 ;
      RECT  1.41 0.75 3.71 0.85 ;
      LAYER V1 ;
      RECT  3.315 0.75 3.415 0.85 ;
      RECT  3.515 0.75 3.615 0.85 ;
      RECT  1.48 0.75 1.58 0.85 ;
      RECT  1.68 0.75 1.78 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3708 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.21 0.22 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.55 1.39 0.74 1.75 ;
      RECT  1.07 1.21 1.26 1.75 ;
      RECT  4.53 1.51 4.735 1.75 ;
      RECT  5.195 1.515 5.405 1.75 ;
      RECT  7.36 1.215 7.51 1.75 ;
      RECT  7.845 1.21 8.02 1.75 ;
      RECT  8.38 1.21 8.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  0.55 0.05 0.74 0.41 ;
      RECT  5.145 0.05 5.325 0.42 ;
      RECT  1.06 0.05 1.21 0.44 ;
      RECT  0.055 0.05 0.22 0.59 ;
      RECT  4.625 0.05 4.815 0.59 ;
      RECT  7.325 0.05 7.51 0.59 ;
      RECT  7.845 0.05 8.02 0.59 ;
      RECT  8.38 0.05 8.545 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.11 0.2 8.29 0.59 ;
      RECT  8.11 0.59 8.25 0.7 ;
      RECT  7.615 0.195 7.75 0.7 ;
      RECT  7.615 0.7 8.25 1.1 ;
      RECT  8.11 1.1 8.25 1.21 ;
      RECT  7.615 1.1 7.75 1.6 ;
      RECT  8.11 1.21 8.29 1.6 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.3 0.145 4.53 0.235 ;
      RECT  3.9 0.235 4.53 0.25 ;
      RECT  2.255 0.235 2.475 0.305 ;
      RECT  1.3 0.235 1.39 0.53 ;
      RECT  3.9 0.25 4.03 0.415 ;
      RECT  4.41 0.25 4.53 0.95 ;
      RECT  0.83 0.2 0.97 0.53 ;
      RECT  0.83 0.53 1.39 0.62 ;
      RECT  0.83 0.62 0.98 0.68 ;
      RECT  0.89 0.68 0.98 1.03 ;
      RECT  3.615 0.95 4.53 1.04 ;
      RECT  0.83 1.03 1.755 1.12 ;
      RECT  3.615 1.04 3.785 1.21 ;
      RECT  1.59 1.12 1.755 1.435 ;
      RECT  0.83 1.12 0.98 1.6 ;
      RECT  1.69 0.325 2.145 0.395 ;
      RECT  1.69 0.395 3.79 0.415 ;
      RECT  2.825 0.325 3.79 0.395 ;
      RECT  1.69 0.415 2.945 0.44 ;
      RECT  2.055 0.44 2.945 0.485 ;
      RECT  2.825 0.485 2.945 0.865 ;
      RECT  2.13 0.865 3.045 0.955 ;
      RECT  2.13 0.955 2.32 1.11 ;
      RECT  2.945 0.955 3.045 1.26 ;
      RECT  2.11 1.11 2.32 1.29 ;
      RECT  2.13 1.29 2.295 1.435 ;
      RECT  5.415 0.195 5.865 0.405 ;
      RECT  5.615 0.405 5.715 1.025 ;
      RECT  5.3 1.025 5.715 1.135 ;
      RECT  6.805 0.32 7.035 0.475 ;
      RECT  6.945 0.475 7.035 1.065 ;
      RECT  6.36 1.065 7.035 1.155 ;
      RECT  6.36 1.155 6.74 1.28 ;
      RECT  6.36 1.28 6.555 1.44 ;
      RECT  0.31 0.16 0.46 0.5 ;
      RECT  0.31 0.5 0.66 0.59 ;
      RECT  0.56 0.59 0.66 0.755 ;
      RECT  0.56 0.755 0.77 0.945 ;
      RECT  0.56 0.945 0.66 1.07 ;
      RECT  0.56 1.07 0.74 1.21 ;
      RECT  0.31 1.21 0.74 1.3 ;
      RECT  0.31 1.3 0.46 1.64 ;
      RECT  4.125 0.36 4.295 0.505 ;
      RECT  3.135 0.505 4.295 0.595 ;
      RECT  3.135 0.595 3.225 1.09 ;
      RECT  3.135 1.09 3.44 1.37 ;
      RECT  2.645 1.06 2.785 1.37 ;
      RECT  2.645 1.37 4.03 1.46 ;
      RECT  3.885 1.22 4.03 1.37 ;
      RECT  6.225 0.36 6.405 0.665 ;
      RECT  5.805 0.665 6.405 0.755 ;
      RECT  5.805 0.755 5.975 1.245 ;
      RECT  5.31 1.245 5.975 1.31 ;
      RECT  4.345 1.31 5.975 1.335 ;
      RECT  4.345 1.335 5.4 1.4 ;
      RECT  4.345 1.4 4.435 1.55 ;
      RECT  1.48 0.37 1.6 0.53 ;
      RECT  1.48 0.53 1.955 0.575 ;
      RECT  1.48 0.575 2.715 0.62 ;
      RECT  1.87 0.62 2.715 0.665 ;
      RECT  1.87 0.665 2.005 1.55 ;
      RECT  1.35 1.21 1.5 1.55 ;
      RECT  1.35 1.55 4.435 1.64 ;
      RECT  2.41 1.205 2.555 1.55 ;
      RECT  7.125 0.745 7.505 0.95 ;
      RECT  7.125 0.95 7.23 1.55 ;
      RECT  5.955 0.14 7.235 0.23 ;
      RECT  5.955 0.23 6.69 0.25 ;
      RECT  7.125 0.23 7.235 0.59 ;
      RECT  6.495 0.25 6.69 0.445 ;
      RECT  5.955 0.25 6.13 0.575 ;
      RECT  6.495 0.445 6.585 0.845 ;
      RECT  6.15 0.845 6.585 0.935 ;
      RECT  6.15 0.935 6.27 1.55 ;
      RECT  5.525 1.44 5.735 1.55 ;
      RECT  5.525 1.55 7.23 1.64 ;
      RECT  4.92 0.2 5.04 0.98 ;
      RECT  4.815 0.98 5.04 1.13 ;
      RECT  4.145 1.13 5.04 1.22 ;
      RECT  4.145 1.22 4.235 1.455 ;
      LAYER M2 ;
      RECT  0.54 1.15 2.36 1.25 ;
      RECT  3.05 1.15 6.79 1.25 ;
      LAYER V1 ;
      RECT  0.64 1.15 0.74 1.25 ;
      RECT  2.165 1.15 2.265 1.25 ;
      RECT  3.14 1.15 3.24 1.25 ;
      RECT  3.34 1.15 3.44 1.25 ;
      RECT  6.36 1.15 6.46 1.25 ;
      RECT  6.56 1.15 6.66 1.25 ;
  END
END SEN_EN3_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_DG_1
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_DG_1
  CLASS CORE ;
  FOREIGN SEN_EN3_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 3.85 0.69 ;
      RECT  3.75 0.69 3.85 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.69 2.94 1.05 ;
      RECT  1.15 0.67 1.25 1.09 ;
      LAYER M2 ;
      RECT  1.11 0.75 2.89 0.85 ;
      LAYER V1 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0837 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.69 0.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.415 0.45 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.85 1.415 0.97 1.75 ;
      RECT  4.23 1.445 4.4 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  4.21 0.05 4.33 0.23 ;
      RECT  0.33 0.05 0.45 0.385 ;
      RECT  0.85 0.05 0.97 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.31 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.03 0.14 2.96 0.23 ;
      RECT  2.03 0.23 2.235 0.335 ;
      RECT  2.86 0.23 2.96 0.35 ;
      RECT  2.145 0.335 2.235 0.825 ;
      RECT  2.145 0.825 2.44 0.915 ;
      RECT  2.32 0.915 2.44 1.3 ;
      RECT  1.53 1.22 1.645 1.3 ;
      RECT  1.53 1.3 2.44 1.39 ;
      RECT  3.05 0.14 3.925 0.23 ;
      RECT  3.05 0.23 3.14 0.46 ;
      RECT  2.59 0.33 2.69 0.46 ;
      RECT  2.59 0.46 3.14 0.55 ;
      RECT  3.05 0.55 3.14 1.56 ;
      RECT  2.59 1.325 2.69 1.56 ;
      RECT  2.59 1.56 3.315 1.66 ;
      RECT  1.34 0.2 1.94 0.32 ;
      RECT  1.34 0.32 1.44 1.48 ;
      RECT  1.34 1.48 1.94 1.6 ;
      RECT  0.565 0.245 0.745 0.365 ;
      RECT  0.645 0.365 0.745 1.44 ;
      RECT  0.565 1.44 0.745 1.56 ;
      RECT  3.43 0.32 4.45 0.42 ;
      RECT  4.35 0.42 4.45 1.25 ;
      RECT  3.985 1.25 4.45 1.355 ;
      RECT  3.985 1.355 4.075 1.57 ;
      RECT  3.5 1.43 3.6 1.57 ;
      RECT  3.5 1.57 4.075 1.66 ;
      RECT  0.07 0.2 0.19 0.48 ;
      RECT  0.07 0.48 0.545 0.57 ;
      RECT  0.445 0.57 0.545 1.235 ;
      RECT  0.07 1.235 0.545 1.325 ;
      RECT  0.07 1.325 0.19 1.485 ;
      RECT  1.11 0.215 1.23 0.49 ;
      RECT  0.905 0.49 1.23 0.58 ;
      RECT  0.905 0.58 1.005 1.2 ;
      RECT  0.905 1.2 1.23 1.29 ;
      RECT  1.11 1.29 1.23 1.53 ;
      RECT  2.325 0.34 2.44 0.645 ;
      RECT  2.325 0.645 2.65 0.735 ;
      RECT  2.55 0.735 2.65 1.14 ;
      RECT  2.55 1.14 2.95 1.235 ;
      RECT  2.85 1.235 2.95 1.45 ;
      RECT  1.95 0.48 2.055 0.9 ;
      RECT  3.41 0.875 3.51 1.01 ;
      RECT  3.41 1.01 4.095 1.105 ;
      RECT  3.975 0.51 4.095 1.01 ;
      RECT  3.975 1.105 4.095 1.16 ;
      RECT  1.53 0.41 1.645 1.015 ;
      RECT  1.53 1.015 2.215 1.13 ;
      RECT  3.23 0.34 3.32 1.21 ;
      RECT  3.23 1.21 3.815 1.3 ;
      RECT  3.725 1.3 3.815 1.385 ;
      RECT  3.23 1.3 3.41 1.45 ;
      RECT  3.725 1.385 3.895 1.48 ;
      LAYER M2 ;
      RECT  0.865 0.55 2.09 0.65 ;
      RECT  0.405 0.95 2.69 1.05 ;
      RECT  0.605 1.15 2.465 1.25 ;
      RECT  1.3 1.35 3.43 1.45 ;
      LAYER V1 ;
      RECT  0.905 0.55 1.005 0.65 ;
      RECT  1.95 0.55 2.05 0.65 ;
      RECT  0.445 0.95 0.545 1.05 ;
      RECT  1.54 0.95 1.64 1.05 ;
      RECT  2.55 0.95 2.65 1.05 ;
      RECT  0.645 1.15 0.745 1.25 ;
      RECT  2.325 1.15 2.425 1.25 ;
      RECT  1.34 1.35 1.44 1.45 ;
      RECT  3.27 1.35 3.37 1.45 ;
  END
END SEN_EN3_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_DG_2
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_DG_2
  CLASS CORE ;
  FOREIGN SEN_EN3_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 3.85 0.69 ;
      RECT  3.55 0.69 3.65 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.67 2.85 0.73 ;
      RECT  2.645 0.73 2.85 0.9 ;
      RECT  2.75 0.9 2.85 1.09 ;
      RECT  1.15 0.67 1.25 1.09 ;
      LAYER M2 ;
      RECT  1.11 0.75 2.85 0.85 ;
      LAYER V1 ;
      RECT  2.71 0.75 2.81 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0927 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.69 0.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.415 0.45 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.85 1.415 0.97 1.75 ;
      RECT  2.94 1.585 3.06 1.75 ;
      RECT  4.255 1.585 4.375 1.75 ;
      RECT  4.815 1.415 4.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  2.94 0.05 3.06 0.215 ;
      RECT  4.27 0.05 4.36 0.215 ;
      RECT  0.33 0.05 0.45 0.385 ;
      RECT  0.85 0.05 0.97 0.385 ;
      RECT  4.81 0.05 4.94 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.53 0.51 4.85 0.69 ;
      RECT  4.75 0.69 4.85 1.11 ;
      RECT  4.535 1.11 4.85 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.96 0.14 2.835 0.205 ;
      RECT  1.865 0.205 2.835 0.23 ;
      RECT  1.865 0.23 2.07 0.345 ;
      RECT  1.98 0.345 2.07 0.69 ;
      RECT  1.98 0.69 2.275 0.78 ;
      RECT  2.155 0.78 2.275 1.17 ;
      RECT  2.145 1.17 2.275 1.26 ;
      RECT  2.16 1.26 2.275 1.375 ;
      RECT  3.73 0.17 3.85 0.31 ;
      RECT  3.73 0.31 4.285 0.4 ;
      RECT  4.195 0.4 4.285 0.785 ;
      RECT  4.195 0.785 4.625 0.895 ;
      RECT  4.195 0.895 4.285 1.35 ;
      RECT  3.705 1.35 4.285 1.455 ;
      RECT  1.57 0.2 1.775 0.32 ;
      RECT  1.57 0.32 1.66 0.785 ;
      RECT  1.57 0.785 1.7 0.875 ;
      RECT  1.61 0.875 1.7 1.31 ;
      RECT  1.61 1.31 1.785 1.53 ;
      RECT  2.97 0.305 3.615 0.32 ;
      RECT  2.39 0.32 3.615 0.41 ;
      RECT  2.97 0.41 3.615 0.42 ;
      RECT  2.97 0.42 3.06 1.39 ;
      RECT  2.39 1.39 3.06 1.395 ;
      RECT  2.39 1.395 3.285 1.495 ;
      RECT  3.195 1.495 3.285 1.545 ;
      RECT  3.195 1.545 4.145 1.66 ;
      RECT  0.565 0.245 0.745 0.365 ;
      RECT  0.645 0.365 0.745 1.44 ;
      RECT  0.565 1.44 0.745 1.56 ;
      RECT  1.11 0.215 1.23 0.49 ;
      RECT  0.905 0.49 1.23 0.58 ;
      RECT  0.905 0.58 1.005 1.2 ;
      RECT  0.905 1.2 1.23 1.29 ;
      RECT  1.11 1.29 1.23 1.53 ;
      RECT  2.16 0.32 2.275 0.5 ;
      RECT  2.16 0.5 2.485 0.59 ;
      RECT  2.385 0.59 2.485 1.195 ;
      RECT  2.385 1.195 2.835 1.3 ;
      RECT  0.045 0.48 0.545 0.6 ;
      RECT  0.445 0.6 0.545 1.205 ;
      RECT  0.045 1.205 0.545 1.325 ;
      RECT  1.79 0.435 1.89 0.855 ;
      RECT  1.365 0.41 1.48 0.95 ;
      RECT  1.34 0.95 1.52 1.05 ;
      RECT  3.22 0.51 3.34 0.99 ;
      RECT  3.22 0.99 3.915 1.08 ;
      RECT  3.815 0.78 3.915 0.99 ;
      RECT  3.22 1.08 3.34 1.26 ;
      RECT  4.005 0.49 4.105 1.17 ;
      RECT  3.47 1.17 4.105 1.26 ;
      RECT  3.47 1.26 3.59 1.35 ;
      RECT  3.4 1.35 3.59 1.45 ;
      RECT  1.34 1.15 1.52 1.455 ;
      RECT  1.875 0.945 2.055 1.57 ;
      LAYER M2 ;
      RECT  0.865 0.55 1.93 0.65 ;
      RECT  0.405 0.95 2.525 1.05 ;
      RECT  1.42 1.15 2.3 1.25 ;
      RECT  1.42 1.25 1.52 1.35 ;
      RECT  0.605 1.35 1.52 1.45 ;
      RECT  1.645 1.35 3.58 1.45 ;
      LAYER V1 ;
      RECT  0.905 0.55 1.005 0.65 ;
      RECT  1.79 0.55 1.89 0.65 ;
      RECT  0.445 0.95 0.545 1.05 ;
      RECT  1.38 0.95 1.48 1.05 ;
      RECT  1.915 0.95 2.015 1.05 ;
      RECT  2.385 0.95 2.485 1.05 ;
      RECT  2.16 1.15 2.26 1.25 ;
      RECT  0.645 1.35 0.745 1.45 ;
      RECT  1.38 1.35 1.48 1.45 ;
      RECT  1.685 1.35 1.785 1.45 ;
      RECT  3.44 1.35 3.54 1.45 ;
  END
END SEN_EN3_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_DG_3
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_DG_3
  CLASS CORE ;
  FOREIGN SEN_EN3_DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.715 0.51 4.05 0.69 ;
      RECT  3.715 0.69 3.885 0.715 ;
      LAYER M2 ;
      RECT  3.245 0.55 4.13 0.65 ;
      LAYER V1 ;
      RECT  3.75 0.55 3.85 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0759 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.815 0.71 3.115 0.9 ;
      RECT  1.34 0.67 1.44 1.09 ;
      LAYER M2 ;
      RECT  1.3 0.75 2.955 0.85 ;
      LAYER V1 ;
      RECT  2.815 0.75 2.915 0.85 ;
      RECT  1.34 0.75 1.44 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1239 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.415 0.175 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  0.575 1.415 0.695 1.75 ;
      RECT  1.07 1.45 1.24 1.75 ;
      RECT  3.175 1.585 3.295 1.75 ;
      RECT  4.46 1.44 4.56 1.75 ;
      RECT  4.965 1.415 5.085 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  3.18 0.05 3.295 0.215 ;
      RECT  4.405 0.05 4.525 0.215 ;
      RECT  0.575 0.05 0.695 0.345 ;
      RECT  0.055 0.05 0.175 0.36 ;
      RECT  1.095 0.05 1.215 0.365 ;
      RECT  4.965 0.05 5.085 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.68 0.51 5.33 0.68 ;
      RECT  4.68 0.68 5.25 0.69 ;
      RECT  5.15 0.69 5.25 1.015 ;
      RECT  5.15 1.015 5.33 1.11 ;
      RECT  4.685 1.11 5.33 1.185 ;
      RECT  4.685 1.185 5.25 1.29 ;
    END
    ANTENNADIFFAREA 0.356 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.19 0.14 3.06 0.205 ;
      RECT  2.095 0.205 3.06 0.23 ;
      RECT  2.095 0.23 2.3 0.335 ;
      RECT  2.21 0.335 2.3 0.71 ;
      RECT  2.21 0.71 2.505 0.8 ;
      RECT  2.385 0.8 2.505 1.35 ;
      RECT  3.66 0.23 3.83 0.305 ;
      RECT  3.23 0.305 3.83 0.32 ;
      RECT  2.62 0.32 3.83 0.42 ;
      RECT  2.62 0.42 3.34 0.44 ;
      RECT  3.23 0.44 3.34 1.375 ;
      RECT  2.62 1.375 3.34 1.395 ;
      RECT  2.62 1.395 3.5 1.495 ;
      RECT  3.41 1.495 3.5 1.545 ;
      RECT  3.41 1.545 4.36 1.66 ;
      RECT  4.19 1.54 4.36 1.545 ;
      RECT  1.805 0.2 2.005 0.32 ;
      RECT  1.805 0.32 1.905 1.31 ;
      RECT  1.805 1.31 2.005 1.49 ;
      RECT  3.92 0.305 4.505 0.42 ;
      RECT  4.415 0.42 4.505 0.785 ;
      RECT  4.415 0.785 5.045 0.895 ;
      RECT  4.415 0.895 4.505 1.22 ;
      RECT  3.92 1.22 4.505 1.325 ;
      RECT  1.355 0.215 1.46 0.49 ;
      RECT  1.15 0.49 1.46 0.58 ;
      RECT  1.15 0.58 1.25 1.2 ;
      RECT  1.15 1.2 1.46 1.29 ;
      RECT  1.355 1.29 1.46 1.53 ;
      RECT  2.39 0.33 2.505 0.53 ;
      RECT  2.39 0.53 2.715 0.62 ;
      RECT  2.615 0.62 2.715 1.165 ;
      RECT  2.615 1.165 3.05 1.285 ;
      RECT  0.29 0.435 0.71 0.555 ;
      RECT  0.62 0.555 0.71 0.73 ;
      RECT  0.62 0.73 0.845 0.9 ;
      RECT  0.62 0.9 0.72 1.205 ;
      RECT  0.29 1.205 0.72 1.325 ;
      RECT  0.81 0.435 1.035 0.555 ;
      RECT  0.935 0.555 1.035 1.22 ;
      RECT  0.84 1.22 1.035 1.35 ;
      RECT  0.84 1.35 0.96 1.49 ;
      RECT  1.995 0.425 2.12 0.845 ;
      RECT  3.465 0.51 3.57 0.86 ;
      RECT  3.465 0.86 4.13 0.95 ;
      RECT  4.025 0.78 4.13 0.86 ;
      RECT  3.465 0.95 3.565 1.26 ;
      RECT  4.225 0.51 4.325 1.04 ;
      RECT  3.685 1.04 4.325 1.13 ;
      RECT  3.685 1.13 3.805 1.35 ;
      RECT  3.615 1.35 3.805 1.45 ;
      RECT  1.615 0.41 1.715 1.09 ;
      RECT  1.55 1.18 1.705 1.555 ;
      RECT  2.115 0.95 2.295 1.58 ;
      LAYER M2 ;
      RECT  1.11 0.55 2.155 0.65 ;
      RECT  0.58 0.95 2.755 1.05 ;
      RECT  1.605 1.15 2.53 1.25 ;
      RECT  1.605 1.25 1.705 1.35 ;
      RECT  0.81 1.35 1.745 1.45 ;
      RECT  1.865 1.35 3.795 1.45 ;
      LAYER V1 ;
      RECT  1.15 0.55 1.25 0.65 ;
      RECT  2.015 0.55 2.115 0.65 ;
      RECT  0.62 0.95 0.72 1.05 ;
      RECT  1.615 0.95 1.715 1.05 ;
      RECT  2.155 0.95 2.255 1.05 ;
      RECT  2.615 0.95 2.715 1.05 ;
      RECT  2.39 1.15 2.49 1.25 ;
      RECT  0.85 1.35 0.95 1.45 ;
      RECT  1.605 1.35 1.705 1.45 ;
      RECT  1.905 1.35 2.005 1.45 ;
      RECT  3.655 1.35 3.755 1.45 ;
  END
END SEN_EN3_DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_DG_4
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_DG_4
  CLASS CORE ;
  FOREIGN SEN_EN3_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.6 0.51 4.05 0.68 ;
      RECT  3.6 0.68 3.69 0.89 ;
      LAYER M2 ;
      RECT  3.185 0.55 4.07 0.65 ;
      LAYER V1 ;
      RECT  3.67 0.55 3.77 0.65 ;
      RECT  3.87 0.55 3.97 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.755 0.71 3.055 0.9 ;
      RECT  1.34 0.67 1.44 1.09 ;
      LAYER M2 ;
      RECT  1.3 0.75 2.895 0.85 ;
      LAYER V1 ;
      RECT  2.755 0.75 2.855 0.85 ;
      RECT  1.34 0.75 1.44 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.36 1.31 4.53 1.4 ;
      RECT  4.435 1.4 4.53 1.75 ;
      RECT  0.055 1.415 0.175 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.575 1.415 0.695 1.75 ;
      RECT  1.07 1.45 1.24 1.75 ;
      RECT  3.115 1.585 3.235 1.75 ;
      RECT  4.905 1.415 5.025 1.75 ;
      RECT  5.42 1.44 5.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  3.12 0.05 3.235 0.215 ;
      RECT  4.345 0.05 4.465 0.215 ;
      RECT  0.575 0.05 0.695 0.345 ;
      RECT  0.055 0.05 0.175 0.36 ;
      RECT  1.095 0.05 1.215 0.365 ;
      RECT  5.42 0.05 5.545 0.365 ;
      RECT  4.905 0.05 5.025 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.62 0.51 5.45 0.69 ;
      RECT  5.35 0.69 5.45 1.11 ;
      RECT  4.625 1.11 5.45 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.13 0.14 3.03 0.205 ;
      RECT  2.035 0.205 3.03 0.23 ;
      RECT  2.035 0.23 2.24 0.335 ;
      RECT  2.15 0.335 2.24 0.71 ;
      RECT  2.15 0.71 2.445 0.8 ;
      RECT  2.325 0.8 2.445 1.35 ;
      RECT  3.6 0.23 3.77 0.305 ;
      RECT  3.17 0.305 3.77 0.32 ;
      RECT  2.56 0.32 3.77 0.42 ;
      RECT  2.56 0.42 3.28 0.44 ;
      RECT  3.17 0.44 3.28 1.375 ;
      RECT  2.56 1.375 3.28 1.395 ;
      RECT  2.56 1.395 3.44 1.495 ;
      RECT  3.35 1.495 3.44 1.545 ;
      RECT  3.35 1.545 4.33 1.66 ;
      RECT  1.745 0.2 1.945 0.32 ;
      RECT  1.745 0.32 1.845 1.35 ;
      RECT  1.745 1.35 1.985 1.45 ;
      RECT  3.86 0.305 4.475 0.42 ;
      RECT  4.385 0.42 4.475 0.785 ;
      RECT  4.385 0.785 4.985 0.895 ;
      RECT  4.385 0.895 4.475 1.13 ;
      RECT  4.14 1.13 4.475 1.22 ;
      RECT  4.14 1.22 4.23 1.365 ;
      RECT  3.86 1.365 4.23 1.455 ;
      RECT  1.355 0.19 1.46 0.49 ;
      RECT  1.15 0.49 1.46 0.58 ;
      RECT  1.15 0.58 1.25 1.2 ;
      RECT  1.15 1.2 1.46 1.29 ;
      RECT  1.355 1.29 1.46 1.61 ;
      RECT  2.33 0.33 2.445 0.53 ;
      RECT  2.33 0.53 2.655 0.62 ;
      RECT  2.555 0.62 2.655 1.165 ;
      RECT  2.555 1.165 2.99 1.285 ;
      RECT  0.29 0.435 0.71 0.555 ;
      RECT  0.62 0.555 0.71 0.755 ;
      RECT  0.62 0.755 0.845 0.925 ;
      RECT  0.62 0.925 0.72 1.205 ;
      RECT  0.29 1.205 0.72 1.325 ;
      RECT  0.81 0.435 1.035 0.555 ;
      RECT  0.935 0.555 1.035 1.22 ;
      RECT  0.84 1.22 1.035 1.35 ;
      RECT  0.84 1.35 0.96 1.49 ;
      RECT  4.17 0.51 4.295 0.68 ;
      RECT  4.195 0.68 4.295 0.95 ;
      RECT  3.96 0.95 4.295 1.04 ;
      RECT  3.96 1.04 4.05 1.185 ;
      RECT  3.64 1.185 4.05 1.275 ;
      RECT  3.64 1.275 3.735 1.35 ;
      RECT  3.555 1.35 3.735 1.45 ;
      RECT  3.78 0.77 4.105 0.86 ;
      RECT  3.78 0.86 3.87 1.0 ;
      RECT  3.405 0.51 3.51 1.0 ;
      RECT  3.405 1.0 3.87 1.09 ;
      RECT  3.405 1.09 3.505 1.26 ;
      RECT  1.935 0.425 2.035 0.88 ;
      RECT  1.555 0.41 1.655 1.09 ;
      RECT  2.135 0.91 2.235 1.41 ;
      RECT  2.075 1.41 2.235 1.58 ;
      RECT  1.555 1.18 1.655 1.54 ;
      RECT  1.555 1.54 1.77 1.66 ;
      LAYER M2 ;
      RECT  1.11 0.55 2.075 0.65 ;
      RECT  0.58 0.95 2.695 1.05 ;
      RECT  1.555 1.15 2.47 1.25 ;
      RECT  1.555 1.25 1.655 1.35 ;
      RECT  0.81 1.35 1.695 1.45 ;
      RECT  1.8 1.35 3.735 1.45 ;
      LAYER V1 ;
      RECT  1.15 0.55 1.25 0.65 ;
      RECT  1.935 0.55 2.035 0.65 ;
      RECT  0.62 0.95 0.72 1.05 ;
      RECT  1.555 0.95 1.655 1.05 ;
      RECT  2.135 0.95 2.235 1.05 ;
      RECT  2.555 0.95 2.655 1.05 ;
      RECT  2.33 1.15 2.43 1.25 ;
      RECT  0.85 1.35 0.95 1.45 ;
      RECT  1.555 1.35 1.655 1.45 ;
      RECT  1.84 1.35 1.94 1.45 ;
      RECT  3.595 1.35 3.695 1.45 ;
  END
END SEN_EN3_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EN3_DG_8
#      Description : "3-Input exclusive NOR"
#      Equation    : X=!((A1^A2)^A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EN3_DG_8
  CLASS CORE ;
  FOREIGN SEN_EN3_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.51 6.45 0.71 ;
      RECT  5.73 0.71 6.45 0.8 ;
      RECT  5.73 0.8 6.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1914 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.67 4.85 1.09 ;
      RECT  2.84 0.685 2.94 1.105 ;
      LAYER M2 ;
      RECT  2.8 0.95 4.89 1.05 ;
      LAYER V1 ;
      RECT  4.75 0.95 4.85 1.05 ;
      RECT  2.84 0.95 2.94 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3174 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.4 1.85 ;
      RECT  0.58 1.415 0.71 1.75 ;
      RECT  1.1 1.415 1.23 1.75 ;
      RECT  1.62 1.415 1.75 1.75 ;
      RECT  2.145 1.21 2.265 1.75 ;
      RECT  5.52 1.44 5.645 1.75 ;
      RECT  7.15 1.21 7.255 1.75 ;
      RECT  7.65 1.41 7.78 1.75 ;
      RECT  8.17 1.41 8.3 1.75 ;
      RECT  8.69 1.41 8.82 1.75 ;
      RECT  9.215 1.21 9.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      RECT  5.5 0.05 5.67 0.305 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.1 0.05 1.23 0.385 ;
      RECT  1.62 0.05 1.75 0.385 ;
      RECT  7.65 0.05 7.78 0.39 ;
      RECT  8.17 0.05 8.3 0.39 ;
      RECT  8.69 0.05 8.82 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  2.145 0.05 2.265 0.59 ;
      RECT  7.15 0.05 7.255 0.59 ;
      RECT  9.215 0.05 9.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.37 0.49 9.06 0.62 ;
      RECT  8.89 0.62 9.06 1.11 ;
      RECT  7.35 1.11 9.06 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.77 0.23 7.06 0.35 ;
      RECT  6.97 0.35 7.06 0.77 ;
      RECT  6.97 0.77 8.715 0.895 ;
      RECT  6.97 0.895 7.06 1.55 ;
      RECT  5.735 1.55 7.06 1.66 ;
      RECT  2.63 0.24 3.815 0.36 ;
      RECT  3.695 0.36 3.815 0.41 ;
      RECT  2.63 0.36 2.74 1.44 ;
      RECT  2.63 1.44 3.84 1.56 ;
      RECT  4.0 0.35 4.9 0.47 ;
      RECT  4.0 0.47 4.1 0.5 ;
      RECT  3.41 0.5 4.1 0.62 ;
      RECT  4.0 0.62 4.1 1.215 ;
      RECT  2.865 1.215 4.36 1.335 ;
      RECT  6.545 0.44 6.88 0.56 ;
      RECT  6.79 0.56 6.88 1.34 ;
      RECT  5.735 1.34 6.88 1.455 ;
      RECT  0.275 0.475 1.23 0.595 ;
      RECT  1.14 0.595 1.23 0.78 ;
      RECT  1.14 0.78 1.865 0.9 ;
      RECT  1.685 0.75 1.865 0.78 ;
      RECT  1.14 0.9 1.23 1.195 ;
      RECT  0.275 1.195 1.23 1.315 ;
      RECT  1.34 0.475 2.055 0.595 ;
      RECT  1.955 0.595 2.055 1.195 ;
      RECT  1.32 1.195 2.055 1.315 ;
      RECT  2.865 0.475 3.13 0.595 ;
      RECT  3.03 0.595 3.13 1.0 ;
      RECT  3.03 1.0 3.605 1.12 ;
      RECT  4.19 0.56 4.58 0.68 ;
      RECT  4.48 0.68 4.58 1.215 ;
      RECT  4.48 1.215 4.9 1.335 ;
      RECT  3.22 0.51 3.32 0.785 ;
      RECT  3.22 0.785 3.905 0.895 ;
      RECT  6.595 0.715 6.695 0.895 ;
      RECT  6.35 0.895 6.695 0.98 ;
      RECT  5.24 0.575 5.435 0.68 ;
      RECT  5.24 0.68 5.34 0.98 ;
      RECT  5.24 0.98 6.695 0.985 ;
      RECT  5.24 0.985 6.45 1.07 ;
      RECT  5.24 1.07 5.385 1.17 ;
      RECT  6.595 1.08 6.7 1.16 ;
      RECT  5.51 1.16 6.7 1.25 ;
      RECT  5.51 1.25 5.6 1.26 ;
      RECT  3.905 0.14 5.135 0.26 ;
      RECT  5.015 0.26 5.135 0.395 ;
      RECT  5.015 0.395 5.66 0.44 ;
      RECT  5.015 0.44 6.23 0.485 ;
      RECT  5.56 0.485 6.23 0.56 ;
      RECT  5.015 0.485 5.135 1.26 ;
      RECT  5.015 1.26 5.6 1.35 ;
      RECT  5.015 1.35 5.135 1.44 ;
      RECT  3.93 1.44 5.135 1.56 ;
      RECT  2.405 0.455 2.525 1.225 ;
      LAYER M2 ;
      RECT  2.375 0.55 3.36 0.65 ;
      RECT  1.685 0.75 4.62 0.85 ;
      RECT  1.915 1.15 4.14 1.25 ;
      RECT  2.595 1.35 5.915 1.45 ;
      LAYER V1 ;
      RECT  2.415 0.55 2.515 0.65 ;
      RECT  3.22 0.55 3.32 0.65 ;
      RECT  1.725 0.75 1.825 0.85 ;
      RECT  3.03 0.75 3.13 0.85 ;
      RECT  4.48 0.75 4.58 0.85 ;
      RECT  1.955 1.15 2.055 1.25 ;
      RECT  4.0 1.15 4.1 1.25 ;
      RECT  2.635 1.35 2.735 1.45 ;
      RECT  5.775 1.35 5.875 1.45 ;
  END
END SEN_EN3_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_0P5
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_0P5
  CLASS CORE ;
  FOREIGN SEN_EO2_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.36 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0477 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.445 0.44 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.815 1.41 1.94 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.815 0.05 1.94 0.39 ;
      RECT  0.31 0.05 0.42 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.32 1.05 1.035 ;
      RECT  0.95 1.035 1.23 1.125 ;
      RECT  1.13 1.125 1.23 1.43 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.51 0.14 1.3 0.23 ;
      RECT  1.21 0.23 1.3 0.425 ;
      RECT  0.51 0.23 0.6 0.485 ;
      RECT  1.21 0.425 1.41 0.515 ;
      RECT  0.055 0.29 0.18 0.485 ;
      RECT  0.055 0.485 0.6 0.575 ;
      RECT  1.32 0.515 1.41 1.19 ;
      RECT  0.51 0.575 0.6 1.18 ;
      RECT  0.055 1.18 0.6 1.27 ;
      RECT  1.32 1.19 1.48 1.365 ;
      RECT  0.055 1.27 0.175 1.61 ;
      RECT  1.57 0.18 1.66 0.75 ;
      RECT  1.5 0.75 1.66 0.92 ;
      RECT  1.57 0.92 1.66 1.415 ;
      RECT  1.57 1.415 1.68 1.57 ;
      RECT  0.68 1.57 1.68 1.66 ;
      RECT  0.69 0.32 0.78 1.27 ;
      RECT  0.69 1.27 1.0 1.37 ;
      RECT  0.55 1.37 1.0 1.39 ;
      RECT  0.55 1.39 0.78 1.46 ;
  END
END SEN_EO2_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_1
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_1
  CLASS CORE ;
  FOREIGN SEN_EO2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.36 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.41 0.435 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.82 1.41 1.94 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.31 0.05 0.42 0.39 ;
      RECT  1.82 0.05 1.94 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.8 ;
      RECT  0.95 0.8 1.23 0.89 ;
      RECT  1.13 0.89 1.23 1.39 ;
    END
    ANTENNADIFFAREA 0.198 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.51 0.24 1.41 0.36 ;
      RECT  0.51 0.36 0.6 0.48 ;
      RECT  1.32 0.36 1.41 1.02 ;
      RECT  0.055 0.19 0.18 0.48 ;
      RECT  0.055 0.48 0.6 0.57 ;
      RECT  0.51 0.57 0.6 1.18 ;
      RECT  1.32 1.02 1.48 1.195 ;
      RECT  0.055 1.18 0.6 1.27 ;
      RECT  0.055 1.27 0.175 1.61 ;
      RECT  1.57 0.21 1.66 0.75 ;
      RECT  1.5 0.75 1.66 0.92 ;
      RECT  1.57 0.92 1.66 1.41 ;
      RECT  1.57 1.41 1.68 1.57 ;
      RECT  0.68 1.57 1.68 1.66 ;
      RECT  0.69 0.455 0.78 1.1 ;
      RECT  0.69 1.1 1.0 1.22 ;
      RECT  0.69 1.22 0.78 1.37 ;
      RECT  0.55 1.37 0.78 1.46 ;
  END
END SEN_EO2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_2
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_2
  CLASS CORE ;
  FOREIGN SEN_EO2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 2.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.18 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.57 1.41 0.7 1.75 ;
      RECT  1.09 1.41 1.22 1.75 ;
      RECT  2.825 1.41 2.945 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  0.57 0.05 0.7 0.345 ;
      RECT  1.09 0.05 1.21 0.365 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  2.825 0.05 2.945 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.3 0.225 2.485 0.345 ;
      RECT  2.35 0.345 2.485 0.4 ;
      RECT  2.35 0.4 2.45 1.31 ;
      RECT  1.855 1.31 2.485 1.38 ;
      RECT  1.325 1.38 2.485 1.49 ;
      RECT  1.325 1.49 1.445 1.61 ;
      RECT  2.365 1.49 2.485 1.61 ;
    END
    ANTENNADIFFAREA 0.46 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.29 0.44 0.65 0.56 ;
      RECT  0.55 0.56 0.65 0.785 ;
      RECT  0.55 0.785 1.0 0.885 ;
      RECT  0.55 0.885 0.65 1.195 ;
      RECT  0.26 1.195 1.735 1.285 ;
      RECT  2.015 0.44 2.25 0.56 ;
      RECT  2.015 0.56 2.115 0.74 ;
      RECT  0.78 0.46 1.925 0.58 ;
      RECT  1.115 0.58 1.205 1.0 ;
      RECT  1.835 0.58 1.925 1.095 ;
      RECT  0.78 1.0 1.205 1.105 ;
      RECT  1.835 1.095 2.25 1.215 ;
      RECT  1.565 0.71 1.675 0.95 ;
      RECT  1.565 0.95 1.745 1.05 ;
      RECT  2.555 0.49 2.66 1.25 ;
      LAYER M2 ;
      RECT  0.51 0.55 2.155 0.65 ;
      RECT  1.565 0.95 2.705 1.05 ;
      LAYER V1 ;
      RECT  0.55 0.55 0.65 0.65 ;
      RECT  2.015 0.55 2.115 0.65 ;
      RECT  1.605 0.95 1.705 1.05 ;
      RECT  2.555 0.95 2.655 1.05 ;
  END
END SEN_EO2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_3
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_3
  CLASS CORE ;
  FOREIGN SEN_EO2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 4.05 0.89 ;
      RECT  3.55 0.89 3.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.27 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.41 0.44 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.83 1.44 0.96 1.75 ;
      RECT  1.35 1.435 1.48 1.75 ;
      RECT  3.67 1.44 3.8 1.75 ;
      RECT  4.21 1.44 4.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  4.19 0.05 4.32 0.345 ;
      RECT  0.31 0.05 0.44 0.385 ;
      RECT  0.83 0.05 0.96 0.385 ;
      RECT  1.35 0.05 1.48 0.385 ;
      RECT  3.67 0.05 3.8 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.645 0.5 3.31 0.62 ;
      RECT  2.645 0.62 3.05 0.69 ;
      RECT  2.95 0.69 3.05 1.11 ;
      RECT  2.645 1.11 3.285 1.29 ;
      RECT  2.645 1.29 2.755 1.345 ;
      RECT  2.07 1.345 2.755 1.46 ;
      RECT  1.85 0.46 2.25 0.58 ;
      RECT  2.15 0.58 2.25 0.69 ;
      LAYER M2 ;
      RECT  2.11 0.55 2.785 0.65 ;
      LAYER V1 ;
      RECT  2.645 0.55 2.745 0.65 ;
      RECT  2.15 0.55 2.25 0.65 ;
    END
    ANTENNADIFFAREA 0.714 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.445 0.215 3.57 0.335 ;
      RECT  2.445 0.335 2.535 1.14 ;
      RECT  1.16 0.785 1.895 0.895 ;
      RECT  1.79 0.895 1.895 1.0 ;
      RECT  1.79 1.0 1.94 1.09 ;
      RECT  1.835 1.09 1.94 1.14 ;
      RECT  1.835 1.14 2.535 1.255 ;
      RECT  0.055 0.16 0.175 0.485 ;
      RECT  0.055 0.485 0.85 0.605 ;
      RECT  0.75 0.605 0.85 1.21 ;
      RECT  0.055 1.21 0.85 1.31 ;
      RECT  0.055 1.31 0.175 1.63 ;
      RECT  3.905 0.435 4.25 0.55 ;
      RECT  4.15 0.55 4.25 1.23 ;
      RECT  3.88 1.23 4.25 1.35 ;
      RECT  1.985 0.78 2.355 0.89 ;
      RECT  2.155 0.89 2.355 1.05 ;
      RECT  2.905 1.415 3.57 1.535 ;
      RECT  2.905 1.535 3.025 1.55 ;
      RECT  1.615 0.24 2.31 0.36 ;
      RECT  1.615 0.36 1.735 0.485 ;
      RECT  0.98 0.485 1.735 0.605 ;
      RECT  0.98 0.605 1.07 1.225 ;
      RECT  0.98 1.225 1.735 1.345 ;
      RECT  1.615 1.345 1.735 1.55 ;
      RECT  1.615 1.55 3.025 1.66 ;
      LAYER M2 ;
      RECT  0.71 0.95 1.935 1.05 ;
      RECT  2.155 0.95 4.29 1.05 ;
      LAYER V1 ;
      RECT  0.75 0.95 0.85 1.05 ;
      RECT  1.795 0.95 1.895 1.05 ;
      RECT  2.195 0.95 2.295 1.05 ;
      RECT  4.15 0.95 4.25 1.05 ;
  END
END SEN_EO2_3
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_4
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_4
  CLASS CORE ;
  FOREIGN SEN_EO2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 4.85 0.71 ;
      RECT  4.75 0.71 5.05 0.92 ;
      RECT  3.775 0.71 4.36 0.92 ;
      LAYER M2 ;
      RECT  3.98 0.75 5.09 0.85 ;
      LAYER V1 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
      RECT  4.02 0.75 4.12 0.85 ;
      RECT  4.22 0.75 4.32 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.36 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  0.59 1.255 0.71 1.75 ;
      RECT  1.11 1.255 1.23 1.75 ;
      RECT  1.63 1.255 1.75 1.75 ;
      RECT  2.15 1.24 2.27 1.75 ;
      RECT  4.69 1.41 4.81 1.75 ;
      RECT  5.21 1.41 5.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  0.585 0.05 0.715 0.345 ;
      RECT  1.105 0.05 1.235 0.345 ;
      RECT  1.625 0.05 1.755 0.365 ;
      RECT  2.145 0.05 2.265 0.365 ;
      RECT  4.69 0.05 4.81 0.39 ;
      RECT  5.21 0.05 5.33 0.39 ;
      RECT  0.07 0.05 0.19 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.355 0.225 4.57 0.345 ;
      RECT  4.46 0.345 4.57 0.51 ;
      RECT  4.46 0.51 4.65 0.615 ;
      RECT  4.55 0.615 4.65 1.195 ;
      RECT  4.46 1.195 4.65 1.29 ;
      RECT  4.46 1.29 4.58 1.31 ;
      RECT  3.55 1.31 4.58 1.38 ;
      RECT  2.38 1.38 4.58 1.49 ;
      RECT  2.38 1.49 2.5 1.61 ;
    END
    ANTENNADIFFAREA 0.884 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.95 0.37 5.07 0.48 ;
      RECT  4.95 0.48 5.25 0.59 ;
      RECT  5.15 0.59 5.25 1.17 ;
      RECT  4.89 1.17 5.25 1.29 ;
      RECT  0.305 0.44 1.255 0.56 ;
      RECT  1.155 0.56 1.255 0.785 ;
      RECT  1.155 0.785 1.93 0.885 ;
      RECT  1.155 0.885 1.255 1.04 ;
      RECT  0.34 1.04 1.255 1.16 ;
      RECT  0.34 1.16 0.45 1.26 ;
      RECT  3.575 0.44 4.37 0.56 ;
      RECT  3.575 0.56 3.675 0.69 ;
      RECT  1.345 0.46 3.485 0.58 ;
      RECT  2.17 0.58 2.26 1.04 ;
      RECT  3.395 0.58 3.485 1.095 ;
      RECT  1.345 1.04 2.26 1.145 ;
      RECT  3.395 1.095 4.35 1.215 ;
      RECT  2.63 0.825 3.16 0.935 ;
      RECT  3.06 0.935 3.16 0.95 ;
      RECT  3.06 0.95 3.285 1.05 ;
      RECT  2.36 0.91 2.46 1.14 ;
      RECT  2.36 1.14 3.305 1.26 ;
      LAYER M2 ;
      RECT  1.115 0.55 3.715 0.65 ;
      RECT  1.115 0.95 2.5 1.05 ;
      RECT  3.02 0.95 5.29 1.05 ;
      LAYER V1 ;
      RECT  1.155 0.55 1.255 0.65 ;
      RECT  3.575 0.55 3.675 0.65 ;
      RECT  1.155 0.95 1.255 1.05 ;
      RECT  2.36 0.95 2.46 1.05 ;
      RECT  3.12 0.95 3.22 1.05 ;
      RECT  5.15 0.95 5.25 1.05 ;
  END
END SEN_EO2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_5
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_5
  CLASS CORE ;
  FOREIGN SEN_EO2_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.96 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.85 0.89 ;
      RECT  5.35 0.89 5.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4125 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.415 0.44 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.83 1.415 0.96 1.75 ;
      RECT  1.355 1.21 1.475 1.75 ;
      RECT  1.87 1.435 2.0 1.75 ;
      RECT  2.39 1.435 2.52 1.75 ;
      RECT  5.395 1.44 5.525 1.75 ;
      RECT  6.035 1.44 6.165 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  0.31 0.05 0.44 0.385 ;
      RECT  0.83 0.05 0.96 0.385 ;
      RECT  1.87 0.05 2.0 0.385 ;
      RECT  2.39 0.05 2.52 0.385 ;
      RECT  5.695 0.05 5.825 0.395 ;
      RECT  6.215 0.05 6.34 0.45 ;
      RECT  1.355 0.05 1.475 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.435 0.5 5.165 0.62 ;
      RECT  4.435 0.62 4.655 0.69 ;
      RECT  4.545 0.69 4.655 1.11 ;
      RECT  4.015 1.11 5.14 1.29 ;
      RECT  4.015 1.29 4.125 1.345 ;
      RECT  2.865 1.345 4.125 1.46 ;
      RECT  2.865 0.46 4.1 0.58 ;
      RECT  3.75 0.58 4.1 0.69 ;
      LAYER M2 ;
      RECT  3.71 0.55 4.58 0.65 ;
      LAYER V1 ;
      RECT  4.44 0.55 4.54 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  3.95 0.55 4.05 0.65 ;
    END
    ANTENNADIFFAREA 0.978 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.23 0.215 5.43 0.335 ;
      RECT  4.23 0.335 4.34 0.91 ;
      RECT  3.82 0.91 4.34 1.02 ;
      RECT  3.82 1.02 3.925 1.14 ;
      RECT  2.2 0.785 2.985 0.895 ;
      RECT  2.875 0.895 2.985 1.14 ;
      RECT  2.875 1.14 3.925 1.255 ;
      RECT  0.055 0.17 0.175 0.485 ;
      RECT  0.055 0.485 1.215 0.605 ;
      RECT  1.095 0.605 1.215 0.785 ;
      RECT  1.095 0.785 1.93 0.895 ;
      RECT  1.095 0.895 1.215 1.195 ;
      RECT  0.055 1.195 1.215 1.315 ;
      RECT  0.055 1.315 0.175 1.62 ;
      RECT  5.395 0.485 6.105 0.6 ;
      RECT  6.005 0.6 6.105 1.23 ;
      RECT  5.645 1.23 6.105 1.35 ;
      RECT  3.075 0.785 3.65 0.895 ;
      RECT  3.55 0.895 3.65 0.95 ;
      RECT  3.55 0.95 3.73 1.05 ;
      RECT  4.215 1.415 4.905 1.535 ;
      RECT  4.215 1.535 4.335 1.55 ;
      RECT  2.655 0.24 3.865 0.36 ;
      RECT  2.655 0.36 2.775 0.485 ;
      RECT  1.565 0.485 2.775 0.605 ;
      RECT  2.02 0.605 2.11 1.225 ;
      RECT  1.59 1.225 2.775 1.345 ;
      RECT  2.655 1.345 2.775 1.55 ;
      RECT  2.655 1.55 4.335 1.66 ;
      LAYER M2 ;
      RECT  3.55 0.95 6.145 1.05 ;
      LAYER V1 ;
      RECT  3.59 0.95 3.69 1.05 ;
      RECT  6.005 0.95 6.105 1.05 ;
  END
END SEN_EO2_5
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_6
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_6
  CLASS CORE ;
  FOREIGN SEN_EO2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.25 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.51 6.85 0.71 ;
      RECT  6.75 0.71 7.25 0.91 ;
      RECT  5.55 0.71 6.4 0.91 ;
      LAYER M2 ;
      RECT  6.06 0.75 7.09 0.85 ;
      LAYER V1 ;
      RECT  6.75 0.75 6.85 0.85 ;
      RECT  6.95 0.75 7.05 0.85 ;
      RECT  6.1 0.75 6.2 0.85 ;
      RECT  6.3 0.75 6.4 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5004 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.59 1.255 0.71 1.75 ;
      RECT  1.11 1.255 1.23 1.75 ;
      RECT  1.63 1.21 1.75 1.75 ;
      RECT  2.15 1.255 2.27 1.75 ;
      RECT  2.67 1.255 2.79 1.75 ;
      RECT  3.19 1.255 3.31 1.75 ;
      RECT  7.025 1.45 7.155 1.75 ;
      RECT  7.565 1.45 7.695 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  0.585 0.05 0.715 0.345 ;
      RECT  1.105 0.05 1.235 0.345 ;
      RECT  7.285 0.05 7.415 0.355 ;
      RECT  2.145 0.05 2.275 0.365 ;
      RECT  2.665 0.05 2.795 0.365 ;
      RECT  3.185 0.05 3.305 0.365 ;
      RECT  6.765 0.05 6.895 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  1.63 0.05 1.75 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.395 0.22 6.65 0.35 ;
      RECT  6.52 0.35 6.65 1.11 ;
      RECT  4.95 1.11 6.65 1.29 ;
      RECT  4.95 1.29 5.05 1.35 ;
      RECT  3.89 1.35 5.05 1.46 ;
    END
    ANTENNADIFFAREA 1.141 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.96 0.44 6.43 0.56 ;
      RECT  4.96 0.56 5.08 0.675 ;
      RECT  4.72 0.675 5.08 0.795 ;
      RECT  4.72 0.795 4.84 1.14 ;
      RECT  3.62 0.91 3.72 1.14 ;
      RECT  3.62 1.14 4.84 1.26 ;
      RECT  6.98 0.45 7.67 0.56 ;
      RECT  7.55 0.56 7.67 1.24 ;
      RECT  6.74 1.24 7.67 1.36 ;
      RECT  0.28 0.435 1.515 0.565 ;
      RECT  1.385 0.565 1.515 0.77 ;
      RECT  1.385 0.77 2.845 0.9 ;
      RECT  1.385 0.9 1.515 1.035 ;
      RECT  0.34 1.035 1.515 1.165 ;
      RECT  0.34 1.165 0.45 1.285 ;
      RECT  1.84 0.455 4.865 0.585 ;
      RECT  3.4 0.585 3.53 1.035 ;
      RECT  1.84 1.035 3.53 1.165 ;
      RECT  3.4 1.165 3.53 1.55 ;
      RECT  3.4 1.55 6.45 1.56 ;
      RECT  5.19 1.44 6.45 1.55 ;
      RECT  3.4 1.56 5.3 1.66 ;
      RECT  3.84 0.82 4.52 0.93 ;
      RECT  4.42 0.93 4.52 0.95 ;
      RECT  4.42 0.95 4.63 1.05 ;
      LAYER M2 ;
      RECT  1.375 0.95 3.76 1.05 ;
      RECT  4.45 0.95 7.69 1.05 ;
      LAYER V1 ;
      RECT  1.415 0.95 1.515 1.05 ;
      RECT  3.62 0.95 3.72 1.05 ;
      RECT  4.49 0.95 4.59 1.05 ;
      RECT  7.55 0.95 7.65 1.05 ;
  END
END SEN_EO2_6
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_8
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_8
  CLASS CORE ;
  FOREIGN SEN_EO2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.35 0.51 8.45 0.71 ;
      RECT  8.35 0.71 8.89 0.87 ;
      RECT  7.18 0.87 8.89 0.98 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.666 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.215 0.19 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.59 1.255 0.71 1.75 ;
      RECT  1.11 1.255 1.23 1.75 ;
      RECT  1.63 1.255 1.75 1.75 ;
      RECT  2.15 1.215 2.27 1.75 ;
      RECT  2.67 1.255 2.79 1.75 ;
      RECT  3.19 1.255 3.31 1.75 ;
      RECT  3.71 1.255 3.83 1.75 ;
      RECT  4.26 1.565 4.435 1.75 ;
      RECT  8.38 1.215 8.495 1.75 ;
      RECT  8.895 1.45 9.015 1.75 ;
      RECT  9.415 1.215 9.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  0.59 0.05 0.71 0.345 ;
      RECT  1.11 0.05 1.23 0.345 ;
      RECT  1.63 0.05 1.75 0.345 ;
      RECT  8.38 0.05 8.495 0.36 ;
      RECT  8.895 0.05 9.015 0.36 ;
      RECT  2.67 0.05 2.79 0.365 ;
      RECT  3.19 0.05 3.31 0.365 ;
      RECT  3.71 0.05 3.83 0.365 ;
      RECT  9.415 0.05 9.535 0.56 ;
      RECT  4.23 0.05 4.35 0.565 ;
      RECT  0.07 0.05 0.19 0.585 ;
      RECT  2.15 0.05 2.27 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.845 0.51 8.05 0.69 ;
      RECT  6.92 0.69 7.09 1.11 ;
      RECT  4.75 0.51 6.475 0.69 ;
      RECT  6.3 0.69 6.475 1.11 ;
      RECT  6.3 1.11 8.06 1.29 ;
      RECT  6.3 1.29 6.45 1.34 ;
      RECT  4.74 1.34 6.45 1.46 ;
    END
    ANTENNADIFFAREA 1.466 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.585 0.24 8.29 0.36 ;
      RECT  6.585 0.36 6.7 0.505 ;
      RECT  4.505 0.235 6.21 0.365 ;
      RECT  4.505 0.365 4.64 0.68 ;
      RECT  2.385 0.455 4.105 0.585 ;
      RECT  3.93 0.585 4.105 0.68 ;
      RECT  3.93 0.68 4.64 0.82 ;
      RECT  3.93 0.82 4.105 1.035 ;
      RECT  2.385 1.035 4.105 1.165 ;
      RECT  3.96 1.165 4.105 1.34 ;
      RECT  3.96 1.34 4.64 1.47 ;
      RECT  4.525 1.47 4.64 1.55 ;
      RECT  4.525 1.55 8.29 1.56 ;
      RECT  6.545 1.44 8.29 1.55 ;
      RECT  4.525 1.56 6.655 1.66 ;
      RECT  1.88 0.31 2.05 0.435 ;
      RECT  0.305 0.435 2.05 0.565 ;
      RECT  1.88 0.565 2.05 0.75 ;
      RECT  1.88 0.75 3.715 0.92 ;
      RECT  1.88 0.92 2.05 1.035 ;
      RECT  0.34 1.035 2.05 1.165 ;
      RECT  0.34 1.165 0.45 1.285 ;
      RECT  8.595 0.45 9.275 0.57 ;
      RECT  9.155 0.57 9.275 1.24 ;
      RECT  8.61 1.24 9.275 1.36 ;
      RECT  4.865 0.86 5.89 0.95 ;
      RECT  4.865 0.95 5.975 0.98 ;
      RECT  5.79 0.98 5.975 1.05 ;
      RECT  4.505 0.91 4.625 1.14 ;
      RECT  4.505 1.14 6.21 1.25 ;
      LAYER M2 ;
      RECT  1.91 0.35 6.725 0.45 ;
      RECT  1.91 0.95 4.65 1.05 ;
      RECT  5.795 0.95 9.31 1.05 ;
      LAYER V1 ;
      RECT  1.95 0.35 2.05 0.45 ;
      RECT  6.585 0.35 6.685 0.45 ;
      RECT  1.95 0.95 2.05 1.05 ;
      RECT  4.51 0.95 4.61 1.05 ;
      RECT  5.835 0.95 5.935 1.05 ;
      RECT  9.17 0.95 9.27 1.05 ;
  END
END SEN_EO2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_S_2
#      Description : "2-Input exclusive OR, symmetric rise/fall"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_S_2
  CLASS CORE ;
  FOREIGN SEN_EO2_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.345 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.35 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0651 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.44 0.175 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.41 1.615 1.58 1.75 ;
      RECT  1.9 1.41 2.025 1.75 ;
      RECT  2.415 1.41 2.54 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.41 0.05 1.58 0.23 ;
      RECT  0.055 0.05 0.175 0.39 ;
      RECT  2.135 0.05 2.255 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.345 0.31 2.54 0.49 ;
      RECT  2.345 0.49 2.45 1.11 ;
      RECT  2.15 1.11 2.45 1.29 ;
    END
    ANTENNADIFFAREA 0.164 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.33 0.14 1.13 0.23 ;
      RECT  0.33 0.23 0.465 0.41 ;
      RECT  0.37 0.41 0.465 1.41 ;
      RECT  0.33 1.41 0.465 1.59 ;
      RECT  0.81 0.32 2.015 0.41 ;
      RECT  1.925 0.41 2.015 0.7 ;
      RECT  0.81 0.41 0.91 1.46 ;
      RECT  1.925 0.7 2.255 0.8 ;
      RECT  1.11 0.5 1.63 0.615 ;
      RECT  1.54 0.615 1.63 1.255 ;
      RECT  1.1 1.255 1.63 1.345 ;
      RECT  1.72 0.505 1.81 1.435 ;
      RECT  1.155 1.435 1.81 1.525 ;
      RECT  1.155 1.525 1.245 1.57 ;
      RECT  0.555 0.445 0.665 1.57 ;
      RECT  0.555 1.57 1.245 1.66 ;
  END
END SEN_EO2_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_S_4
#      Description : "2-Input exclusive OR, symmetric rise/fall"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_S_4
  CLASS CORE ;
  FOREIGN SEN_EO2_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.455 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.32 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.46 1.44 1.59 1.75 ;
      RECT  1.97 1.41 2.1 1.75 ;
      RECT  2.49 1.41 2.62 1.75 ;
      RECT  3.015 1.21 3.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  1.44 0.05 1.61 0.185 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  2.235 0.05 2.365 0.39 ;
      RECT  2.835 0.05 2.965 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.54 0.31 2.66 0.495 ;
      RECT  2.54 0.495 2.865 0.585 ;
      RECT  2.745 0.585 2.865 1.11 ;
      RECT  2.25 1.11 2.865 1.29 ;
    END
    ANTENNADIFFAREA 0.3 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.18 1.1 0.27 ;
      RECT  0.34 0.27 0.475 0.39 ;
      RECT  1.01 0.27 1.1 0.73 ;
      RECT  0.38 0.39 0.475 1.34 ;
      RECT  1.01 0.73 1.2 0.9 ;
      RECT  0.34 1.34 0.475 1.535 ;
      RECT  1.195 0.19 1.315 0.295 ;
      RECT  1.195 0.295 1.685 0.385 ;
      RECT  1.595 0.385 1.685 1.015 ;
      RECT  1.12 1.015 1.685 1.105 ;
      RECT  1.995 0.7 2.64 0.8 ;
      RECT  1.995 0.8 2.095 1.29 ;
      RECT  1.79 0.245 1.88 1.255 ;
      RECT  1.165 1.255 1.88 1.345 ;
      RECT  1.165 1.345 1.255 1.48 ;
      RECT  0.565 0.38 0.675 1.48 ;
      RECT  0.565 1.48 1.255 1.57 ;
      RECT  0.82 0.43 0.92 1.36 ;
      LAYER M2 ;
      RECT  0.78 1.15 2.135 1.25 ;
      LAYER V1 ;
      RECT  0.82 1.15 0.92 1.25 ;
      RECT  1.995 1.15 2.095 1.25 ;
  END
END SEN_EO2_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_S_8
#      Description : "2-Input exclusive OR, symmetric rise/fall"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_S_8
  CLASS CORE ;
  FOREIGN SEN_EO2_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.025 0.51 1.125 0.66 ;
      RECT  1.025 0.66 1.445 0.77 ;
      RECT  0.15 0.51 0.25 1.12 ;
      LAYER M2 ;
      RECT  0.11 0.55 1.165 0.65 ;
      LAYER V1 ;
      RECT  1.025 0.55 1.125 0.65 ;
      RECT  0.15 0.55 0.25 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  1.535 1.615 1.705 1.75 ;
      RECT  2.075 1.615 2.245 1.75 ;
      RECT  2.63 1.415 2.755 1.75 ;
      RECT  3.145 1.41 3.275 1.75 ;
      RECT  3.665 1.41 3.795 1.75 ;
      RECT  4.205 1.21 4.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  2.095 0.05 2.225 0.225 ;
      RECT  3.125 0.05 3.295 0.305 ;
      RECT  3.645 0.05 3.815 0.305 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  2.625 0.05 2.755 0.39 ;
      RECT  4.2 0.05 4.33 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.89 0.19 3.01 0.395 ;
      RECT  2.89 0.395 4.06 0.485 ;
      RECT  3.41 0.19 3.53 0.395 ;
      RECT  3.93 0.19 4.06 0.395 ;
      RECT  3.94 0.485 4.06 1.1 ;
      RECT  2.885 1.1 4.06 1.3 ;
    END
    ANTENNADIFFAREA 0.612 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.07 0.14 1.75 0.215 ;
      RECT  0.48 0.215 1.75 0.23 ;
      RECT  0.48 0.23 1.195 0.32 ;
      RECT  0.605 0.32 1.195 0.335 ;
      RECT  0.605 0.335 0.7 1.11 ;
      RECT  0.605 1.11 1.195 1.215 ;
      RECT  1.095 1.215 1.195 1.29 ;
      RECT  1.285 0.32 2.515 0.41 ;
      RECT  2.425 0.41 2.515 1.435 ;
      RECT  0.74 1.435 2.515 1.525 ;
      RECT  0.34 0.41 0.51 0.58 ;
      RECT  0.41 0.58 0.51 1.24 ;
      RECT  0.3 1.24 0.51 1.36 ;
      RECT  1.535 0.5 1.975 0.59 ;
      RECT  1.535 0.59 1.625 0.86 ;
      RECT  0.79 0.425 0.91 0.86 ;
      RECT  0.79 0.86 1.625 0.95 ;
      RECT  1.535 0.95 1.625 1.235 ;
      RECT  1.285 1.235 2.32 1.33 ;
      RECT  2.23 0.62 2.32 1.235 ;
      RECT  2.625 0.575 3.83 0.67 ;
      RECT  2.625 0.67 2.725 1.29 ;
      LAYER M2 ;
      RECT  1.055 1.15 2.765 1.25 ;
      LAYER V1 ;
      RECT  1.095 1.15 1.195 1.25 ;
      RECT  2.625 1.15 2.725 1.25 ;
  END
END SEN_EO2_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_DG_1
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_DG_1
  CLASS CORE ;
  FOREIGN SEN_EO2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.625 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.755 0.16 1.65 0.33 ;
      RECT  1.55 0.33 1.65 0.69 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.735 1.44 1.865 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.32 0.05 0.45 0.345 ;
      RECT  1.74 0.05 1.86 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.12 0.49 ;
      RECT  1.95 0.49 2.05 1.11 ;
      RECT  1.95 1.11 2.12 1.29 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.195 0.18 0.435 ;
      RECT  0.07 0.435 0.505 0.535 ;
      RECT  0.4 0.535 0.505 1.235 ;
      RECT  0.07 1.235 0.505 1.325 ;
      RECT  0.07 1.325 0.18 1.585 ;
      RECT  1.315 0.52 1.46 0.69 ;
      RECT  1.315 0.69 1.415 1.05 ;
      RECT  1.315 1.05 1.57 1.16 ;
      RECT  1.76 0.74 1.86 1.25 ;
      RECT  1.44 1.25 1.86 1.35 ;
      RECT  1.44 1.35 1.54 1.45 ;
      RECT  0.84 0.42 0.96 1.45 ;
      RECT  0.84 1.45 1.54 1.55 ;
      RECT  1.12 0.42 1.225 1.335 ;
      RECT  0.595 0.42 0.71 1.565 ;
      LAYER M2 ;
      RECT  0.36 1.15 1.26 1.25 ;
      LAYER V1 ;
      RECT  0.4 1.15 0.5 1.25 ;
      RECT  1.12 1.15 1.22 1.25 ;
  END
END SEN_EO2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_DG_16
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_DG_16
  CLASS CORE ;
  FOREIGN SEN_EO2_DG_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.72 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 4.85 1.13 ;
      RECT  3.42 0.49 3.52 0.71 ;
      RECT  2.91 0.71 3.52 0.89 ;
      LAYER M2 ;
      RECT  3.38 0.55 4.89 0.65 ;
      LAYER V1 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.42 0.55 3.52 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.105 1.21 1.225 1.75 ;
      RECT  1.62 1.44 1.75 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  4.71 1.48 4.88 1.75 ;
      RECT  5.23 1.48 5.4 1.75 ;
      RECT  5.77 1.41 5.9 1.75 ;
      RECT  6.29 1.41 6.42 1.75 ;
      RECT  6.81 1.41 6.94 1.75 ;
      RECT  7.33 1.41 7.46 1.75 ;
      RECT  7.85 1.41 7.98 1.75 ;
      RECT  8.37 1.41 8.5 1.75 ;
      RECT  8.89 1.41 9.02 1.75 ;
      RECT  9.415 1.21 9.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  0.58 0.05 0.71 0.35 ;
      RECT  7.33 0.05 7.46 0.35 ;
      RECT  7.85 0.05 7.98 0.35 ;
      RECT  8.37 0.05 8.5 0.35 ;
      RECT  8.89 0.05 9.02 0.35 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  4.73 0.05 4.86 0.39 ;
      RECT  5.77 0.05 5.9 0.39 ;
      RECT  6.29 0.05 6.42 0.39 ;
      RECT  6.81 0.05 6.94 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.105 0.05 1.225 0.59 ;
      RECT  5.255 0.05 5.375 0.59 ;
      RECT  9.415 0.05 9.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.345 0.44 8.845 0.49 ;
      RECT  5.515 0.49 8.845 0.51 ;
      RECT  5.515 0.51 9.275 0.69 ;
      RECT  8.53 0.69 8.85 1.04 ;
      RECT  7.625 1.04 8.85 1.11 ;
      RECT  5.515 1.11 9.275 1.29 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.44 0.99 0.56 ;
      RECT  0.89 0.56 0.99 0.785 ;
      RECT  0.89 0.785 1.945 0.895 ;
      RECT  0.89 0.895 0.99 1.225 ;
      RECT  0.28 1.225 0.99 1.35 ;
      RECT  1.315 0.45 3.33 0.56 ;
      RECT  2.335 0.56 2.425 1.24 ;
      RECT  1.315 1.24 4.385 1.35 ;
      RECT  3.61 0.44 4.385 0.56 ;
      RECT  3.61 0.56 3.71 1.04 ;
      RECT  2.64 0.91 2.74 1.04 ;
      RECT  2.64 1.04 3.71 1.15 ;
      RECT  3.88 0.785 4.25 0.895 ;
      RECT  4.15 0.895 4.25 1.09 ;
      RECT  5.255 0.8 8.385 0.91 ;
      RECT  5.255 0.91 7.505 0.97 ;
      RECT  5.255 0.97 5.425 1.22 ;
      RECT  2.36 0.24 4.605 0.35 ;
      RECT  4.485 0.35 4.605 1.22 ;
      RECT  4.485 1.22 5.425 1.39 ;
      RECT  4.485 1.39 4.59 1.44 ;
      RECT  2.36 1.44 4.59 1.56 ;
      RECT  4.995 0.415 5.14 1.03 ;
      RECT  4.97 1.03 5.14 1.12 ;
      LAYER M2 ;
      RECT  0.85 0.95 2.78 1.05 ;
      RECT  4.11 0.95 5.14 1.05 ;
      LAYER V1 ;
      RECT  0.89 0.95 0.99 1.05 ;
      RECT  2.64 0.95 2.74 1.05 ;
      RECT  4.15 0.95 4.25 1.05 ;
      RECT  5.0 0.95 5.1 1.05 ;
  END
END SEN_EO2_DG_16
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_DG_2
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_DG_2
  CLASS CORE ;
  FOREIGN SEN_EO2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.64 0.25 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.45 1.665 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.435 0.44 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.67 1.44 1.8 1.75 ;
      RECT  2.22 1.41 2.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.31 0.05 0.44 0.36 ;
      RECT  1.67 0.05 1.8 0.36 ;
      RECT  2.225 0.05 2.345 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.05 0.5 ;
      RECT  1.95 0.5 2.25 0.59 ;
      RECT  2.15 0.59 2.25 1.11 ;
      RECT  1.95 1.11 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.06 0.27 0.17 0.45 ;
      RECT  0.06 0.45 0.5 0.55 ;
      RECT  0.4 0.55 0.5 1.245 ;
      RECT  0.055 1.245 0.5 1.345 ;
      RECT  0.055 1.345 0.175 1.465 ;
      RECT  1.77 0.785 2.04 0.895 ;
      RECT  1.77 0.895 1.86 1.25 ;
      RECT  1.46 1.25 1.86 1.35 ;
      RECT  1.46 1.35 1.57 1.41 ;
      RECT  0.845 0.47 0.965 1.41 ;
      RECT  0.845 1.41 1.57 1.53 ;
      RECT  1.33 0.49 1.46 1.05 ;
      RECT  1.33 1.05 1.57 1.16 ;
      RECT  1.11 0.435 1.21 1.29 ;
      RECT  0.59 0.415 0.7 1.505 ;
      LAYER M2 ;
      RECT  0.36 1.15 1.25 1.25 ;
      LAYER V1 ;
      RECT  0.4 1.15 0.5 1.25 ;
      RECT  1.11 1.15 1.21 1.25 ;
  END
END SEN_EO2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_DG_4
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_DG_4
  CLASS CORE ;
  FOREIGN SEN_EO2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.65 0.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.805 0.51 2.05 0.69 ;
      RECT  1.805 0.69 1.915 0.96 ;
      RECT  0.78 0.45 0.88 0.955 ;
      LAYER M2 ;
      RECT  0.74 0.55 2.07 0.65 ;
      LAYER V1 ;
      RECT  1.93 0.55 2.03 0.65 ;
      RECT  0.78 0.55 0.88 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.45 0.45 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.91 1.465 2.08 1.75 ;
      RECT  2.45 1.41 2.58 1.75 ;
      RECT  3.015 1.21 3.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.32 0.05 0.45 0.345 ;
      RECT  1.905 0.05 2.035 0.39 ;
      RECT  2.45 0.05 2.58 0.39 ;
      RECT  3.015 0.05 3.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.85 0.69 ;
      RECT  2.75 0.69 2.85 1.11 ;
      RECT  2.205 1.11 2.85 1.29 ;
    END
    ANTENNADIFFAREA 0.476 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.33 0.185 0.44 ;
      RECT  0.065 0.44 0.51 0.56 ;
      RECT  0.41 0.56 0.51 1.24 ;
      RECT  0.07 1.24 0.51 1.36 ;
      RECT  0.07 1.36 0.18 1.465 ;
      RECT  0.97 0.445 1.24 0.555 ;
      RECT  0.97 0.555 1.06 1.045 ;
      RECT  0.835 1.045 1.06 1.135 ;
      RECT  0.835 1.135 0.955 1.29 ;
      RECT  2.025 0.78 2.64 0.89 ;
      RECT  2.025 0.89 2.115 1.255 ;
      RECT  0.795 0.23 1.475 0.34 ;
      RECT  1.37 0.34 1.475 1.255 ;
      RECT  1.045 1.255 2.115 1.365 ;
      RECT  1.15 0.645 1.28 1.09 ;
      RECT  1.615 0.215 1.715 1.16 ;
      RECT  0.6 0.415 0.69 1.46 ;
      RECT  0.6 1.46 1.525 1.57 ;
      LAYER M2 ;
      RECT  1.095 0.95 1.765 1.05 ;
      RECT  0.37 1.15 0.995 1.25 ;
      LAYER V1 ;
      RECT  1.15 0.95 1.25 1.05 ;
      RECT  1.615 0.95 1.715 1.05 ;
      RECT  0.41 1.15 0.51 1.25 ;
      RECT  0.855 1.15 0.955 1.25 ;
  END
END SEN_EO2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_DG_8
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_DG_8
  CLASS CORE ;
  FOREIGN SEN_EO2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.645 0.45 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.835 0.71 2.94 0.785 ;
      RECT  2.64 0.785 2.94 0.92 ;
      RECT  1.51 0.69 1.85 0.91 ;
      LAYER M2 ;
      RECT  1.47 0.75 2.98 0.85 ;
      LAYER V1 ;
      RECT  2.84 0.75 2.94 0.85 ;
      RECT  1.53 0.75 1.63 0.85 ;
      RECT  1.73 0.75 1.83 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.1 1.44 1.225 1.75 ;
      RECT  2.93 1.44 3.06 1.75 ;
      RECT  3.45 1.41 3.58 1.75 ;
      RECT  3.97 1.41 4.1 1.75 ;
      RECT  4.49 1.41 4.62 1.75 ;
      RECT  5.015 1.21 5.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.91 0.05 3.08 0.305 ;
      RECT  0.58 0.05 0.71 0.355 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  3.45 0.05 3.58 0.39 ;
      RECT  3.97 0.05 4.1 0.39 ;
      RECT  4.49 0.05 4.62 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.015 0.05 5.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.21 0.51 4.88 0.69 ;
      RECT  4.28 0.69 4.45 1.11 ;
      RECT  3.21 1.11 4.865 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.32 0.245 2.82 0.355 ;
      RECT  2.73 0.355 2.82 0.395 ;
      RECT  2.73 0.395 3.12 0.485 ;
      RECT  3.03 0.485 3.12 0.785 ;
      RECT  3.03 0.785 4.19 0.895 ;
      RECT  3.03 0.895 3.12 1.24 ;
      RECT  2.485 1.24 3.12 1.34 ;
      RECT  2.485 1.34 2.6 1.445 ;
      RECT  1.315 1.445 2.6 1.555 ;
      RECT  0.275 0.445 0.73 0.555 ;
      RECT  0.63 0.555 0.73 0.79 ;
      RECT  0.63 0.79 0.945 0.9 ;
      RECT  0.63 0.9 0.73 1.23 ;
      RECT  0.28 1.23 0.73 1.35 ;
      RECT  1.94 0.445 2.24 0.555 ;
      RECT  2.13 0.555 2.24 0.615 ;
      RECT  1.94 0.555 2.04 1.045 ;
      RECT  1.55 1.045 2.04 1.155 ;
      RECT  0.82 0.45 1.785 0.57 ;
      RECT  1.28 0.57 1.37 1.245 ;
      RECT  0.82 1.245 2.3 1.35 ;
      RECT  2.33 0.575 2.75 0.67 ;
      RECT  2.33 0.67 2.43 1.05 ;
      RECT  2.33 1.05 2.8 1.15 ;
      LAYER M2 ;
      RECT  0.59 0.55 2.11 0.65 ;
      LAYER V1 ;
      RECT  0.63 0.55 0.73 0.65 ;
      RECT  1.94 0.55 2.04 0.65 ;
  END
END SEN_EO2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_S_0P5
#      Description : "2-Input exclusive OR, symmetric rise/fall"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_S_0P5
  CLASS CORE ;
  FOREIGN SEN_EO2_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.335 0.93 ;
      RECT  1.15 0.93 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0492 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.28 0.205 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.125 1.495 1.295 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  1.17 0.05 1.29 0.595 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.44 0.755 0.56 ;
      RECT  0.55 0.56 0.65 1.285 ;
      RECT  0.55 1.285 0.77 1.405 ;
    END
    ANTENNADIFFAREA 0.122 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.14 1.08 0.23 ;
      RECT  0.98 0.23 1.08 0.38 ;
      RECT  0.34 0.23 0.46 1.435 ;
      RECT  0.87 0.48 0.99 1.225 ;
      RECT  1.425 0.4 1.545 1.315 ;
      RECT  0.91 1.315 1.545 1.405 ;
      RECT  0.91 1.405 1.0 1.55 ;
      RECT  0.44 1.55 1.0 1.66 ;
  END
END SEN_EO2_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_S_1
#      Description : "2-Input exclusive OR, symmetric rise/fall"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_S_1
  CLASS CORE ;
  FOREIGN SEN_EO2_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.285 0.71 0.45 0.925 ;
      RECT  0.35 0.925 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0633 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0927 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.345 1.385 0.475 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  2.015 1.41 2.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.33 0.05 0.455 0.385 ;
      RECT  1.78 0.05 1.91 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.25 0.69 ;
      RECT  1.15 0.69 1.25 1.11 ;
      RECT  1.15 1.11 1.365 1.29 ;
    END
    ANTENNADIFFAREA 0.196 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.545 0.245 1.435 0.365 ;
      RECT  0.545 0.365 0.635 0.495 ;
      RECT  1.345 0.365 1.435 0.8 ;
      RECT  0.065 0.495 0.635 0.585 ;
      RECT  0.54 0.585 0.635 0.925 ;
      RECT  0.065 0.585 0.185 1.26 ;
      RECT  1.345 0.8 1.605 0.89 ;
      RECT  1.495 0.89 1.605 1.325 ;
      RECT  1.525 0.285 1.645 0.6 ;
      RECT  1.525 0.6 1.79 0.69 ;
      RECT  1.695 0.69 1.79 1.44 ;
      RECT  1.695 1.44 1.925 1.46 ;
      RECT  0.915 0.78 1.015 1.46 ;
      RECT  0.915 1.46 1.925 1.56 ;
      RECT  0.725 0.48 0.825 1.34 ;
  END
END SEN_EO2_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_S_3
#      Description : "2-Input exclusive OR, symmetric rise/fall"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_S_3
  CLASS CORE ;
  FOREIGN SEN_EO2_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.72 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1899 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.73 0.71 4.25 0.925 ;
      RECT  4.15 0.925 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2778 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  1.365 1.24 1.485 1.75 ;
      RECT  3.685 1.21 3.805 1.75 ;
      RECT  4.205 1.21 4.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  3.685 0.05 3.81 0.385 ;
      RECT  4.205 0.05 4.325 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.835 0.24 3.58 0.36 ;
      RECT  3.35 0.36 3.45 1.11 ;
      RECT  2.71 1.11 3.45 1.29 ;
      RECT  2.71 1.29 2.815 1.35 ;
      RECT  2.08 1.35 2.815 1.47 ;
    END
    ANTENNADIFFAREA 0.633 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.385 0.185 0.485 ;
      RECT  0.065 0.485 0.935 0.605 ;
      RECT  0.845 0.605 0.935 0.71 ;
      RECT  0.845 0.71 1.16 0.93 ;
      RECT  0.845 0.93 0.935 1.195 ;
      RECT  0.065 1.195 0.935 1.315 ;
      RECT  0.065 1.315 0.185 1.415 ;
      RECT  2.53 0.485 3.26 0.605 ;
      RECT  3.155 0.605 3.26 0.69 ;
      RECT  2.53 0.605 2.62 1.13 ;
      RECT  1.43 0.71 1.925 0.93 ;
      RECT  1.835 0.93 1.925 1.13 ;
      RECT  1.835 1.13 2.62 1.25 ;
      RECT  3.54 0.485 4.11 0.605 ;
      RECT  3.54 0.605 3.64 1.03 ;
      RECT  3.54 1.03 4.06 1.12 ;
      RECT  3.945 1.12 4.06 1.465 ;
      RECT  2.025 0.71 2.44 0.93 ;
      RECT  2.915 1.415 3.595 1.535 ;
      RECT  2.915 1.535 3.035 1.57 ;
      RECT  1.05 0.485 2.315 0.6 ;
      RECT  1.05 0.6 1.34 0.605 ;
      RECT  1.25 0.605 1.34 1.03 ;
      RECT  1.055 1.03 1.745 1.15 ;
      RECT  1.625 1.15 1.745 1.57 ;
      RECT  1.625 1.57 3.035 1.66 ;
      LAYER M2 ;
      RECT  1.02 0.75 1.57 0.85 ;
      RECT  2.1 0.75 3.68 0.85 ;
      LAYER V1 ;
      RECT  1.06 0.75 1.16 0.85 ;
      RECT  1.43 0.75 1.53 0.85 ;
      RECT  2.14 0.75 2.24 0.85 ;
      RECT  2.34 0.75 2.44 0.85 ;
      RECT  3.54 0.75 3.64 0.85 ;
  END
END SEN_EO2_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_S_5
#      Description : "2-Input exclusive OR, symmetric rise/fall"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_S_5
  CLASS CORE ;
  FOREIGN SEN_EO2_S_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.06 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3165 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.51 5.45 0.71 ;
      RECT  4.745 0.71 5.66 0.82 ;
      RECT  4.745 0.82 5.25 0.89 ;
      RECT  5.55 0.82 5.66 0.91 ;
      RECT  5.55 0.91 6.05 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.456 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.42 1.415 0.55 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.94 1.415 1.07 1.75 ;
      RECT  1.465 1.21 1.585 1.75 ;
      RECT  1.985 1.24 2.105 1.75 ;
      RECT  2.505 1.24 2.625 1.75 ;
      RECT  5.35 1.41 5.48 1.75 ;
      RECT  5.88 1.41 6.01 1.75 ;
      RECT  6.4 1.41 6.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.42 0.05 0.55 0.385 ;
      RECT  0.94 0.05 1.07 0.385 ;
      RECT  1.98 0.05 2.11 0.385 ;
      RECT  2.5 0.05 2.63 0.385 ;
      RECT  5.88 0.05 6.01 0.385 ;
      RECT  1.465 0.05 1.585 0.59 ;
      RECT  6.405 0.05 6.525 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.545 0.46 5.26 0.58 ;
      RECT  4.545 0.58 4.655 1.11 ;
      RECT  4.125 1.11 5.25 1.29 ;
      RECT  4.125 1.29 4.235 1.345 ;
      RECT  5.15 1.29 5.25 1.49 ;
      RECT  2.98 1.345 4.235 1.46 ;
      RECT  2.975 0.46 4.25 0.58 ;
      RECT  3.95 0.58 4.25 0.69 ;
      LAYER M2 ;
      RECT  3.91 0.55 4.69 0.65 ;
      LAYER V1 ;
      RECT  4.55 0.55 4.65 0.65 ;
      RECT  3.95 0.55 4.05 0.65 ;
      RECT  4.15 0.55 4.25 0.65 ;
    END
    ANTENNADIFFAREA 1.032 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.34 0.24 5.54 0.36 ;
      RECT  4.34 0.36 4.45 0.91 ;
      RECT  3.925 0.91 4.45 1.02 ;
      RECT  3.925 1.02 4.035 1.14 ;
      RECT  2.31 0.75 3.095 0.895 ;
      RECT  2.985 0.895 3.095 1.14 ;
      RECT  2.985 1.14 4.035 1.255 ;
      RECT  0.115 0.485 1.325 0.605 ;
      RECT  1.205 0.605 1.325 0.75 ;
      RECT  1.205 0.75 2.04 0.895 ;
      RECT  1.205 0.895 1.325 1.195 ;
      RECT  0.115 1.195 1.325 1.315 ;
      RECT  5.575 0.485 6.26 0.605 ;
      RECT  6.145 0.605 6.26 1.2 ;
      RECT  5.35 0.91 5.45 1.2 ;
      RECT  5.35 1.2 6.26 1.29 ;
      RECT  5.615 1.29 5.735 1.535 ;
      RECT  6.145 1.29 6.26 1.535 ;
      RECT  3.185 0.785 3.755 0.895 ;
      RECT  3.655 0.895 3.755 0.95 ;
      RECT  3.655 0.95 3.835 1.05 ;
      RECT  4.325 1.415 5.02 1.535 ;
      RECT  4.325 1.535 4.445 1.55 ;
      RECT  2.765 0.24 3.98 0.36 ;
      RECT  2.765 0.36 2.885 0.485 ;
      RECT  1.68 0.485 2.885 0.605 ;
      RECT  2.13 0.605 2.22 1.03 ;
      RECT  1.68 1.03 2.885 1.15 ;
      RECT  2.765 1.15 2.885 1.55 ;
      RECT  2.765 1.55 4.445 1.66 ;
      LAYER M2 ;
      RECT  1.66 0.75 2.69 0.85 ;
      RECT  3.655 0.95 5.49 1.05 ;
      LAYER V1 ;
      RECT  1.7 0.75 1.8 0.85 ;
      RECT  1.9 0.75 2.0 0.85 ;
      RECT  2.35 0.75 2.45 0.85 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  3.695 0.95 3.795 1.05 ;
      RECT  5.35 0.95 5.45 1.05 ;
  END
END SEN_EO2_S_5
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_S_6
#      Description : "2-Input exclusive OR, symmetric rise/fall"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_S_6
  CLASS CORE ;
  FOREIGN SEN_EO2_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.25 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3798 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.98 0.71 7.45 0.935 ;
      RECT  6.98 0.935 7.08 1.09 ;
      RECT  5.55 0.71 6.45 0.935 ;
      RECT  6.35 0.935 6.45 1.09 ;
      LAYER M2 ;
      RECT  6.31 0.95 7.12 1.05 ;
      LAYER V1 ;
      RECT  6.98 0.95 7.08 1.05 ;
      RECT  6.35 0.95 6.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5553 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.0 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.625 1.21 1.745 1.75 ;
      RECT  2.145 1.24 2.265 1.75 ;
      RECT  2.665 1.24 2.785 1.75 ;
      RECT  3.185 1.24 3.305 1.75 ;
      RECT  7.015 1.41 7.145 1.75 ;
      RECT  7.58 1.21 7.7 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.1 0.05 1.23 0.385 ;
      RECT  2.14 0.05 2.27 0.385 ;
      RECT  2.66 0.05 2.79 0.385 ;
      RECT  3.18 0.05 3.31 0.385 ;
      RECT  6.78 0.05 6.91 0.385 ;
      RECT  7.3 0.05 7.43 0.385 ;
      RECT  7.82 0.05 7.945 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.625 0.05 1.745 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.41 0.225 6.67 0.355 ;
      RECT  6.54 0.355 6.67 1.18 ;
      RECT  4.95 1.11 6.255 1.18 ;
      RECT  4.95 1.18 6.67 1.3 ;
      RECT  3.825 1.3 6.67 1.31 ;
      RECT  3.825 1.31 5.08 1.43 ;
    END
    ANTENNADIFFAREA 1.27 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.25 0.465 6.45 0.585 ;
      RECT  5.25 0.585 5.38 0.735 ;
      RECT  4.73 0.735 5.38 0.865 ;
      RECT  4.73 0.865 4.86 1.07 ;
      RECT  2.62 0.735 3.745 0.905 ;
      RECT  3.615 0.905 3.745 1.07 ;
      RECT  3.615 1.07 4.86 1.2 ;
      RECT  1.835 0.475 4.91 0.595 ;
      RECT  2.4 0.595 4.91 0.605 ;
      RECT  2.4 0.605 2.53 1.02 ;
      RECT  2.4 1.02 3.525 1.03 ;
      RECT  1.835 1.03 3.525 1.15 ;
      RECT  3.395 1.15 3.525 1.53 ;
      RECT  3.395 1.53 6.385 1.535 ;
      RECT  5.17 1.415 6.385 1.53 ;
      RECT  3.395 1.535 5.3 1.66 ;
      RECT  6.76 0.485 7.735 0.6 ;
      RECT  6.76 0.6 6.89 1.185 ;
      RECT  6.76 1.185 7.45 1.305 ;
      RECT  0.275 0.485 1.49 0.605 ;
      RECT  1.36 0.605 1.49 0.735 ;
      RECT  1.36 0.735 2.31 0.905 ;
      RECT  1.36 0.905 1.49 1.19 ;
      RECT  0.275 1.19 1.49 1.31 ;
      RECT  3.945 0.71 4.63 0.89 ;
      LAYER M2 ;
      RECT  1.93 0.75 3.0 0.85 ;
      RECT  4.29 0.75 6.9 0.85 ;
      LAYER V1 ;
      RECT  1.97 0.75 2.07 0.85 ;
      RECT  2.17 0.75 2.27 0.85 ;
      RECT  2.66 0.75 2.76 0.85 ;
      RECT  2.86 0.75 2.96 0.85 ;
      RECT  4.33 0.75 4.43 0.85 ;
      RECT  4.53 0.75 4.63 0.85 ;
      RECT  6.76 0.75 6.86 0.85 ;
  END
END SEN_EO2_S_6
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_G_1
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_G_1
  CLASS CORE ;
  FOREIGN SEN_EO2_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.51 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.45 1.45 0.98 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.33 0.455 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.7 1.44 1.83 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  1.72 0.05 1.825 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.095 0.555 ;
      RECT  1.95 0.555 2.05 1.09 ;
      RECT  1.95 1.09 2.095 1.315 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.71 0.22 1.63 0.33 ;
      RECT  1.54 0.33 1.63 1.07 ;
      RECT  1.35 1.07 1.63 1.17 ;
      RECT  0.605 0.42 0.725 0.98 ;
      RECT  0.26 0.98 0.725 1.15 ;
      RECT  0.605 1.15 0.725 1.5 ;
      RECT  1.75 0.72 1.86 1.26 ;
      RECT  1.495 1.26 1.86 1.35 ;
      RECT  1.495 1.35 1.585 1.55 ;
      RECT  0.865 0.45 0.985 1.55 ;
      RECT  0.865 1.55 1.585 1.64 ;
      RECT  0.065 0.22 0.17 1.31 ;
      RECT  0.065 1.31 0.245 1.49 ;
      RECT  1.125 0.45 1.24 1.35 ;
      RECT  1.125 1.35 1.305 1.45 ;
      LAYER M2 ;
      RECT  0.105 1.35 1.305 1.45 ;
      LAYER V1 ;
      RECT  0.145 1.35 0.245 1.45 ;
      RECT  1.165 1.35 1.265 1.45 ;
  END
END SEN_EO2_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_G_2
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_G_2
  CLASS CORE ;
  FOREIGN SEN_EO2_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.515 0.71 0.65 1.145 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.315 0.925 ;
      RECT  1.15 0.925 1.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.85 1.465 2.02 1.75 ;
      RECT  2.395 1.41 2.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.32 0.05 0.45 0.345 ;
      RECT  2.4 0.05 2.53 0.39 ;
      RECT  1.875 0.05 1.995 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.135 0.51 2.45 0.69 ;
      RECT  2.35 0.69 2.45 1.11 ;
      RECT  2.14 1.11 2.45 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.31 0.69 0.45 ;
      RECT  0.315 0.45 0.69 0.54 ;
      RECT  0.315 0.54 0.405 0.755 ;
      RECT  0.26 0.755 0.405 0.925 ;
      RECT  0.315 0.925 0.405 1.235 ;
      RECT  0.315 1.235 0.7 1.325 ;
      RECT  0.59 1.325 0.7 1.55 ;
      RECT  0.59 1.55 1.5 1.64 ;
      RECT  1.33 1.465 1.5 1.55 ;
      RECT  0.97 0.445 1.265 0.565 ;
      RECT  0.97 0.565 1.06 1.015 ;
      RECT  0.835 1.015 1.06 1.105 ;
      RECT  0.835 1.105 0.955 1.31 ;
      RECT  1.95 0.785 2.24 0.895 ;
      RECT  1.95 0.895 2.05 1.25 ;
      RECT  0.79 0.245 1.5 0.355 ;
      RECT  1.41 0.355 1.5 1.24 ;
      RECT  1.045 1.24 1.5 1.25 ;
      RECT  1.045 1.25 2.05 1.36 ;
      RECT  0.78 0.445 0.88 0.925 ;
      RECT  0.07 0.44 0.17 1.11 ;
      RECT  0.07 1.11 0.225 1.29 ;
      RECT  1.61 0.21 1.72 1.16 ;
      LAYER M2 ;
      RECT  0.74 0.55 1.76 0.65 ;
      RECT  0.085 1.15 0.985 1.25 ;
      LAYER V1 ;
      RECT  0.78 0.55 0.88 0.65 ;
      RECT  1.62 0.55 1.72 0.65 ;
      RECT  0.125 1.15 0.225 1.25 ;
      RECT  0.845 1.15 0.945 1.25 ;
  END
END SEN_EO2_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_G_4
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_G_4
  CLASS CORE ;
  FOREIGN SEN_EO2_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.0 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.455 0.78 ;
      RECT  2.35 0.78 2.685 0.895 ;
      RECT  2.35 0.895 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.585 1.21 0.7 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  2.96 1.455 3.09 1.75 ;
      RECT  3.48 1.41 3.61 1.75 ;
      RECT  4.005 1.21 4.125 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  2.94 0.05 3.11 0.305 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  3.48 0.05 3.61 0.4 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  0.585 0.05 0.7 0.59 ;
      RECT  4.005 0.05 4.125 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.85 0.69 ;
      RECT  3.75 0.69 3.85 1.11 ;
      RECT  3.15 1.11 3.85 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.385 0.16 2.85 0.25 ;
      RECT  1.385 0.25 1.505 0.345 ;
      RECT  2.76 0.25 2.85 0.395 ;
      RECT  1.905 0.25 2.025 0.42 ;
      RECT  2.44 0.25 2.56 0.42 ;
      RECT  2.76 0.395 3.06 0.485 ;
      RECT  2.96 0.485 3.06 0.785 ;
      RECT  2.96 0.785 3.64 0.895 ;
      RECT  2.96 0.895 3.06 1.275 ;
      RECT  2.78 1.275 3.06 1.365 ;
      RECT  2.78 1.365 2.87 1.445 ;
      RECT  1.335 1.445 2.87 1.555 ;
      RECT  2.14 0.34 2.35 0.46 ;
      RECT  2.14 0.46 2.23 1.045 ;
      RECT  1.595 1.045 2.23 1.155 ;
      RECT  0.79 0.45 1.815 0.55 ;
      RECT  0.79 0.55 0.88 0.755 ;
      RECT  1.35 0.55 1.45 1.245 ;
      RECT  0.525 0.755 0.88 0.925 ;
      RECT  0.79 0.925 0.88 1.245 ;
      RECT  0.79 1.245 1.02 1.355 ;
      RECT  1.35 1.245 2.34 1.355 ;
      RECT  2.57 0.51 2.67 0.575 ;
      RECT  2.57 0.575 2.87 0.69 ;
      RECT  2.78 0.69 2.87 1.04 ;
      RECT  2.655 1.04 2.87 1.16 ;
      RECT  1.95 0.51 2.05 0.775 ;
      RECT  1.6 0.775 2.05 0.895 ;
      RECT  0.335 0.29 0.435 1.23 ;
      LAYER M2 ;
      RECT  0.295 0.35 2.32 0.45 ;
      RECT  1.91 0.55 2.71 0.65 ;
      LAYER V1 ;
      RECT  0.335 0.35 0.435 0.45 ;
      RECT  2.18 0.35 2.28 0.45 ;
      RECT  1.95 0.55 2.05 0.65 ;
      RECT  2.57 0.55 2.67 0.65 ;
  END
END SEN_EO2_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EO2_G_8
#      Description : "2-Input exclusive OR"
#      Equation    : X=A1^A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO2_G_8
  CLASS CORE ;
  FOREIGN SEN_EO2_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.705 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.45 0.925 ;
      RECT  4.35 0.925 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.18 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  0.58 1.45 0.71 1.75 ;
      RECT  1.105 1.21 1.225 1.75 ;
      RECT  1.62 1.45 1.75 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  4.74 1.455 4.865 1.75 ;
      RECT  5.255 1.455 5.385 1.75 ;
      RECT  5.775 1.41 5.905 1.75 ;
      RECT  6.295 1.41 6.425 1.75 ;
      RECT  6.815 1.41 6.945 1.75 ;
      RECT  7.36 1.21 7.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  0.58 0.05 0.71 0.35 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.155 0.05 2.285 0.36 ;
      RECT  5.775 0.05 5.905 0.39 ;
      RECT  6.295 0.05 6.425 0.39 ;
      RECT  6.815 0.05 6.945 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.105 0.05 1.225 0.59 ;
      RECT  4.74 0.05 4.86 0.59 ;
      RECT  5.26 0.05 5.38 0.59 ;
      RECT  7.36 0.05 7.48 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.52 0.51 7.25 0.69 ;
      RECT  6.68 0.69 6.85 1.11 ;
      RECT  5.52 1.11 7.25 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.56 0.445 3.3 0.555 ;
      RECT  3.19 0.555 3.3 0.635 ;
      RECT  2.56 0.555 2.66 1.09 ;
      RECT  3.58 0.445 4.4 0.555 ;
      RECT  3.58 0.555 3.67 1.055 ;
      RECT  3.35 1.055 3.67 1.145 ;
      RECT  3.35 1.145 3.45 1.24 ;
      RECT  1.315 0.45 2.43 0.57 ;
      RECT  2.34 0.57 2.43 1.24 ;
      RECT  1.315 1.24 3.45 1.35 ;
      RECT  0.275 0.44 0.99 0.56 ;
      RECT  0.89 0.56 0.99 0.78 ;
      RECT  0.89 0.78 2.16 0.89 ;
      RECT  2.06 0.89 2.16 1.09 ;
      RECT  0.89 0.89 0.99 1.24 ;
      RECT  0.275 1.24 0.99 1.36 ;
      RECT  4.975 0.505 5.17 0.625 ;
      RECT  4.975 0.625 5.075 1.0 ;
      RECT  4.975 1.0 5.145 1.105 ;
      RECT  3.39 0.51 3.49 0.725 ;
      RECT  2.95 0.725 3.49 0.905 ;
      RECT  5.235 0.78 6.57 0.95 ;
      RECT  5.235 0.95 5.405 1.195 ;
      RECT  2.375 0.24 4.65 0.355 ;
      RECT  4.55 0.355 4.65 1.195 ;
      RECT  4.55 1.195 5.405 1.365 ;
      RECT  4.55 1.365 4.65 1.445 ;
      RECT  2.36 1.445 4.65 1.555 ;
      RECT  3.76 0.91 3.86 1.245 ;
      RECT  3.655 1.245 4.4 1.355 ;
      LAYER M2 ;
      RECT  3.35 0.55 5.115 0.65 ;
      RECT  2.02 0.95 3.9 1.05 ;
      LAYER V1 ;
      RECT  3.39 0.55 3.49 0.65 ;
      RECT  4.975 0.55 5.075 0.65 ;
      RECT  2.06 0.95 2.16 1.05 ;
      RECT  2.56 0.95 2.66 1.05 ;
      RECT  3.76 0.95 3.86 1.05 ;
  END
END SEN_EO2_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_3
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_3
  CLASS CORE ;
  FOREIGN SEN_EO3_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.65 0.89 ;
      RECT  7.15 0.89 7.25 0.945 ;
      RECT  7.55 0.89 7.65 1.09 ;
      RECT  6.75 0.945 7.25 1.045 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2061 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.665 2.25 0.91 ;
      RECT  2.15 0.91 2.45 0.945 ;
      RECT  2.15 0.945 3.09 1.09 ;
      RECT  4.26 0.715 5.165 0.85 ;
      LAYER M2 ;
      RECT  4.26 0.75 4.545 0.85 ;
      RECT  4.26 0.85 4.36 0.95 ;
      RECT  2.8 0.95 4.36 1.05 ;
      LAYER V1 ;
      RECT  2.84 0.95 2.94 1.05 ;
      RECT  4.405 0.75 4.505 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.393 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.095 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.42 0.45 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  1.36 1.415 1.49 1.75 ;
      RECT  5.245 1.415 5.37 1.75 ;
      RECT  5.765 1.21 5.885 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  1.36 0.05 1.49 0.35 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  5.24 0.05 5.37 0.36 ;
      RECT  0.845 0.05 0.965 0.59 ;
      RECT  5.765 0.05 5.885 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.545 0.375 6.665 0.47 ;
      RECT  6.545 0.47 7.85 0.59 ;
      RECT  7.75 0.59 7.85 1.315 ;
      RECT  6.49 1.315 7.85 1.405 ;
    END
    ANTENNADIFFAREA 0.55 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.665 0.17 3.295 0.26 ;
      RECT  2.665 0.26 2.785 0.35 ;
      RECT  3.185 0.26 3.295 1.14 ;
      RECT  3.185 1.14 3.4 1.18 ;
      RECT  2.72 1.18 3.4 1.285 ;
      RECT  3.295 1.285 3.4 1.33 ;
      RECT  6.3 0.175 6.925 0.265 ;
      RECT  6.3 0.265 6.45 0.37 ;
      RECT  6.805 0.265 6.925 0.38 ;
      RECT  6.35 0.37 6.45 1.035 ;
      RECT  6.265 1.035 6.45 1.125 ;
      RECT  6.265 1.125 6.375 1.495 ;
      RECT  6.265 1.495 6.945 1.6 ;
      RECT  3.385 0.23 4.06 0.35 ;
      RECT  3.385 0.35 3.49 0.83 ;
      RECT  3.385 0.83 3.6 0.945 ;
      RECT  3.49 0.945 3.6 1.45 ;
      RECT  3.49 1.45 4.17 1.56 ;
      RECT  3.49 1.56 3.6 1.57 ;
      RECT  1.625 0.23 2.315 0.35 ;
      RECT  1.625 0.35 1.745 0.44 ;
      RECT  1.055 0.44 1.745 0.56 ;
      RECT  1.625 0.56 1.745 1.205 ;
      RECT  0.275 0.785 0.935 0.895 ;
      RECT  0.845 0.895 0.935 1.205 ;
      RECT  0.845 1.205 1.745 1.325 ;
      RECT  1.625 1.325 1.745 1.465 ;
      RECT  1.625 1.465 2.29 1.555 ;
      RECT  2.12 1.555 2.29 1.57 ;
      RECT  2.12 1.57 3.6 1.66 ;
      RECT  4.355 0.23 5.05 0.35 ;
      RECT  4.93 0.35 5.05 0.45 ;
      RECT  4.93 0.45 5.405 0.57 ;
      RECT  5.285 0.57 5.405 0.945 ;
      RECT  5.04 0.945 5.405 1.065 ;
      RECT  5.04 1.065 5.155 1.45 ;
      RECT  4.475 1.45 5.155 1.57 ;
      RECT  7.315 0.23 8.05 0.35 ;
      RECT  7.94 0.35 8.05 1.495 ;
      RECT  7.375 1.495 8.05 1.6 ;
      RECT  2.915 0.35 3.095 0.44 ;
      RECT  1.885 0.44 3.095 0.56 ;
      RECT  1.885 0.56 2.005 1.255 ;
      RECT  1.885 1.255 2.59 1.375 ;
      RECT  2.47 1.375 3.205 1.48 ;
      RECT  3.58 0.44 4.815 0.56 ;
      RECT  3.74 0.56 3.86 1.24 ;
      RECT  3.74 1.24 4.95 1.36 ;
      RECT  4.285 1.36 4.385 1.51 ;
      RECT  0.065 0.45 0.745 0.565 ;
      RECT  0.565 0.565 0.745 0.65 ;
      RECT  0.065 0.565 0.185 1.21 ;
      RECT  0.065 1.21 0.755 1.33 ;
      RECT  6.055 0.17 6.175 0.565 ;
      RECT  6.055 0.565 6.26 0.735 ;
      RECT  6.055 0.735 6.175 1.13 ;
      RECT  6.025 1.13 6.175 1.315 ;
      RECT  6.54 0.705 6.985 0.815 ;
      RECT  6.54 0.815 6.63 1.135 ;
      RECT  6.54 1.135 7.46 1.225 ;
      RECT  7.36 0.99 7.46 1.135 ;
      RECT  2.525 0.705 3.095 0.85 ;
      RECT  3.97 0.675 4.08 0.945 ;
      RECT  3.97 0.945 4.84 1.055 ;
      RECT  5.505 0.31 5.625 1.38 ;
      LAYER M2 ;
      RECT  2.915 0.35 6.49 0.45 ;
      RECT  0.565 0.55 5.43 0.65 ;
      RECT  2.91 0.75 4.115 0.85 ;
      RECT  4.66 0.95 5.645 1.05 ;
      RECT  4.245 1.35 8.085 1.45 ;
      LAYER V1 ;
      RECT  2.955 0.35 3.055 0.45 ;
      RECT  6.35 0.35 6.45 0.45 ;
      RECT  0.605 0.55 0.705 0.65 ;
      RECT  3.195 0.55 3.295 0.65 ;
      RECT  5.29 0.55 5.39 0.65 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  3.975 0.75 4.075 0.85 ;
      RECT  4.7 0.95 4.8 1.05 ;
      RECT  5.505 0.95 5.605 1.05 ;
      RECT  4.285 1.35 4.385 1.45 ;
      RECT  7.945 1.35 8.045 1.45 ;
  END
END SEN_EO3_3
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_6
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_6
  CLASS CORE ;
  FOREIGN SEN_EO3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.95 0.51 12.05 0.71 ;
      RECT  10.51 0.71 12.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3834 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 0.71 9.12 0.92 ;
      RECT  8.55 0.92 8.65 1.09 ;
      RECT  4.915 0.71 5.26 0.79 ;
      RECT  4.175 0.79 5.26 0.89 ;
      RECT  5.16 0.89 5.26 1.105 ;
      LAYER M2 ;
      RECT  5.12 0.95 8.69 1.05 ;
      LAYER V1 ;
      RECT  8.55 0.95 8.65 1.05 ;
      RECT  5.16 0.95 5.26 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7311 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.25 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 13.6 1.85 ;
      RECT  0.58 1.415 0.71 1.75 ;
      RECT  1.1 1.415 1.23 1.75 ;
      RECT  1.62 1.415 1.75 1.75 ;
      RECT  2.14 1.415 2.27 1.75 ;
      RECT  2.66 1.415 2.79 1.75 ;
      RECT  3.185 1.21 3.305 1.75 ;
      RECT  3.7 1.41 3.83 1.75 ;
      RECT  9.805 1.515 9.935 1.75 ;
      RECT  10.425 1.515 10.55 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 13.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
      RECT  11.85 1.75 11.95 1.85 ;
      RECT  12.45 1.75 12.55 1.85 ;
      RECT  13.05 1.75 13.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 13.6 0.05 ;
      RECT  9.885 0.05 10.015 0.29 ;
      RECT  10.425 0.05 10.555 0.29 ;
      RECT  3.7 0.05 3.83 0.35 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.1 0.05 1.23 0.385 ;
      RECT  1.62 0.05 1.75 0.385 ;
      RECT  2.14 0.05 2.27 0.385 ;
      RECT  2.66 0.05 2.79 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.185 0.05 3.305 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 13.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
      RECT  11.85 -0.05 11.95 0.05 ;
      RECT  12.45 -0.05 12.55 0.05 ;
      RECT  13.05 -0.05 13.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.87 0.23 12.26 0.35 ;
      RECT  12.14 0.35 12.26 0.54 ;
      RECT  12.14 0.54 13.3 0.655 ;
      RECT  13.15 0.655 13.3 1.34 ;
      RECT  10.885 1.34 13.3 1.455 ;
    END
    ANTENNADIFFAREA 1.027 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.795 0.33 8.245 0.35 ;
      RECT  6.795 0.35 9.34 0.45 ;
      RECT  8.125 0.45 9.34 0.47 ;
      RECT  6.795 0.45 6.91 0.5 ;
      RECT  9.235 0.47 9.34 0.56 ;
      RECT  5.73 0.5 6.91 0.62 ;
      RECT  9.235 0.56 9.85 0.68 ;
      RECT  6.795 0.62 6.91 1.215 ;
      RECT  4.69 1.215 8.25 1.335 ;
      RECT  4.42 0.24 6.705 0.36 ;
      RECT  4.42 0.36 4.6 0.45 ;
      RECT  12.35 0.33 13.535 0.45 ;
      RECT  13.415 0.45 13.535 1.545 ;
      RECT  10.615 1.35 10.795 1.45 ;
      RECT  10.69 1.45 10.795 1.545 ;
      RECT  10.69 1.545 13.535 1.66 ;
      RECT  3.395 0.44 4.085 0.56 ;
      RECT  3.965 0.56 4.085 1.14 ;
      RECT  3.395 1.14 4.085 1.26 ;
      RECT  7.0 0.54 8.04 0.56 ;
      RECT  7.0 0.56 8.45 0.66 ;
      RECT  7.895 0.66 8.45 0.68 ;
      RECT  8.35 0.68 8.45 1.215 ;
      RECT  8.35 1.215 9.33 1.335 ;
      RECT  4.195 0.46 4.315 0.575 ;
      RECT  4.195 0.575 5.45 0.595 ;
      RECT  4.69 0.475 5.45 0.575 ;
      RECT  4.195 0.595 4.79 0.665 ;
      RECT  5.35 0.595 5.45 1.0 ;
      RECT  5.35 1.0 6.42 1.12 ;
      RECT  0.275 0.475 1.75 0.595 ;
      RECT  1.65 0.595 1.75 0.78 ;
      RECT  1.65 0.78 2.855 0.9 ;
      RECT  1.65 0.9 1.75 1.195 ;
      RECT  0.275 1.195 1.75 1.315 ;
      RECT  1.84 0.475 3.095 0.595 ;
      RECT  2.995 0.595 3.095 1.195 ;
      RECT  1.84 1.195 3.095 1.315 ;
      RECT  5.54 0.49 5.64 0.75 ;
      RECT  5.54 0.75 6.695 0.895 ;
      RECT  7.105 0.75 7.795 0.79 ;
      RECT  7.105 0.79 8.14 0.895 ;
      RECT  12.22 0.775 13.04 0.895 ;
      RECT  12.22 0.895 12.32 0.98 ;
      RECT  10.135 0.56 10.335 0.68 ;
      RECT  10.135 0.68 10.235 0.98 ;
      RECT  10.135 0.98 12.32 1.07 ;
      RECT  10.135 1.07 10.28 1.245 ;
      RECT  10.405 1.16 12.97 1.25 ;
      RECT  10.405 1.25 10.495 1.335 ;
      RECT  7.24 0.14 9.565 0.24 ;
      RECT  8.345 0.24 9.565 0.26 ;
      RECT  9.445 0.26 9.565 0.38 ;
      RECT  9.445 0.38 10.555 0.44 ;
      RECT  9.445 0.44 11.86 0.47 ;
      RECT  10.455 0.47 11.86 0.56 ;
      RECT  9.94 0.47 10.045 1.26 ;
      RECT  9.445 1.26 10.045 1.335 ;
      RECT  9.445 1.335 10.495 1.425 ;
      RECT  9.445 1.425 9.565 1.44 ;
      RECT  7.25 1.44 9.565 1.56 ;
      RECT  4.415 1.29 4.525 1.425 ;
      RECT  4.415 1.425 6.71 1.545 ;
      LAYER M2 ;
      RECT  4.42 0.35 12.53 0.45 ;
      RECT  3.935 0.55 5.68 0.65 ;
      RECT  5.78 0.55 7.645 0.65 ;
      RECT  5.78 0.65 5.88 0.75 ;
      RECT  1.61 0.75 5.88 0.85 ;
      RECT  6.245 0.75 7.46 0.85 ;
      RECT  2.955 1.15 6.935 1.25 ;
      RECT  4.38 1.35 10.795 1.45 ;
      LAYER V1 ;
      RECT  4.46 0.35 4.56 0.45 ;
      RECT  12.39 0.35 12.49 0.45 ;
      RECT  3.975 0.55 4.075 0.65 ;
      RECT  5.54 0.55 5.64 0.65 ;
      RECT  7.14 0.55 7.24 0.65 ;
      RECT  7.505 0.55 7.605 0.65 ;
      RECT  1.65 0.75 1.75 0.85 ;
      RECT  5.35 0.75 5.45 0.85 ;
      RECT  6.285 0.75 6.385 0.85 ;
      RECT  6.555 0.75 6.655 0.85 ;
      RECT  7.32 0.75 7.42 0.85 ;
      RECT  2.995 1.15 3.095 1.25 ;
      RECT  6.795 1.15 6.895 1.25 ;
      RECT  4.42 1.35 4.52 1.45 ;
      RECT  10.655 1.35 10.755 1.45 ;
  END
END SEN_EO3_6
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_1
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_1
  CLASS CORE ;
  FOREIGN SEN_EO3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 2.68 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0732 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.34 0.51 2.45 1.07 ;
      RECT  2.315 1.07 2.45 1.31 ;
      RECT  1.455 0.865 1.555 1.35 ;
      RECT  0.815 0.925 0.925 1.17 ;
      RECT  0.815 1.17 0.915 1.4 ;
      LAYER M2 ;
      RECT  0.71 1.15 2.49 1.25 ;
      LAYER V1 ;
      RECT  2.315 1.15 2.415 1.25 ;
      RECT  1.455 1.15 1.555 1.25 ;
      RECT  0.815 1.15 0.915 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1119 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.67 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.59 0.485 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  2.39 1.58 2.6 1.75 ;
      RECT  3.725 1.255 3.855 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.335 0.05 0.465 0.38 ;
      RECT  2.455 0.05 2.585 0.4 ;
      RECT  3.745 0.05 3.86 0.5 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.3 4.13 0.6 ;
      RECT  3.95 0.6 4.05 1.2 ;
      RECT  3.95 1.2 4.13 1.5 ;
    END
    ANTENNADIFFAREA 0.185 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.625 0.14 1.935 0.23 ;
      RECT  1.845 0.23 1.935 0.46 ;
      RECT  0.625 0.23 0.725 1.3 ;
      RECT  1.845 0.46 2.055 0.675 ;
      RECT  1.845 0.675 1.935 1.24 ;
      RECT  1.845 1.24 1.995 1.48 ;
      RECT  2.695 0.24 2.875 0.36 ;
      RECT  2.77 0.36 2.875 0.77 ;
      RECT  2.77 0.77 2.935 0.97 ;
      RECT  2.77 0.97 2.87 1.2 ;
      RECT  2.65 1.2 2.87 1.31 ;
      RECT  2.155 0.26 2.365 0.38 ;
      RECT  2.155 0.38 2.25 0.765 ;
      RECT  2.085 0.765 2.25 0.985 ;
      RECT  2.085 0.985 2.225 1.26 ;
      RECT  0.825 0.34 1.47 0.45 ;
      RECT  0.825 0.45 1.165 0.46 ;
      RECT  1.075 0.46 1.165 1.25 ;
      RECT  1.005 1.25 1.165 1.445 ;
      RECT  3.18 0.33 3.62 0.45 ;
      RECT  3.5 0.45 3.62 0.59 ;
      RECT  3.5 0.59 3.86 0.69 ;
      RECT  3.77 0.69 3.86 1.075 ;
      RECT  3.54 1.075 3.86 1.165 ;
      RECT  3.54 1.165 3.63 1.425 ;
      RECT  3.405 1.425 3.63 1.545 ;
      RECT  2.98 0.41 3.085 0.54 ;
      RECT  2.98 0.54 3.115 0.64 ;
      RECT  3.025 0.64 3.115 1.4 ;
      RECT  2.11 1.4 3.115 1.49 ;
      RECT  2.11 1.49 2.2 1.57 ;
      RECT  1.645 0.42 1.735 1.57 ;
      RECT  1.645 1.57 2.2 1.66 ;
      RECT  1.255 0.54 1.46 0.65 ;
      RECT  1.255 0.65 1.365 1.555 ;
      RECT  0.065 0.3 0.185 0.47 ;
      RECT  0.065 0.47 0.535 0.56 ;
      RECT  0.445 0.56 0.535 1.41 ;
      RECT  0.065 1.41 0.69 1.5 ;
      RECT  0.6 1.5 0.69 1.555 ;
      RECT  0.065 1.5 0.185 1.62 ;
      RECT  0.6 1.555 1.365 1.645 ;
      RECT  3.205 0.54 3.385 0.78 ;
      RECT  3.205 0.78 3.68 0.87 ;
      RECT  3.52 0.87 3.68 0.985 ;
      RECT  3.205 0.87 3.3 1.48 ;
      LAYER M2 ;
      RECT  1.02 0.35 3.59 0.45 ;
      LAYER V1 ;
      RECT  1.095 0.35 1.195 0.45 ;
      RECT  1.295 0.35 1.395 0.45 ;
      RECT  3.22 0.35 3.32 0.45 ;
      RECT  3.42 0.35 3.52 0.45 ;
  END
END SEN_EO3_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_2
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_2
  CLASS CORE ;
  FOREIGN SEN_EO3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.64 0.5 5.78 0.75 ;
      RECT  5.64 0.75 6.06 0.925 ;
      RECT  4.71 0.68 4.885 1.1 ;
      LAYER M2 ;
      RECT  4.71 0.75 6.06 0.85 ;
      LAYER V1 ;
      RECT  5.68 0.75 5.78 0.85 ;
      RECT  5.88 0.75 5.98 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1464 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.445 0.68 4.6 1.145 ;
      RECT  2.98 0.68 3.08 1.185 ;
      RECT  2.21 0.7 2.59 0.9 ;
      RECT  1.35 0.7 1.85 0.9 ;
      RECT  1.35 0.9 1.62 0.985 ;
      LAYER M2 ;
      RECT  1.46 0.75 4.59 0.85 ;
      LAYER V1 ;
      RECT  4.445 0.75 4.545 0.85 ;
      RECT  2.98 0.75 3.08 0.85 ;
      RECT  2.25 0.75 2.35 0.85 ;
      RECT  2.45 0.75 2.55 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2238 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.09 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  0.565 1.615 0.745 1.75 ;
      RECT  1.11 1.615 1.29 1.75 ;
      RECT  3.985 1.615 4.19 1.75 ;
      RECT  4.565 1.615 4.745 1.75 ;
      RECT  5.105 1.615 5.285 1.75 ;
      RECT  6.68 1.2 6.8 1.75 ;
      RECT  7.2 1.21 7.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  1.105 0.05 1.295 0.21 ;
      RECT  0.065 0.05 0.185 0.39 ;
      RECT  0.58 0.05 0.71 0.4 ;
      RECT  6.37 0.05 6.5 0.41 ;
      RECT  6.65 0.05 6.78 0.41 ;
      RECT  4.46 0.05 4.58 0.59 ;
      RECT  7.2 0.05 7.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.5 7.05 1.3 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.68 0.14 3.795 0.23 ;
      RECT  1.68 0.23 1.8 0.3 ;
      RECT  3.625 0.23 3.795 0.51 ;
      RECT  0.81 0.3 1.8 0.39 ;
      RECT  0.81 0.39 1.24 0.41 ;
      RECT  1.15 0.41 1.24 1.075 ;
      RECT  3.625 0.51 3.715 1.27 ;
      RECT  0.87 1.075 1.83 1.165 ;
      RECT  0.87 1.165 0.99 1.325 ;
      RECT  3.45 1.27 3.715 1.37 ;
      RECT  1.965 0.32 2.765 0.41 ;
      RECT  1.965 0.41 2.065 0.5 ;
      RECT  1.365 0.5 2.065 0.59 ;
      RECT  1.965 0.59 2.065 1.13 ;
      RECT  1.965 1.13 2.61 1.22 ;
      RECT  1.965 1.22 2.065 1.255 ;
      RECT  1.34 1.255 2.065 1.345 ;
      RECT  4.72 0.37 4.84 0.5 ;
      RECT  4.72 0.5 5.065 0.59 ;
      RECT  4.975 0.59 5.065 0.75 ;
      RECT  4.975 0.75 5.19 0.95 ;
      RECT  4.975 0.95 5.065 1.235 ;
      RECT  4.81 1.235 5.065 1.325 ;
      RECT  5.205 0.335 5.37 0.505 ;
      RECT  5.28 0.505 5.37 1.28 ;
      RECT  5.16 1.28 5.835 1.37 ;
      RECT  5.16 1.37 5.25 1.415 ;
      RECT  3.95 0.37 4.07 0.6 ;
      RECT  3.805 0.6 4.07 0.69 ;
      RECT  3.805 0.69 3.895 1.415 ;
      RECT  3.805 1.415 5.25 1.48 ;
      RECT  2.875 0.32 3.535 0.41 ;
      RECT  3.425 0.41 3.535 0.7 ;
      RECT  3.24 0.7 3.535 0.79 ;
      RECT  3.24 0.79 3.34 1.48 ;
      RECT  3.24 1.48 5.25 1.49 ;
      RECT  2.665 1.49 5.25 1.505 ;
      RECT  2.665 1.505 3.895 1.58 ;
      RECT  5.87 0.335 5.975 0.55 ;
      RECT  5.87 0.55 6.85 0.65 ;
      RECT  6.76 0.65 6.85 1.02 ;
      RECT  6.465 1.02 6.85 1.11 ;
      RECT  6.465 1.11 6.555 1.28 ;
      RECT  6.105 1.28 6.555 1.37 ;
      RECT  2.305 0.5 3.315 0.59 ;
      RECT  2.78 0.59 2.87 1.3 ;
      RECT  2.78 1.3 3.13 1.31 ;
      RECT  2.17 1.31 3.13 1.4 ;
      RECT  2.17 1.4 2.29 1.435 ;
      RECT  0.325 0.3 0.445 0.5 ;
      RECT  0.325 0.5 0.755 0.59 ;
      RECT  0.665 0.59 0.755 0.79 ;
      RECT  0.665 0.79 1.06 0.89 ;
      RECT  0.665 0.89 0.755 1.435 ;
      RECT  0.325 1.3 0.445 1.435 ;
      RECT  0.325 1.435 2.29 1.525 ;
      RECT  4.2 0.43 4.32 0.8 ;
      RECT  4.005 0.8 4.32 0.89 ;
      RECT  4.005 0.89 4.095 1.235 ;
      RECT  4.005 1.235 4.5 1.325 ;
      RECT  6.21 0.81 6.67 0.91 ;
      RECT  6.21 0.91 6.3 1.08 ;
      RECT  4.97 0.155 6.23 0.245 ;
      RECT  5.46 0.245 5.6 0.4 ;
      RECT  4.97 0.245 5.09 0.41 ;
      RECT  6.115 0.245 6.23 0.42 ;
      RECT  5.46 0.4 5.55 1.08 ;
      RECT  5.46 1.08 6.3 1.17 ;
      RECT  5.925 1.17 6.015 1.48 ;
      RECT  5.365 1.48 6.59 1.57 ;
      LAYER M2 ;
      RECT  1.87 0.55 6.47 0.65 ;
      LAYER V1 ;
      RECT  1.965 0.55 2.065 0.65 ;
      RECT  6.08 0.55 6.18 0.65 ;
      RECT  6.28 0.55 6.38 0.65 ;
  END
END SEN_EO3_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_4
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_4
  CLASS CORE ;
  FOREIGN SEN_EO3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.92 7.26 1.06 ;
      LAYER M2 ;
      RECT  6.5 0.95 7.3 1.05 ;
      LAYER V1 ;
      RECT  6.75 0.95 6.85 1.05 ;
      RECT  6.95 0.95 7.05 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2928 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.25 0.635 5.35 1.07 ;
      RECT  3.15 0.7 3.6 0.915 ;
      RECT  2.98 0.915 3.6 0.93 ;
      RECT  2.98 0.93 3.25 1.05 ;
      RECT  1.55 0.7 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.1 ;
      LAYER M2 ;
      RECT  1.5 0.75 5.5 0.85 ;
      LAYER V1 ;
      RECT  5.25 0.75 5.35 0.85 ;
      RECT  3.23 0.75 3.33 0.85 ;
      RECT  3.43 0.75 3.53 0.85 ;
      RECT  1.7 0.75 1.8 0.85 ;
      RECT  1.9 0.75 2.0 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4476 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.36 1.435 1.49 1.75 ;
      RECT  5.215 1.6 5.395 1.75 ;
      RECT  5.755 1.6 5.935 1.75 ;
      RECT  6.31 1.43 6.44 1.75 ;
      RECT  8.575 1.21 8.695 1.75 ;
      RECT  9.09 1.41 9.22 1.75 ;
      RECT  9.615 1.21 9.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  5.21 0.05 5.39 0.185 ;
      RECT  5.91 0.05 6.09 0.185 ;
      RECT  6.525 0.05 6.705 0.185 ;
      RECT  8.545 0.05 8.725 0.305 ;
      RECT  0.32 0.05 0.445 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      RECT  9.09 0.05 9.22 0.39 ;
      RECT  9.615 0.05 9.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.85 0.51 9.46 0.69 ;
      RECT  9.35 0.69 9.46 1.11 ;
      RECT  8.85 1.11 9.46 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.18 0.16 5.105 0.23 ;
      RECT  2.0 0.23 5.105 0.25 ;
      RECT  5.015 0.25 5.105 0.275 ;
      RECT  2.0 0.25 3.285 0.33 ;
      RECT  5.015 0.275 6.895 0.36 ;
      RECT  2.605 0.33 2.695 0.7 ;
      RECT  5.015 0.36 7.995 0.365 ;
      RECT  6.805 0.365 7.995 0.46 ;
      RECT  7.885 0.46 7.995 0.575 ;
      RECT  7.885 0.575 8.54 0.665 ;
      RECT  7.975 0.665 8.065 1.11 ;
      RECT  2.15 0.7 2.695 0.79 ;
      RECT  2.15 0.79 2.25 1.21 ;
      RECT  7.35 1.11 8.065 1.15 ;
      RECT  6.78 1.15 8.065 1.2 ;
      RECT  6.78 1.2 7.475 1.25 ;
      RECT  1.835 1.21 3.085 1.31 ;
      RECT  6.78 1.25 6.905 1.365 ;
      RECT  6.985 0.16 8.205 0.25 ;
      RECT  8.085 0.25 8.205 0.395 ;
      RECT  8.085 0.395 8.74 0.485 ;
      RECT  8.65 0.485 8.74 0.79 ;
      RECT  8.155 0.79 9.24 0.89 ;
      RECT  8.155 0.89 8.255 1.31 ;
      RECT  7.58 1.31 8.255 1.4 ;
      RECT  7.58 1.4 7.685 1.44 ;
      RECT  6.99 1.44 7.685 1.54 ;
      RECT  3.605 0.34 4.905 0.43 ;
      RECT  4.815 0.43 4.905 0.455 ;
      RECT  4.815 0.455 6.69 0.545 ;
      RECT  6.6 0.545 6.69 0.56 ;
      RECT  5.75 0.545 5.85 1.35 ;
      RECT  6.6 0.56 7.47 0.65 ;
      RECT  5.47 1.35 5.85 1.4 ;
      RECT  4.485 1.4 5.85 1.47 ;
      RECT  3.405 1.47 5.85 1.49 ;
      RECT  3.405 1.49 4.66 1.57 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 0.92 0.59 ;
      RECT  0.82 0.59 0.92 0.78 ;
      RECT  0.82 0.78 1.24 0.9 ;
      RECT  0.82 0.9 0.92 1.21 ;
      RECT  0.065 1.21 0.92 1.31 ;
      RECT  0.065 1.31 0.185 1.43 ;
      RECT  2.805 0.44 3.495 0.52 ;
      RECT  2.805 0.52 4.08 0.53 ;
      RECT  3.34 0.53 4.08 0.61 ;
      RECT  3.72 0.61 4.08 0.63 ;
      RECT  3.72 0.63 3.81 1.11 ;
      RECT  3.34 1.11 3.81 1.195 ;
      RECT  3.195 1.195 3.81 1.29 ;
      RECT  3.195 1.29 3.295 1.43 ;
      RECT  2.61 1.43 3.295 1.53 ;
      RECT  1.05 0.49 2.495 0.59 ;
      RECT  1.35 0.59 1.44 1.21 ;
      RECT  1.11 1.21 1.44 1.22 ;
      RECT  1.11 1.22 1.735 1.31 ;
      RECT  1.635 1.31 1.735 1.45 ;
      RECT  1.11 1.31 1.22 1.51 ;
      RECT  1.635 1.45 2.32 1.55 ;
      RECT  4.37 0.54 4.705 0.63 ;
      RECT  4.615 0.63 4.705 0.635 ;
      RECT  4.615 0.635 5.14 0.725 ;
      RECT  4.615 0.725 4.705 1.125 ;
      RECT  4.615 1.125 4.85 1.14 ;
      RECT  4.1 1.14 4.85 1.26 ;
      RECT  4.745 1.26 4.85 1.31 ;
      RECT  6.22 0.635 6.45 0.73 ;
      RECT  6.36 0.73 6.45 0.74 ;
      RECT  6.36 0.74 7.825 0.83 ;
      RECT  7.72 0.83 7.825 0.99 ;
      RECT  6.36 0.83 6.45 1.21 ;
      RECT  6.0 1.21 6.69 1.31 ;
      RECT  6.575 1.31 6.69 1.62 ;
      RECT  5.46 0.635 5.66 0.735 ;
      RECT  5.56 0.735 5.66 1.16 ;
      RECT  4.94 0.88 5.05 1.16 ;
      RECT  4.94 1.16 5.66 1.26 ;
      RECT  3.905 0.74 4.525 0.84 ;
      RECT  3.905 0.84 4.01 1.14 ;
      RECT  2.785 0.62 2.88 0.9 ;
      RECT  2.345 0.9 2.88 1.07 ;
      RECT  8.345 1.27 8.455 1.49 ;
      RECT  7.775 1.49 8.455 1.59 ;
      LAYER M2 ;
      RECT  2.46 0.95 5.12 1.05 ;
      RECT  0.73 1.15 3.75 1.25 ;
      RECT  3.9 1.15 4.54 1.25 ;
      RECT  3.9 1.25 4.0 1.35 ;
      RECT  1.03 1.35 4.0 1.45 ;
      RECT  5.46 1.35 8.49 1.45 ;
      LAYER V1 ;
      RECT  2.53 0.95 2.63 1.05 ;
      RECT  2.73 0.95 2.83 1.05 ;
      RECT  3.91 0.95 4.01 1.05 ;
      RECT  4.945 0.95 5.045 1.05 ;
      RECT  0.82 1.15 0.92 1.25 ;
      RECT  3.35 1.15 3.45 1.25 ;
      RECT  3.55 1.15 3.65 1.25 ;
      RECT  4.14 1.15 4.24 1.25 ;
      RECT  4.34 1.15 4.44 1.25 ;
      RECT  1.115 1.35 1.215 1.45 ;
      RECT  5.55 1.35 5.65 1.45 ;
      RECT  5.75 1.35 5.85 1.45 ;
      RECT  8.35 1.35 8.45 1.45 ;
  END
END SEN_EO3_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_DG_1
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_DG_1
  CLASS CORE ;
  FOREIGN SEN_EO3_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 3.85 0.69 ;
      RECT  3.55 0.69 3.65 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0492 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.67 2.85 0.73 ;
      RECT  2.645 0.73 2.85 0.9 ;
      RECT  2.75 0.9 2.85 1.09 ;
      RECT  1.15 0.67 1.25 1.09 ;
      LAYER M2 ;
      RECT  1.11 0.75 2.85 0.85 ;
      LAYER V1 ;
      RECT  2.71 0.75 2.81 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.69 0.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.415 0.45 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.85 1.415 0.97 1.75 ;
      RECT  2.94 1.585 3.06 1.75 ;
      RECT  4.255 1.585 4.375 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  2.94 0.05 3.06 0.215 ;
      RECT  4.245 0.05 4.375 0.215 ;
      RECT  0.33 0.05 0.45 0.385 ;
      RECT  0.85 0.05 0.97 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.47 4.675 1.29 ;
    END
    ANTENNADIFFAREA 0.175 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.96 0.14 2.835 0.205 ;
      RECT  1.865 0.205 2.835 0.23 ;
      RECT  1.865 0.23 2.07 0.345 ;
      RECT  1.98 0.345 2.07 0.69 ;
      RECT  1.98 0.69 2.275 0.78 ;
      RECT  2.155 0.78 2.275 1.17 ;
      RECT  2.145 1.17 2.275 1.26 ;
      RECT  2.16 1.26 2.275 1.51 ;
      RECT  3.73 0.215 3.85 0.31 ;
      RECT  3.73 0.31 4.285 0.4 ;
      RECT  4.195 0.4 4.285 0.785 ;
      RECT  4.195 0.785 4.455 0.895 ;
      RECT  4.195 0.895 4.285 1.35 ;
      RECT  3.705 1.35 4.285 1.455 ;
      RECT  1.57 0.2 1.775 0.32 ;
      RECT  1.57 0.32 1.66 0.785 ;
      RECT  1.57 0.785 1.7 0.875 ;
      RECT  1.61 0.875 1.7 1.31 ;
      RECT  1.61 1.31 1.785 1.61 ;
      RECT  2.97 0.305 3.615 0.32 ;
      RECT  2.39 0.32 3.615 0.41 ;
      RECT  2.97 0.41 3.615 0.42 ;
      RECT  2.97 0.42 3.06 1.39 ;
      RECT  2.76 1.39 3.06 1.395 ;
      RECT  2.76 1.395 3.285 1.405 ;
      RECT  2.39 1.405 3.285 1.495 ;
      RECT  3.195 1.495 3.285 1.545 ;
      RECT  3.195 1.545 4.145 1.66 ;
      RECT  0.565 0.245 0.745 0.365 ;
      RECT  0.645 0.365 0.745 1.44 ;
      RECT  0.565 1.44 0.745 1.56 ;
      RECT  0.07 0.245 0.19 0.48 ;
      RECT  0.07 0.48 0.545 0.6 ;
      RECT  0.445 0.6 0.545 1.205 ;
      RECT  0.07 1.205 0.545 1.325 ;
      RECT  0.07 1.325 0.235 1.49 ;
      RECT  1.11 0.215 1.23 0.49 ;
      RECT  0.905 0.49 1.23 0.58 ;
      RECT  0.905 0.58 1.005 1.2 ;
      RECT  0.905 1.2 1.23 1.29 ;
      RECT  1.11 1.29 1.23 1.6 ;
      RECT  2.16 0.32 2.275 0.5 ;
      RECT  2.16 0.5 2.485 0.59 ;
      RECT  2.385 0.59 2.485 1.195 ;
      RECT  2.385 1.195 2.855 1.3 ;
      RECT  1.79 0.435 1.89 0.855 ;
      RECT  1.365 0.41 1.48 0.95 ;
      RECT  1.34 0.95 1.52 1.05 ;
      RECT  3.22 0.51 3.34 0.99 ;
      RECT  3.22 0.99 3.915 1.08 ;
      RECT  3.815 0.78 3.915 0.99 ;
      RECT  3.22 1.08 3.34 1.26 ;
      RECT  4.005 0.49 4.105 1.17 ;
      RECT  3.47 1.17 4.105 1.26 ;
      RECT  3.47 1.26 3.59 1.35 ;
      RECT  3.4 1.35 3.59 1.45 ;
      RECT  1.34 1.15 1.48 1.605 ;
      RECT  1.875 0.945 2.055 1.61 ;
      LAYER M2 ;
      RECT  0.865 0.55 1.93 0.65 ;
      RECT  0.605 0.95 2.525 1.05 ;
      RECT  1.42 1.15 2.3 1.25 ;
      RECT  1.42 1.25 1.52 1.35 ;
      RECT  0.095 1.35 1.52 1.45 ;
      RECT  1.645 1.35 3.58 1.45 ;
      LAYER V1 ;
      RECT  0.905 0.55 1.005 0.65 ;
      RECT  1.79 0.55 1.89 0.65 ;
      RECT  0.645 0.95 0.745 1.05 ;
      RECT  1.38 0.95 1.48 1.05 ;
      RECT  1.915 0.95 2.015 1.05 ;
      RECT  2.385 0.95 2.485 1.05 ;
      RECT  2.16 1.15 2.26 1.25 ;
      RECT  0.135 1.35 0.235 1.45 ;
      RECT  1.38 1.35 1.48 1.45 ;
      RECT  1.685 1.35 1.785 1.45 ;
      RECT  3.44 1.35 3.54 1.45 ;
  END
END SEN_EO3_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_DG_2
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_DG_2
  CLASS CORE ;
  FOREIGN SEN_EO3_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 3.85 0.69 ;
      RECT  3.55 0.69 3.65 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.057 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.67 2.85 0.73 ;
      RECT  2.645 0.73 2.85 0.9 ;
      RECT  2.75 0.9 2.85 1.09 ;
      RECT  1.15 0.67 1.25 1.09 ;
      LAYER M2 ;
      RECT  1.11 0.75 2.85 0.85 ;
      LAYER V1 ;
      RECT  2.71 0.75 2.81 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0894 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.69 0.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.415 0.45 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.85 1.415 0.97 1.75 ;
      RECT  2.94 1.585 3.06 1.75 ;
      RECT  4.255 1.585 4.375 1.75 ;
      RECT  4.815 1.415 4.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  2.94 0.05 3.06 0.215 ;
      RECT  4.27 0.05 4.36 0.215 ;
      RECT  0.33 0.05 0.45 0.385 ;
      RECT  0.85 0.05 0.97 0.385 ;
      RECT  4.82 0.05 4.94 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.53 0.51 4.85 0.69 ;
      RECT  4.75 0.69 4.85 1.11 ;
      RECT  4.535 1.11 4.85 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.96 0.14 2.835 0.205 ;
      RECT  1.865 0.205 2.835 0.23 ;
      RECT  1.865 0.23 2.07 0.345 ;
      RECT  1.98 0.345 2.07 0.69 ;
      RECT  1.98 0.69 2.275 0.78 ;
      RECT  2.155 0.78 2.275 1.17 ;
      RECT  2.145 1.17 2.275 1.26 ;
      RECT  2.16 1.26 2.275 1.375 ;
      RECT  3.73 0.17 3.85 0.31 ;
      RECT  3.73 0.31 4.285 0.4 ;
      RECT  4.195 0.4 4.285 0.785 ;
      RECT  4.195 0.785 4.625 0.895 ;
      RECT  4.195 0.895 4.285 1.35 ;
      RECT  3.705 1.35 4.285 1.455 ;
      RECT  1.57 0.2 1.775 0.32 ;
      RECT  1.57 0.32 1.66 0.785 ;
      RECT  1.57 0.785 1.7 0.875 ;
      RECT  1.61 0.875 1.7 1.31 ;
      RECT  1.61 1.31 1.785 1.53 ;
      RECT  2.97 0.305 3.615 0.32 ;
      RECT  2.39 0.32 3.615 0.41 ;
      RECT  2.97 0.41 3.615 0.42 ;
      RECT  2.97 0.42 3.06 1.39 ;
      RECT  2.39 1.39 3.06 1.395 ;
      RECT  2.39 1.395 3.285 1.495 ;
      RECT  3.195 1.495 3.285 1.545 ;
      RECT  3.195 1.545 4.145 1.66 ;
      RECT  0.565 0.245 0.745 0.365 ;
      RECT  0.645 0.365 0.745 1.44 ;
      RECT  0.565 1.44 0.745 1.56 ;
      RECT  1.11 0.215 1.23 0.49 ;
      RECT  0.905 0.49 1.23 0.58 ;
      RECT  0.905 0.58 1.005 1.2 ;
      RECT  0.905 1.2 1.23 1.29 ;
      RECT  1.11 1.29 1.23 1.6 ;
      RECT  2.16 0.32 2.275 0.5 ;
      RECT  2.16 0.5 2.485 0.59 ;
      RECT  2.385 0.59 2.485 1.195 ;
      RECT  2.385 1.195 2.835 1.3 ;
      RECT  0.045 0.48 0.545 0.6 ;
      RECT  0.445 0.6 0.545 1.205 ;
      RECT  0.07 1.205 0.545 1.325 ;
      RECT  0.07 1.325 0.235 1.49 ;
      RECT  1.79 0.435 1.89 0.855 ;
      RECT  1.365 0.41 1.48 0.95 ;
      RECT  1.34 0.95 1.52 1.05 ;
      RECT  3.22 0.51 3.34 0.99 ;
      RECT  3.22 0.99 3.915 1.08 ;
      RECT  3.815 0.78 3.915 0.99 ;
      RECT  3.22 1.08 3.34 1.26 ;
      RECT  4.005 0.49 4.105 1.17 ;
      RECT  3.47 1.17 4.105 1.26 ;
      RECT  3.47 1.26 3.59 1.35 ;
      RECT  3.4 1.35 3.59 1.45 ;
      RECT  1.34 1.15 1.52 1.455 ;
      RECT  1.875 0.945 2.055 1.57 ;
      LAYER M2 ;
      RECT  0.865 0.55 1.93 0.65 ;
      RECT  0.605 0.95 2.525 1.05 ;
      RECT  1.42 1.15 2.3 1.25 ;
      RECT  1.42 1.25 1.52 1.35 ;
      RECT  0.095 1.35 1.52 1.45 ;
      RECT  1.645 1.35 3.58 1.45 ;
      LAYER V1 ;
      RECT  0.905 0.55 1.005 0.65 ;
      RECT  1.79 0.55 1.89 0.65 ;
      RECT  0.645 0.95 0.745 1.05 ;
      RECT  1.38 0.95 1.48 1.05 ;
      RECT  1.915 0.95 2.015 1.05 ;
      RECT  2.385 0.95 2.485 1.05 ;
      RECT  2.16 1.15 2.26 1.25 ;
      RECT  0.135 1.35 0.235 1.45 ;
      RECT  1.38 1.35 1.48 1.45 ;
      RECT  1.685 1.35 1.785 1.45 ;
      RECT  3.44 1.35 3.54 1.45 ;
  END
END SEN_EO3_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_DG_4
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_DG_4
  CLASS CORE ;
  FOREIGN SEN_EO3_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.6 0.51 4.045 0.68 ;
      RECT  3.6 0.68 3.69 0.89 ;
      LAYER M2 ;
      RECT  3.185 0.55 4.07 0.65 ;
      LAYER V1 ;
      RECT  3.67 0.55 3.77 0.65 ;
      RECT  3.87 0.55 3.97 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.755 0.71 3.055 0.9 ;
      RECT  1.34 0.67 1.44 1.09 ;
      LAYER M2 ;
      RECT  1.3 0.75 2.895 0.85 ;
      LAYER V1 ;
      RECT  2.755 0.75 2.855 0.85 ;
      RECT  1.34 0.75 1.44 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.36 1.31 4.53 1.4 ;
      RECT  4.435 1.4 4.53 1.75 ;
      RECT  0.055 1.415 0.175 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.575 1.415 0.695 1.75 ;
      RECT  1.07 1.45 1.24 1.75 ;
      RECT  3.115 1.585 3.235 1.75 ;
      RECT  4.905 1.415 5.025 1.75 ;
      RECT  5.42 1.44 5.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  3.12 0.05 3.235 0.215 ;
      RECT  4.345 0.05 4.465 0.215 ;
      RECT  0.575 0.05 0.695 0.345 ;
      RECT  0.055 0.05 0.175 0.36 ;
      RECT  1.095 0.05 1.215 0.365 ;
      RECT  5.42 0.05 5.545 0.365 ;
      RECT  4.905 0.05 5.025 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.62 0.51 5.45 0.69 ;
      RECT  5.35 0.69 5.45 1.11 ;
      RECT  4.625 1.11 5.45 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.13 0.14 3.03 0.205 ;
      RECT  2.035 0.205 3.03 0.23 ;
      RECT  2.035 0.23 2.24 0.335 ;
      RECT  2.15 0.335 2.24 0.71 ;
      RECT  2.15 0.71 2.445 0.8 ;
      RECT  2.325 0.8 2.445 1.35 ;
      RECT  3.6 0.23 3.77 0.305 ;
      RECT  3.17 0.305 3.77 0.32 ;
      RECT  2.56 0.32 3.77 0.42 ;
      RECT  2.56 0.42 3.28 0.44 ;
      RECT  3.17 0.44 3.28 1.375 ;
      RECT  2.56 1.375 3.28 1.395 ;
      RECT  2.56 1.395 3.44 1.495 ;
      RECT  3.35 1.495 3.44 1.545 ;
      RECT  3.35 1.545 4.33 1.66 ;
      RECT  1.745 0.2 1.945 0.32 ;
      RECT  1.745 0.32 1.845 1.35 ;
      RECT  1.745 1.35 1.985 1.45 ;
      RECT  3.86 0.305 4.475 0.42 ;
      RECT  4.385 0.42 4.475 0.785 ;
      RECT  4.385 0.785 4.985 0.895 ;
      RECT  4.385 0.895 4.475 1.13 ;
      RECT  4.14 1.13 4.475 1.22 ;
      RECT  4.14 1.22 4.23 1.365 ;
      RECT  3.86 1.365 4.23 1.455 ;
      RECT  1.355 0.19 1.46 0.49 ;
      RECT  1.15 0.49 1.46 0.58 ;
      RECT  1.15 0.58 1.25 1.2 ;
      RECT  1.15 1.2 1.46 1.29 ;
      RECT  1.355 1.29 1.46 1.61 ;
      RECT  2.33 0.33 2.445 0.53 ;
      RECT  2.33 0.53 2.655 0.62 ;
      RECT  2.555 0.62 2.655 1.165 ;
      RECT  2.555 1.165 2.99 1.285 ;
      RECT  0.29 0.435 0.71 0.555 ;
      RECT  0.62 0.555 0.71 0.755 ;
      RECT  0.62 0.755 0.845 0.925 ;
      RECT  0.62 0.925 0.72 1.205 ;
      RECT  0.315 1.205 0.72 1.325 ;
      RECT  0.315 1.325 0.445 1.49 ;
      RECT  0.81 0.435 1.035 0.555 ;
      RECT  0.935 0.555 1.035 1.22 ;
      RECT  0.84 1.22 1.035 1.35 ;
      RECT  0.84 1.35 0.96 1.44 ;
      RECT  4.17 0.51 4.295 0.68 ;
      RECT  4.195 0.68 4.295 0.95 ;
      RECT  3.96 0.95 4.295 1.04 ;
      RECT  3.96 1.04 4.05 1.185 ;
      RECT  3.64 1.185 4.05 1.275 ;
      RECT  3.64 1.275 3.735 1.35 ;
      RECT  3.555 1.35 3.735 1.45 ;
      RECT  3.78 0.77 4.105 0.86 ;
      RECT  3.78 0.86 3.87 1.0 ;
      RECT  3.405 0.51 3.51 1.0 ;
      RECT  3.405 1.0 3.87 1.09 ;
      RECT  3.405 1.09 3.505 1.26 ;
      RECT  1.935 0.425 2.035 0.96 ;
      RECT  1.555 0.41 1.655 1.09 ;
      RECT  2.135 0.91 2.235 1.41 ;
      RECT  2.075 1.41 2.235 1.58 ;
      RECT  1.555 1.18 1.655 1.54 ;
      RECT  1.555 1.54 1.77 1.66 ;
      LAYER M2 ;
      RECT  1.11 0.55 2.075 0.65 ;
      RECT  0.895 0.95 2.695 1.05 ;
      RECT  1.595 1.15 2.47 1.25 ;
      RECT  1.595 1.25 1.695 1.35 ;
      RECT  0.29 1.35 1.695 1.45 ;
      RECT  1.8 1.35 3.735 1.45 ;
      LAYER V1 ;
      RECT  1.15 0.55 1.25 0.65 ;
      RECT  1.935 0.55 2.035 0.65 ;
      RECT  0.935 0.95 1.035 1.05 ;
      RECT  1.555 0.95 1.655 1.05 ;
      RECT  2.135 0.95 2.235 1.05 ;
      RECT  2.555 0.95 2.655 1.05 ;
      RECT  2.33 1.15 2.43 1.25 ;
      RECT  0.33 1.35 0.43 1.45 ;
      RECT  1.555 1.35 1.655 1.45 ;
      RECT  1.84 1.35 1.94 1.45 ;
      RECT  3.595 1.35 3.695 1.45 ;
  END
END SEN_EO3_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_EO3_DG_8
#      Description : "3-Input exclusive OR"
#      Equation    : X=(A1^A2)^A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO3_DG_8
  CLASS CORE ;
  FOREIGN SEN_EO3_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.51 6.45 0.71 ;
      RECT  5.845 0.71 6.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1914 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.64 4.85 1.09 ;
      RECT  2.88 0.65 2.98 1.09 ;
      LAYER M2 ;
      RECT  2.84 0.95 4.89 1.05 ;
      LAYER V1 ;
      RECT  4.75 0.95 4.85 1.05 ;
      RECT  2.88 0.95 2.98 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3174 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.4 1.85 ;
      RECT  0.58 1.45 0.71 1.75 ;
      RECT  1.1 1.45 1.23 1.75 ;
      RECT  1.62 1.43 1.75 1.75 ;
      RECT  2.14 1.22 2.27 1.75 ;
      RECT  5.53 1.44 5.66 1.75 ;
      RECT  7.115 1.21 7.235 1.75 ;
      RECT  7.63 1.41 7.76 1.75 ;
      RECT  8.15 1.41 8.28 1.75 ;
      RECT  8.67 1.41 8.8 1.75 ;
      RECT  9.21 1.215 9.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      RECT  0.58 0.05 0.71 0.35 ;
      RECT  1.1 0.05 1.23 0.35 ;
      RECT  1.62 0.05 1.75 0.35 ;
      RECT  2.14 0.05 2.27 0.35 ;
      RECT  5.54 0.05 5.665 0.385 ;
      RECT  7.63 0.05 7.76 0.39 ;
      RECT  8.15 0.05 8.28 0.39 ;
      RECT  8.67 0.05 8.8 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  7.115 0.05 7.235 0.59 ;
      RECT  9.21 0.05 9.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.51 9.05 0.69 ;
      RECT  8.485 0.69 8.65 1.11 ;
      RECT  7.35 1.11 9.065 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.655 0.215 3.815 0.335 ;
      RECT  3.695 0.335 3.815 0.385 ;
      RECT  2.655 0.335 2.775 1.405 ;
      RECT  2.655 1.405 3.815 1.505 ;
      RECT  3.695 1.505 3.815 1.61 ;
      RECT  5.755 0.215 7.01 0.335 ;
      RECT  6.92 0.335 7.01 0.785 ;
      RECT  6.92 0.785 8.375 0.895 ;
      RECT  6.92 0.895 7.01 1.54 ;
      RECT  5.75 1.54 7.01 1.66 ;
      RECT  3.925 0.395 4.925 0.485 ;
      RECT  3.925 0.485 4.015 0.495 ;
      RECT  3.45 0.495 4.015 0.665 ;
      RECT  3.925 0.665 4.015 1.205 ;
      RECT  2.87 1.205 4.015 1.315 ;
      RECT  3.925 1.315 4.015 1.33 ;
      RECT  3.925 1.33 4.385 1.45 ;
      RECT  0.28 0.44 1.23 0.555 ;
      RECT  1.14 0.555 1.23 0.785 ;
      RECT  1.14 0.785 1.83 0.895 ;
      RECT  1.14 0.895 1.23 1.22 ;
      RECT  1.14 1.22 2.0 1.24 ;
      RECT  0.28 1.24 2.0 1.34 ;
      RECT  0.28 1.34 1.23 1.36 ;
      RECT  1.9 1.34 2.0 1.51 ;
      RECT  1.32 0.44 2.25 0.56 ;
      RECT  2.15 0.56 2.25 1.01 ;
      RECT  1.32 1.01 2.25 1.13 ;
      RECT  2.87 0.44 3.17 0.56 ;
      RECT  3.07 0.56 3.17 1.005 ;
      RECT  3.07 1.005 3.605 1.115 ;
      RECT  6.54 0.44 6.765 0.56 ;
      RECT  6.54 0.56 6.63 1.13 ;
      RECT  6.03 1.13 6.63 1.25 ;
      RECT  5.555 0.475 6.225 0.595 ;
      RECT  5.555 0.595 5.645 1.26 ;
      RECT  3.92 0.165 5.17 0.285 ;
      RECT  5.08 0.285 5.17 1.26 ;
      RECT  5.08 1.26 5.845 1.34 ;
      RECT  5.08 1.34 6.765 1.35 ;
      RECT  5.75 1.35 6.765 1.45 ;
      RECT  5.08 1.35 5.18 1.54 ;
      RECT  3.905 1.54 5.18 1.66 ;
      RECT  4.16 0.575 4.65 0.68 ;
      RECT  4.55 0.68 4.65 1.24 ;
      RECT  4.55 1.24 4.93 1.36 ;
      RECT  3.26 0.51 3.36 0.79 ;
      RECT  3.26 0.79 3.765 0.9 ;
      RECT  6.72 0.65 6.82 1.11 ;
      RECT  5.275 0.415 5.39 1.17 ;
      RECT  2.405 0.425 2.525 1.315 ;
      LAYER M2 ;
      RECT  2.38 0.55 3.4 0.65 ;
      RECT  2.11 0.75 4.69 0.85 ;
      RECT  5.25 0.95 6.86 1.05 ;
      RECT  2.63 1.15 6.21 1.25 ;
      RECT  1.86 1.35 4.18 1.45 ;
      LAYER V1 ;
      RECT  2.42 0.55 2.52 0.65 ;
      RECT  3.26 0.55 3.36 0.65 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  3.07 0.75 3.17 0.85 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  5.29 0.95 5.39 1.05 ;
      RECT  6.72 0.95 6.82 1.05 ;
      RECT  2.67 1.15 2.77 1.25 ;
      RECT  6.07 1.15 6.17 1.25 ;
      RECT  1.9 1.35 2.0 1.45 ;
      RECT  4.04 1.35 4.14 1.45 ;
  END
END SEN_EO3_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_EO4_DG_1
#      Description : "4-Input exclusive OR"
#      Equation    : X=((A1^A2)^A3)^A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO4_DG_1
  CLASS CORE ;
  FOREIGN SEN_EO4_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.71 5.85 0.91 ;
      RECT  5.55 0.91 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.765 ;
      RECT  0.95 0.765 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.51 4.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.455 0.45 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  1.79 1.465 1.9 1.75 ;
      RECT  3.35 1.415 3.48 1.75 ;
      RECT  3.86 1.42 3.99 1.75 ;
      RECT  5.515 1.43 5.645 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  1.85 0.05 2.02 0.215 ;
      RECT  0.38 0.05 0.5 0.39 ;
      RECT  3.355 0.05 3.48 0.39 ;
      RECT  3.86 0.05 3.99 0.39 ;
      RECT  5.51 0.05 5.64 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.055 0.23 3.265 0.35 ;
      RECT  3.175 0.35 3.265 0.48 ;
      RECT  3.175 0.48 3.45 0.57 ;
      RECT  3.35 0.57 3.45 1.015 ;
      RECT  3.045 1.015 3.45 1.12 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.14 0.14 4.98 0.23 ;
      RECT  4.87 0.23 4.98 0.925 ;
      RECT  4.14 0.23 4.25 1.585 ;
      RECT  2.845 0.18 2.965 0.305 ;
      RECT  1.95 0.305 2.965 0.4 ;
      RECT  1.95 0.4 2.05 1.265 ;
      RECT  1.61 1.265 2.08 1.355 ;
      RECT  1.61 1.355 1.7 1.445 ;
      RECT  1.99 1.355 2.08 1.57 ;
      RECT  1.08 1.445 1.7 1.555 ;
      RECT  1.99 1.57 2.41 1.66 ;
      RECT  1.365 0.19 1.485 0.35 ;
      RECT  1.365 0.35 1.69 0.45 ;
      RECT  1.055 0.27 1.275 0.39 ;
      RECT  1.185 0.39 1.275 0.55 ;
      RECT  1.185 0.55 1.49 0.65 ;
      RECT  0.065 0.215 0.29 0.48 ;
      RECT  0.065 0.48 0.515 0.57 ;
      RECT  0.425 0.57 0.515 1.275 ;
      RECT  0.065 1.275 0.645 1.365 ;
      RECT  0.555 1.365 0.645 1.445 ;
      RECT  0.065 1.365 0.185 1.53 ;
      RECT  0.555 1.445 0.99 1.555 ;
      RECT  3.615 0.2 3.735 0.48 ;
      RECT  3.615 0.48 3.845 0.57 ;
      RECT  3.755 0.57 3.845 1.21 ;
      RECT  2.35 0.755 2.44 1.21 ;
      RECT  2.35 1.21 3.845 1.3 ;
      RECT  3.615 1.3 3.845 1.33 ;
      RECT  3.615 1.33 3.735 1.58 ;
      RECT  5.815 0.22 5.935 0.48 ;
      RECT  5.335 0.48 5.935 0.57 ;
      RECT  5.335 0.57 5.46 0.9 ;
      RECT  5.37 0.9 5.46 1.25 ;
      RECT  5.115 1.25 5.935 1.34 ;
      RECT  5.115 1.34 5.205 1.455 ;
      RECT  5.815 1.34 5.935 1.6 ;
      RECT  4.865 1.455 5.205 1.575 ;
      RECT  2.53 0.495 3.08 0.605 ;
      RECT  2.99 0.605 3.08 0.755 ;
      RECT  2.53 0.605 2.62 1.015 ;
      RECT  2.99 0.755 3.26 0.925 ;
      RECT  2.53 1.015 2.7 1.12 ;
      RECT  4.35 0.32 4.52 0.89 ;
      RECT  1.58 0.54 1.75 0.99 ;
      RECT  0.965 0.99 1.75 1.1 ;
      RECT  1.58 1.1 1.75 1.135 ;
      RECT  5.145 0.22 5.245 0.99 ;
      RECT  5.145 0.99 5.28 1.07 ;
      RECT  4.935 1.07 5.28 1.16 ;
      RECT  4.935 1.16 5.025 1.25 ;
      RECT  4.375 1.25 5.025 1.34 ;
      RECT  4.375 1.34 4.495 1.585 ;
      RECT  0.74 0.2 0.86 1.01 ;
      RECT  0.605 1.01 0.86 1.185 ;
      RECT  0.75 1.185 0.86 1.22 ;
      RECT  0.75 1.22 1.52 1.33 ;
      RECT  2.8 0.695 2.9 1.12 ;
      RECT  3.54 0.67 3.64 1.12 ;
      RECT  4.61 0.32 4.78 1.16 ;
      RECT  2.17 0.49 2.26 1.39 ;
      RECT  2.17 1.39 3.015 1.48 ;
      LAYER M2 ;
      RECT  0.11 0.35 1.69 0.45 ;
      RECT  1.31 0.55 2.09 0.65 ;
      RECT  4.38 0.75 5.5 0.85 ;
      RECT  2.76 0.95 4.8 1.05 ;
      LAYER V1 ;
      RECT  0.15 0.35 0.25 0.45 ;
      RECT  1.55 0.35 1.65 0.45 ;
      RECT  1.35 0.55 1.45 0.65 ;
      RECT  1.95 0.55 2.05 0.65 ;
      RECT  4.42 0.75 4.52 0.85 ;
      RECT  5.36 0.75 5.46 0.85 ;
      RECT  2.8 0.95 2.9 1.05 ;
      RECT  3.54 0.95 3.64 1.05 ;
      RECT  4.66 0.95 4.76 1.05 ;
  END
END SEN_EO4_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_EO4_DG_2
#      Description : "4-Input exclusive OR"
#      Equation    : X=((A1^A2)^A3)^A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO4_DG_2
  CLASS CORE ;
  FOREIGN SEN_EO4_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.69 0.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.69 6.05 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.745 ;
      RECT  0.95 0.745 1.485 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.51 4.25 0.755 ;
      RECT  4.15 0.755 4.32 0.925 ;
      RECT  4.15 0.925 4.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.45 0.46 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  1.83 1.46 1.96 1.75 ;
      RECT  3.14 1.4 3.27 1.75 ;
      RECT  3.66 1.4 3.79 1.75 ;
      RECT  4.17 1.39 4.3 1.75 ;
      RECT  5.74 1.43 5.87 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  1.85 0.05 2.02 0.19 ;
      RECT  0.34 0.05 0.46 0.36 ;
      RECT  3.14 0.05 3.27 0.38 ;
      RECT  3.66 0.05 3.79 0.39 ;
      RECT  4.17 0.05 4.3 0.39 ;
      RECT  5.74 0.05 5.87 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.65 0.69 ;
      RECT  3.55 0.69 3.65 1.0 ;
      RECT  3.38 1.0 3.65 1.12 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.435 0.14 5.265 0.23 ;
      RECT  5.165 0.23 5.265 0.9 ;
      RECT  4.435 0.23 4.555 1.59 ;
      RECT  1.87 0.28 3.05 0.38 ;
      RECT  1.87 0.38 1.97 0.705 ;
      RECT  1.87 0.705 2.115 0.875 ;
      RECT  1.87 0.875 1.96 1.28 ;
      RECT  1.61 1.28 2.14 1.37 ;
      RECT  1.61 1.37 1.7 1.47 ;
      RECT  2.05 1.37 2.14 1.57 ;
      RECT  1.08 1.47 1.7 1.585 ;
      RECT  2.05 1.57 2.51 1.66 ;
      RECT  1.105 0.215 1.24 0.385 ;
      RECT  1.14 0.385 1.24 0.55 ;
      RECT  1.14 0.55 1.37 0.65 ;
      RECT  0.605 0.28 1.015 0.4 ;
      RECT  0.605 0.4 0.71 1.08 ;
      RECT  0.605 1.08 0.845 1.17 ;
      RECT  0.755 1.17 0.845 1.275 ;
      RECT  0.755 1.275 1.52 1.38 ;
      RECT  1.335 0.215 1.515 0.45 ;
      RECT  0.075 0.31 0.25 0.46 ;
      RECT  0.075 0.46 0.465 0.56 ;
      RECT  0.375 0.56 0.465 0.755 ;
      RECT  0.375 0.755 0.515 0.925 ;
      RECT  0.375 0.925 0.465 1.24 ;
      RECT  0.075 1.24 0.465 1.26 ;
      RECT  0.075 1.26 0.645 1.36 ;
      RECT  0.075 1.36 0.195 1.47 ;
      RECT  0.555 1.36 0.645 1.47 ;
      RECT  0.555 1.47 0.99 1.585 ;
      RECT  6.015 0.25 6.135 0.5 ;
      RECT  5.685 0.5 6.135 0.59 ;
      RECT  5.685 0.59 5.795 0.71 ;
      RECT  5.595 0.71 5.795 0.89 ;
      RECT  5.685 0.89 5.795 1.25 ;
      RECT  5.49 1.25 6.135 1.34 ;
      RECT  5.49 1.34 5.58 1.465 ;
      RECT  6.015 1.34 6.135 1.53 ;
      RECT  5.175 1.465 5.58 1.585 ;
      RECT  2.59 0.47 3.255 0.56 ;
      RECT  3.165 0.56 3.255 0.785 ;
      RECT  2.59 0.56 2.71 1.015 ;
      RECT  3.165 0.785 3.46 0.895 ;
      RECT  2.59 1.015 2.76 1.12 ;
      RECT  2.13 0.47 2.32 0.59 ;
      RECT  2.215 0.59 2.32 1.02 ;
      RECT  2.105 1.02 2.32 1.19 ;
      RECT  2.23 1.19 2.32 1.39 ;
      RECT  2.23 1.39 3.05 1.48 ;
      RECT  4.685 0.32 4.805 0.97 ;
      RECT  5.36 0.24 5.48 0.99 ;
      RECT  5.36 0.99 5.58 1.07 ;
      RECT  5.31 1.07 5.58 1.16 ;
      RECT  5.31 1.16 5.4 1.285 ;
      RECT  4.685 1.285 5.4 1.375 ;
      RECT  4.685 1.375 4.805 1.53 ;
      RECT  1.005 0.99 1.115 1.07 ;
      RECT  1.005 1.07 1.725 1.16 ;
      RECT  1.605 0.37 1.725 1.07 ;
      RECT  3.74 0.62 3.85 1.09 ;
      RECT  2.85 0.67 2.955 1.12 ;
      RECT  4.955 0.32 5.075 1.16 ;
      RECT  2.41 0.785 2.5 1.21 ;
      RECT  2.41 1.21 4.045 1.3 ;
      RECT  3.94 0.2 4.045 1.21 ;
      RECT  3.925 1.3 4.045 1.58 ;
      LAYER M2 ;
      RECT  0.11 0.35 1.515 0.45 ;
      RECT  1.19 0.55 2.01 0.65 ;
      RECT  4.66 0.75 5.735 0.85 ;
      RECT  2.815 0.95 5.11 1.05 ;
      LAYER V1 ;
      RECT  0.15 0.35 0.25 0.45 ;
      RECT  1.375 0.35 1.475 0.45 ;
      RECT  1.23 0.55 1.33 0.65 ;
      RECT  1.87 0.55 1.97 0.65 ;
      RECT  4.7 0.75 4.8 0.85 ;
      RECT  5.595 0.75 5.695 0.85 ;
      RECT  2.855 0.95 2.955 1.05 ;
      RECT  3.745 0.95 3.845 1.05 ;
      RECT  4.97 0.95 5.07 1.05 ;
  END
END SEN_EO4_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_EO4_DG_3
#      Description : "4-Input exclusive OR"
#      Equation    : X=((A1^A2)^A3)^A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO4_DG_3
  CLASS CORE ;
  FOREIGN SEN_EO4_DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.71 6.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.825 2.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0759 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.67 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0759 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.215 0.185 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.58 1.45 0.705 1.75 ;
      RECT  1.125 1.45 1.245 1.75 ;
      RECT  2.42 1.57 2.54 1.75 ;
      RECT  4.015 1.44 4.135 1.75 ;
      RECT  4.525 1.44 4.645 1.75 ;
      RECT  5.045 1.44 5.165 1.75 ;
      RECT  6.53 1.575 6.7 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  0.57 0.05 0.74 0.195 ;
      RECT  1.11 0.05 1.28 0.195 ;
      RECT  2.435 0.05 2.605 0.26 ;
      RECT  3.99 0.05 4.16 0.28 ;
      RECT  4.525 0.05 4.645 0.385 ;
      RECT  5.055 0.05 5.175 0.385 ;
      RECT  6.55 0.05 6.67 0.385 ;
      RECT  0.065 0.05 0.185 0.535 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.265 0.51 5.05 0.69 ;
      RECT  4.95 0.69 5.05 1.04 ;
      RECT  4.24 1.04 5.05 1.155 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.315 0.14 6.21 0.23 ;
      RECT  6.12 0.23 6.21 0.925 ;
      RECT  5.315 0.23 5.435 1.17 ;
      RECT  1.455 0.15 2.075 0.26 ;
      RECT  1.455 0.26 1.545 0.285 ;
      RECT  0.3 0.285 1.545 0.38 ;
      RECT  0.3 0.38 0.74 0.385 ;
      RECT  0.65 0.385 0.74 0.785 ;
      RECT  0.65 0.785 1.0 0.895 ;
      RECT  0.65 0.895 0.74 1.235 ;
      RECT  0.3 1.235 0.74 1.25 ;
      RECT  0.3 1.25 1.545 1.36 ;
      RECT  2.955 0.165 3.625 0.28 ;
      RECT  2.955 0.28 3.045 0.35 ;
      RECT  1.635 0.35 3.045 0.44 ;
      RECT  1.635 0.44 2.63 0.455 ;
      RECT  2.54 0.455 2.63 0.785 ;
      RECT  2.54 0.785 2.69 0.955 ;
      RECT  2.54 0.955 2.63 1.39 ;
      RECT  2.155 1.39 2.72 1.44 ;
      RECT  1.635 1.44 2.72 1.48 ;
      RECT  1.635 1.48 2.245 1.56 ;
      RECT  2.63 1.48 2.72 1.57 ;
      RECT  2.63 1.57 3.1 1.66 ;
      RECT  3.2 0.37 4.175 0.46 ;
      RECT  4.085 0.46 4.175 0.785 ;
      RECT  3.2 0.46 3.32 1.0 ;
      RECT  4.085 0.785 4.86 0.895 ;
      RECT  3.2 1.0 3.375 1.12 ;
      RECT  5.58 0.365 5.84 0.485 ;
      RECT  5.74 0.485 5.84 0.73 ;
      RECT  6.825 0.37 6.945 0.51 ;
      RECT  6.5 0.51 6.945 0.6 ;
      RECT  6.5 0.6 6.6 1.38 ;
      RECT  6.5 1.38 6.945 1.395 ;
      RECT  6.1 1.395 6.945 1.485 ;
      RECT  6.825 1.485 6.945 1.56 ;
      RECT  6.1 1.485 6.205 1.61 ;
      RECT  0.84 0.47 1.545 0.59 ;
      RECT  1.155 0.59 1.245 1.04 ;
      RECT  0.83 1.04 1.245 1.07 ;
      RECT  0.83 1.07 2.035 1.16 ;
      RECT  1.925 1.16 2.035 1.34 ;
      RECT  3.555 0.55 3.89 0.66 ;
      RECT  3.555 0.66 3.645 1.21 ;
      RECT  3.01 0.78 3.11 1.21 ;
      RECT  3.01 1.21 3.85 1.3 ;
      RECT  3.745 1.3 3.85 1.515 ;
      RECT  2.155 0.545 2.325 0.665 ;
      RECT  2.155 0.665 2.26 0.855 ;
      RECT  1.45 0.855 2.26 0.965 ;
      RECT  2.155 0.965 2.26 1.23 ;
      RECT  2.81 0.575 2.98 0.665 ;
      RECT  2.81 0.665 2.9 1.13 ;
      RECT  2.72 1.13 2.9 1.3 ;
      RECT  2.81 1.3 2.9 1.39 ;
      RECT  2.81 1.39 3.615 1.48 ;
      RECT  3.495 1.48 3.615 1.61 ;
      RECT  5.93 0.375 6.03 1.015 ;
      RECT  5.74 1.015 6.03 1.125 ;
      RECT  5.74 1.125 5.83 1.26 ;
      RECT  3.745 0.755 3.855 0.985 ;
      RECT  3.745 0.985 4.03 1.075 ;
      RECT  3.94 1.075 4.03 1.26 ;
      RECT  3.94 1.26 5.83 1.35 ;
      RECT  6.3 0.37 6.41 1.215 ;
      RECT  5.92 1.215 6.41 1.305 ;
      RECT  5.92 1.305 6.01 1.465 ;
      RECT  5.52 1.465 6.01 1.585 ;
      LAYER M2 ;
      RECT  5.7 0.55 6.64 0.65 ;
      LAYER V1 ;
      RECT  5.74 0.55 5.84 0.65 ;
      RECT  6.5 0.55 6.6 0.65 ;
  END
END SEN_EO4_DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_EO4_DG_4
#      Description : "4-Input exclusive OR"
#      Equation    : X=((A1^A2)^A3)^A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_EO4_DG_4
  CLASS CORE ;
  FOREIGN SEN_EO4_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.71 6.85 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.835 0.54 2.05 0.65 ;
      RECT  1.95 0.65 2.05 0.925 ;
      LAYER M2 ;
      RECT  1.91 0.75 2.535 0.85 ;
      LAYER V1 ;
      RECT  1.95 0.75 2.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 5.85 0.71 ;
      RECT  5.54 0.71 5.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.58 1.45 0.71 1.75 ;
      RECT  1.08 1.45 1.25 1.75 ;
      RECT  2.39 1.44 2.515 1.75 ;
      RECT  3.935 1.44 4.065 1.75 ;
      RECT  4.455 1.44 4.585 1.75 ;
      RECT  4.995 1.44 5.125 1.75 ;
      RECT  6.545 1.455 6.675 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  3.915 0.05 4.085 0.305 ;
      RECT  0.595 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  6.545 0.05 6.66 0.36 ;
      RECT  4.475 0.05 4.605 0.39 ;
      RECT  5.0 0.05 5.13 0.39 ;
      RECT  2.38 0.05 2.49 0.43 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.235 0.51 5.05 0.69 ;
      RECT  4.95 0.69 5.05 1.04 ;
      RECT  4.145 1.04 5.05 1.16 ;
    END
    ANTENNADIFFAREA 0.454 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.27 0.14 6.21 0.23 ;
      RECT  6.12 0.23 6.21 0.925 ;
      RECT  5.27 0.23 5.39 1.16 ;
      RECT  2.58 0.2 3.61 0.305 ;
      RECT  2.58 0.305 2.68 0.73 ;
      RECT  2.545 0.73 2.68 0.9 ;
      RECT  2.545 0.9 2.635 1.26 ;
      RECT  2.14 1.26 2.695 1.35 ;
      RECT  2.14 1.35 2.23 1.48 ;
      RECT  2.605 1.35 2.695 1.57 ;
      RECT  1.56 1.48 2.23 1.6 ;
      RECT  2.605 1.57 3.025 1.66 ;
      RECT  0.325 0.35 0.505 0.45 ;
      RECT  0.325 0.45 0.645 0.54 ;
      RECT  0.555 0.54 0.645 0.785 ;
      RECT  0.555 0.785 1.02 0.895 ;
      RECT  0.555 0.895 0.645 1.24 ;
      RECT  0.275 1.24 1.5 1.36 ;
      RECT  1.835 0.19 2.015 0.45 ;
      RECT  5.48 0.32 5.665 0.45 ;
      RECT  5.48 0.45 5.6 0.61 ;
      RECT  6.75 0.31 6.93 0.45 ;
      RECT  6.54 0.45 6.93 0.54 ;
      RECT  6.54 0.54 6.63 0.755 ;
      RECT  6.49 0.755 6.63 0.925 ;
      RECT  6.54 0.925 6.63 1.265 ;
      RECT  6.355 1.265 6.93 1.365 ;
      RECT  6.355 1.365 6.445 1.465 ;
      RECT  6.81 1.365 6.93 1.49 ;
      RECT  5.99 1.465 6.445 1.585 ;
      RECT  3.145 0.395 4.145 0.485 ;
      RECT  4.055 0.485 4.145 0.785 ;
      RECT  3.145 0.485 3.265 1.01 ;
      RECT  4.055 0.785 4.665 0.895 ;
      RECT  3.145 1.01 3.34 1.11 ;
      RECT  0.795 0.45 1.52 0.57 ;
      RECT  1.155 0.57 1.245 1.03 ;
      RECT  0.795 1.03 1.68 1.15 ;
      RECT  1.59 1.15 1.68 1.24 ;
      RECT  1.59 1.24 2.05 1.36 ;
      RECT  3.52 0.575 3.83 0.675 ;
      RECT  3.52 0.675 3.61 1.2 ;
      RECT  2.965 0.75 3.055 1.2 ;
      RECT  2.965 1.2 3.785 1.29 ;
      RECT  3.68 1.29 3.785 1.53 ;
      RECT  1.615 0.2 1.735 0.69 ;
      RECT  1.375 0.785 1.86 0.895 ;
      RECT  1.77 0.895 1.86 1.015 ;
      RECT  1.77 1.015 2.27 1.135 ;
      RECT  2.14 0.21 2.27 1.015 ;
      RECT  2.78 0.415 2.875 1.0 ;
      RECT  2.725 1.0 2.875 1.17 ;
      RECT  2.785 1.17 2.875 1.38 ;
      RECT  2.785 1.38 3.59 1.48 ;
      RECT  5.94 0.45 6.03 1.025 ;
      RECT  5.555 1.025 6.03 1.145 ;
      RECT  5.555 1.145 5.645 1.26 ;
      RECT  3.7 0.785 3.965 0.895 ;
      RECT  3.875 0.895 3.965 1.26 ;
      RECT  3.875 1.26 5.645 1.35 ;
      RECT  6.3 0.415 6.4 1.08 ;
      RECT  6.155 1.08 6.4 1.17 ;
      RECT  6.155 1.17 6.245 1.26 ;
      RECT  5.755 1.26 6.245 1.35 ;
      RECT  5.755 1.35 5.845 1.465 ;
      RECT  5.47 1.465 5.845 1.585 ;
      LAYER M2 ;
      RECT  0.325 0.35 2.015 0.45 ;
      RECT  5.48 0.35 6.89 0.45 ;
      RECT  1.585 0.55 2.72 0.65 ;
      LAYER V1 ;
      RECT  0.365 0.35 0.465 0.45 ;
      RECT  1.875 0.35 1.975 0.45 ;
      RECT  5.52 0.35 5.62 0.45 ;
      RECT  6.75 0.35 6.85 0.45 ;
      RECT  1.625 0.55 1.725 0.65 ;
      RECT  2.58 0.55 2.68 0.65 ;
  END
END SEN_EO4_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDAO22PQ_1
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((A1&A2)|(B1&B2))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDAO22PQ_1
  CLASS CORE ;
  FOREIGN SEN_FDAO22PQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END B2
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.072 ;
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.31 5.535 0.485 ;
      RECT  5.35 0.485 5.45 1.115 ;
      RECT  5.35 1.115 5.535 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  2.33 1.615 2.5 1.75 ;
      RECT  3.8 1.51 3.97 1.75 ;
      RECT  4.63 1.395 4.76 1.75 ;
      RECT  5.15 1.38 5.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  4.62 0.05 4.79 0.185 ;
      RECT  2.475 0.05 2.645 0.245 ;
      RECT  3.82 0.05 3.95 0.33 ;
      RECT  1.135 0.05 1.26 0.385 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  5.15 0.05 5.26 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.35 0.14 2.31 0.245 ;
      RECT  2.205 0.245 2.31 0.335 ;
      RECT  2.205 0.335 3.125 0.425 ;
      RECT  2.205 0.425 2.31 0.54 ;
      RECT  3.02 0.425 3.125 1.115 ;
      RECT  2.095 0.54 2.31 0.63 ;
      RECT  2.095 0.63 2.185 1.165 ;
      RECT  2.975 1.115 3.125 1.285 ;
      RECT  4.895 0.215 5.015 0.275 ;
      RECT  4.19 0.275 5.015 0.365 ;
      RECT  4.19 0.365 4.28 0.42 ;
      RECT  4.895 0.365 5.015 1.62 ;
      RECT  3.745 0.42 4.28 0.51 ;
      RECT  3.745 0.51 3.835 1.01 ;
      RECT  1.42 0.335 2.105 0.445 ;
      RECT  1.42 0.445 1.51 0.475 ;
      RECT  0.535 0.24 1.03 0.36 ;
      RECT  0.94 0.36 1.03 0.475 ;
      RECT  0.94 0.475 1.51 0.565 ;
      RECT  1.34 0.565 1.43 1.225 ;
      RECT  0.815 1.225 1.43 1.255 ;
      RECT  0.815 1.255 1.68 1.345 ;
      RECT  3.925 0.64 4.275 0.73 ;
      RECT  3.925 0.73 4.025 1.135 ;
      RECT  3.925 1.135 4.27 1.24 ;
      RECT  2.77 0.515 2.875 0.755 ;
      RECT  2.275 0.755 2.875 0.845 ;
      RECT  2.785 0.845 2.875 1.225 ;
      RECT  2.575 1.225 2.875 1.345 ;
      RECT  4.37 0.5 4.46 0.885 ;
      RECT  4.115 0.885 4.46 0.995 ;
      RECT  4.37 0.995 4.46 1.33 ;
      RECT  3.62 1.33 4.46 1.42 ;
      RECT  3.62 1.42 3.71 1.435 ;
      RECT  1.965 1.435 3.71 1.525 ;
      RECT  1.965 1.525 2.055 1.63 ;
      RECT  2.805 1.525 2.915 1.66 ;
      RECT  2.395 0.975 2.67 1.085 ;
      RECT  2.395 1.085 2.485 1.255 ;
      RECT  1.62 0.54 1.92 0.645 ;
      RECT  1.8 0.645 1.92 1.255 ;
      RECT  1.8 1.255 2.485 1.345 ;
      RECT  5.15 0.51 5.25 1.09 ;
      RECT  3.295 0.51 3.395 1.115 ;
      RECT  3.235 1.115 3.395 1.285 ;
      RECT  3.56 0.515 3.655 1.135 ;
      RECT  3.505 1.135 3.72 1.24 ;
      RECT  1.55 0.735 1.65 1.165 ;
      RECT  0.065 1.26 0.705 1.35 ;
      RECT  0.585 1.35 0.705 1.44 ;
      RECT  0.065 1.35 0.185 1.485 ;
      RECT  0.585 1.44 1.31 1.56 ;
      LAYER M2 ;
      RECT  3.22 0.55 5.32 0.65 ;
      RECT  1.48 0.95 4.09 1.05 ;
      LAYER V1 ;
      RECT  3.295 0.55 3.395 0.65 ;
      RECT  5.15 0.55 5.25 0.65 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  3.925 0.95 4.025 1.05 ;
  END
END SEN_FDAO22PQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNQ_1
#      Description : "D-Flip Flop, neg-edge triggered"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNQ_1
  CLASS CORE ;
  FOREIGN SEN_FDNQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.225 0.65 3.325 1.09 ;
      RECT  0.52 0.85 0.625 0.95 ;
      RECT  0.275 0.95 0.625 1.055 ;
      LAYER M2 ;
      RECT  0.41 0.95 3.39 1.05 ;
      LAYER V1 ;
      RECT  3.225 0.95 3.325 1.05 ;
      RECT  0.48 0.95 0.58 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0915 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.92 0.51 1.05 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.31 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.57 0.2 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.775 1.555 0.925 1.75 ;
      RECT  1.825 1.46 1.955 1.75 ;
      RECT  2.305 1.44 2.475 1.75 ;
      RECT  3.795 1.395 3.9 1.75 ;
      RECT  4.065 1.21 4.185 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  1.985 0.05 2.155 0.35 ;
      RECT  2.475 0.05 2.645 0.355 ;
      RECT  0.795 0.05 0.935 0.36 ;
      RECT  3.475 0.05 3.61 0.36 ;
      RECT  0.32 0.05 0.465 0.58 ;
      RECT  4.065 0.05 4.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.97 0.215 3.335 0.335 ;
      RECT  3.245 0.335 3.335 0.47 ;
      RECT  3.245 0.47 3.705 0.56 ;
      RECT  3.615 0.56 3.705 0.73 ;
      RECT  3.615 0.73 3.795 0.9 ;
      RECT  3.615 0.9 3.705 1.465 ;
      RECT  3.225 1.465 3.705 1.585 ;
      RECT  3.7 0.21 3.885 0.38 ;
      RECT  3.795 0.38 3.885 0.42 ;
      RECT  3.795 0.42 3.975 0.59 ;
      RECT  3.885 0.59 3.975 1.02 ;
      RECT  3.795 1.02 3.975 1.19 ;
      RECT  1.125 0.2 1.23 0.4 ;
      RECT  1.14 0.4 1.23 0.99 ;
      RECT  1.015 0.99 1.23 1.105 ;
      RECT  2.27 0.275 2.385 0.445 ;
      RECT  2.27 0.445 2.505 0.535 ;
      RECT  2.405 0.535 2.505 1.025 ;
      RECT  1.79 0.88 1.885 1.025 ;
      RECT  1.79 1.025 2.505 1.145 ;
      RECT  1.51 0.2 1.63 0.45 ;
      RECT  1.34 0.45 2.125 0.54 ;
      RECT  2.035 0.54 2.125 0.625 ;
      RECT  1.34 0.54 1.44 1.08 ;
      RECT  2.035 0.625 2.28 0.715 ;
      RECT  2.17 0.715 2.28 0.875 ;
      RECT  2.595 0.445 3.125 0.56 ;
      RECT  3.035 0.56 3.125 1.16 ;
      RECT  2.595 0.56 2.715 1.17 ;
      RECT  2.845 0.735 2.945 0.86 ;
      RECT  2.805 0.86 2.945 0.965 ;
      RECT  2.805 0.965 2.895 1.25 ;
      RECT  2.805 1.25 3.525 1.26 ;
      RECT  3.435 1.18 3.525 1.25 ;
      RECT  1.61 0.63 1.85 0.735 ;
      RECT  1.61 0.735 1.7 1.26 ;
      RECT  1.61 1.26 3.525 1.35 ;
      RECT  1.61 1.35 1.7 1.38 ;
      RECT  0.595 0.41 0.715 0.67 ;
      RECT  0.275 0.67 0.805 0.76 ;
      RECT  0.275 0.76 0.365 0.86 ;
      RECT  0.715 0.76 0.805 1.17 ;
      RECT  0.45 1.17 0.805 1.195 ;
      RECT  0.45 1.195 1.285 1.285 ;
      RECT  1.195 1.285 1.285 1.38 ;
      RECT  1.195 1.38 1.7 1.48 ;
      RECT  0.09 0.37 0.18 1.375 ;
      RECT  0.09 1.375 1.105 1.465 ;
      RECT  1.015 1.465 1.105 1.57 ;
      RECT  0.335 1.465 0.455 1.59 ;
      RECT  1.015 1.57 1.67 1.66 ;
  END
END SEN_FDNQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNQ_2
#      Description : "D-Flip Flop, neg-edge triggered"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNQ_2
  CLASS CORE ;
  FOREIGN SEN_FDNQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.665 0.65 3.765 1.09 ;
      RECT  0.455 0.74 0.595 0.92 ;
      RECT  0.455 0.92 0.56 0.95 ;
      RECT  0.275 0.95 0.56 1.05 ;
      LAYER M2 ;
      RECT  0.35 0.95 3.84 1.05 ;
      LAYER V1 ;
      RECT  3.665 0.95 3.765 1.05 ;
      RECT  0.42 0.95 0.52 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1167 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.92 0.51 1.05 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0552 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.31 4.865 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.495 0.47 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.775 1.555 0.91 1.75 ;
      RECT  1.825 1.44 1.955 1.75 ;
      RECT  2.385 1.44 2.555 1.75 ;
      RECT  2.915 1.44 3.07 1.75 ;
      RECT  4.225 1.39 4.335 1.75 ;
      RECT  4.495 1.21 4.615 1.75 ;
      RECT  5.015 1.21 5.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.815 0.05 2.985 0.34 ;
      RECT  2.02 0.05 2.19 0.35 ;
      RECT  3.905 0.05 4.04 0.36 ;
      RECT  0.8 0.05 0.935 0.39 ;
      RECT  0.31 0.05 0.455 0.47 ;
      RECT  5.015 0.05 5.135 0.585 ;
      RECT  4.495 0.05 4.615 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.41 0.215 3.765 0.335 ;
      RECT  3.675 0.335 3.765 0.47 ;
      RECT  3.675 0.47 4.135 0.56 ;
      RECT  4.045 0.56 4.135 0.7 ;
      RECT  4.045 0.7 4.225 0.9 ;
      RECT  4.045 0.9 4.135 1.465 ;
      RECT  3.165 1.465 4.135 1.585 ;
      RECT  4.13 0.21 4.315 0.38 ;
      RECT  4.225 0.38 4.315 0.42 ;
      RECT  4.225 0.42 4.405 0.59 ;
      RECT  4.315 0.59 4.405 1.02 ;
      RECT  4.225 1.02 4.405 1.19 ;
      RECT  1.12 0.2 1.23 0.4 ;
      RECT  1.14 0.4 1.23 0.99 ;
      RECT  1.01 0.99 1.23 1.105 ;
      RECT  2.58 0.31 2.7 0.44 ;
      RECT  2.58 0.44 3.57 0.53 ;
      RECT  2.675 0.53 3.57 0.555 ;
      RECT  3.47 0.555 3.57 1.16 ;
      RECT  2.675 0.555 2.795 1.17 ;
      RECT  1.51 0.2 1.63 0.45 ;
      RECT  1.34 0.45 2.205 0.54 ;
      RECT  2.115 0.54 2.205 0.8 ;
      RECT  1.34 0.54 1.44 1.16 ;
      RECT  2.115 0.8 2.39 0.9 ;
      RECT  2.35 0.19 2.465 0.62 ;
      RECT  2.35 0.62 2.585 0.71 ;
      RECT  2.485 0.71 2.585 1.025 ;
      RECT  1.83 0.88 1.925 1.025 ;
      RECT  1.83 1.025 2.585 1.145 ;
      RECT  3.275 0.735 3.375 0.86 ;
      RECT  3.235 0.86 3.375 0.965 ;
      RECT  3.235 0.965 3.325 1.25 ;
      RECT  3.235 1.25 3.955 1.26 ;
      RECT  3.865 1.15 3.955 1.25 ;
      RECT  1.65 0.63 1.85 0.735 ;
      RECT  1.65 0.735 1.74 1.25 ;
      RECT  0.585 0.385 0.705 0.56 ;
      RECT  0.265 0.56 0.83 0.65 ;
      RECT  0.265 0.65 0.355 0.86 ;
      RECT  0.74 0.65 0.83 1.135 ;
      RECT  0.59 1.135 0.83 1.195 ;
      RECT  0.59 1.195 1.255 1.225 ;
      RECT  0.74 1.225 1.255 1.25 ;
      RECT  0.74 1.25 1.74 1.26 ;
      RECT  0.74 1.26 3.955 1.285 ;
      RECT  1.17 1.285 3.955 1.34 ;
      RECT  1.66 1.34 3.955 1.35 ;
      RECT  0.065 0.34 0.17 1.315 ;
      RECT  0.065 1.315 0.655 1.375 ;
      RECT  0.065 1.375 1.085 1.405 ;
      RECT  0.565 1.405 1.085 1.43 ;
      RECT  0.065 1.405 0.185 1.59 ;
      RECT  0.565 1.43 1.615 1.465 ;
      RECT  0.995 1.465 1.615 1.52 ;
  END
END SEN_FDNQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNQ_4
#      Description : "D-Flip Flop, neg-edge triggered"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNQ_4
  CLASS CORE ;
  FOREIGN SEN_FDNQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.65 4.455 1.11 ;
      RECT  0.455 0.74 0.615 0.92 ;
      RECT  0.455 0.92 0.58 0.95 ;
      RECT  0.275 0.95 0.58 1.05 ;
      LAYER M2 ;
      RECT  0.35 0.95 4.495 1.05 ;
      LAYER V1 ;
      RECT  4.355 0.95 4.455 1.05 ;
      RECT  0.42 0.95 0.52 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1566 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.105 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0714 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.44 0.45 5.565 0.91 ;
      RECT  5.44 0.91 6.075 1.09 ;
      RECT  5.95 0.31 6.075 0.91 ;
      RECT  5.44 1.09 5.565 1.185 ;
      RECT  5.95 1.09 6.075 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.575 0.48 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.86 1.555 0.99 1.75 ;
      RECT  1.905 1.44 2.025 1.75 ;
      RECT  2.19 1.44 2.36 1.75 ;
      RECT  2.73 1.44 2.88 1.75 ;
      RECT  3.25 1.44 3.4 1.75 ;
      RECT  4.915 1.38 5.025 1.75 ;
      RECT  5.185 1.21 5.305 1.75 ;
      RECT  5.705 1.21 5.825 1.75 ;
      RECT  6.22 1.41 6.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  1.04 0.05 1.215 0.24 ;
      RECT  2.095 0.05 2.265 0.35 ;
      RECT  4.595 0.05 4.73 0.36 ;
      RECT  3.17 0.05 3.32 0.39 ;
      RECT  5.18 0.05 5.31 0.39 ;
      RECT  6.22 0.05 6.345 0.39 ;
      RECT  2.66 0.05 2.79 0.45 ;
      RECT  0.32 0.05 0.465 0.47 ;
      RECT  5.705 0.05 5.825 0.68 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.805 0.18 0.915 0.33 ;
      RECT  0.805 0.33 1.455 0.42 ;
      RECT  1.335 0.22 1.455 0.33 ;
      RECT  1.225 0.42 1.455 0.44 ;
      RECT  1.225 0.44 1.315 0.99 ;
      RECT  1.09 0.99 1.315 1.105 ;
      RECT  3.58 0.215 4.455 0.335 ;
      RECT  4.365 0.335 4.455 0.47 ;
      RECT  4.365 0.47 4.825 0.56 ;
      RECT  4.735 0.56 4.825 0.76 ;
      RECT  4.735 0.76 5.17 0.87 ;
      RECT  4.735 0.87 4.825 1.465 ;
      RECT  3.79 1.465 4.825 1.585 ;
      RECT  4.82 0.21 5.02 0.38 ;
      RECT  4.915 0.38 5.02 0.5 ;
      RECT  4.915 0.5 5.35 0.59 ;
      RECT  5.26 0.59 5.35 0.99 ;
      RECT  4.915 0.99 5.35 1.08 ;
      RECT  4.915 1.08 5.02 1.21 ;
      RECT  3.865 0.43 4.035 0.44 ;
      RECT  3.6 0.44 4.255 0.53 ;
      RECT  2.87 0.53 4.255 0.555 ;
      RECT  2.87 0.555 3.69 0.65 ;
      RECT  4.135 0.555 4.255 1.16 ;
      RECT  3.6 0.65 3.69 1.05 ;
      RECT  2.95 1.05 3.69 1.17 ;
      RECT  1.595 0.2 1.715 0.45 ;
      RECT  1.555 0.45 2.29 0.54 ;
      RECT  2.2 0.54 2.29 0.745 ;
      RECT  1.555 0.54 1.645 0.905 ;
      RECT  2.2 0.745 2.515 0.845 ;
      RECT  1.42 0.905 1.645 0.995 ;
      RECT  1.42 0.995 1.53 1.16 ;
      RECT  2.405 0.26 2.525 0.565 ;
      RECT  2.405 0.565 2.72 0.655 ;
      RECT  2.625 0.655 2.72 0.77 ;
      RECT  2.625 0.77 3.32 0.88 ;
      RECT  2.625 0.88 2.72 1.025 ;
      RECT  1.915 0.88 2.015 1.025 ;
      RECT  1.915 1.025 2.72 1.145 ;
      RECT  3.815 0.69 4.02 0.8 ;
      RECT  3.815 0.8 3.905 1.25 ;
      RECT  3.815 1.25 4.645 1.26 ;
      RECT  4.555 1.15 4.645 1.25 ;
      RECT  1.735 0.63 1.94 0.735 ;
      RECT  1.735 0.735 1.825 1.25 ;
      RECT  0.605 0.42 0.715 0.56 ;
      RECT  0.265 0.56 0.85 0.65 ;
      RECT  0.265 0.65 0.355 0.86 ;
      RECT  0.76 0.65 0.85 1.165 ;
      RECT  0.55 1.165 0.85 1.195 ;
      RECT  0.55 1.195 1.335 1.25 ;
      RECT  0.55 1.25 1.825 1.26 ;
      RECT  0.55 1.26 4.645 1.285 ;
      RECT  1.25 1.285 4.645 1.34 ;
      RECT  1.745 1.34 4.645 1.35 ;
      RECT  0.065 0.35 0.17 1.375 ;
      RECT  0.065 1.375 1.165 1.43 ;
      RECT  0.065 1.43 1.7 1.465 ;
      RECT  1.075 1.465 1.7 1.52 ;
  END
END SEN_FDNQ_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNQ_D_1
#      Description : "D-Flip Flop, neg-edge triggered"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FDNQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.34 0.31 3.46 1.29 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.8 1.415 0.93 1.75 ;
      RECT  1.785 1.575 1.91 1.75 ;
      RECT  2.79 1.56 2.92 1.75 ;
      RECT  3.6 1.21 3.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.795 0.05 0.925 0.39 ;
      RECT  1.8 0.05 1.925 0.39 ;
      RECT  2.79 0.05 2.92 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.6 0.05 3.72 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.25 0.185 1.71 0.3 ;
      RECT  1.62 0.3 1.71 0.74 ;
      RECT  1.39 0.74 1.98 0.83 ;
      RECT  1.88 0.66 1.98 0.74 ;
      RECT  1.39 0.83 1.48 1.31 ;
      RECT  1.24 1.31 1.48 1.43 ;
      RECT  2.27 0.22 2.55 0.34 ;
      RECT  2.46 0.34 2.55 0.88 ;
      RECT  2.46 0.88 2.975 0.97 ;
      RECT  2.875 0.97 2.975 1.33 ;
      RECT  2.27 1.33 2.975 1.45 ;
      RECT  1.42 0.39 1.53 0.55 ;
      RECT  1.2 0.55 1.53 0.65 ;
      RECT  1.2 0.65 1.3 0.97 ;
      RECT  3.065 0.26 3.185 0.59 ;
      RECT  2.64 0.59 3.185 0.705 ;
      RECT  3.065 0.705 3.185 0.755 ;
      RECT  3.065 0.755 3.25 0.925 ;
      RECT  3.065 0.925 3.185 1.46 ;
      RECT  0.34 0.505 0.51 0.91 ;
      RECT  0.34 0.91 0.45 1.39 ;
      RECT  2.26 0.485 2.36 1.105 ;
      RECT  2.26 1.105 2.64 1.215 ;
      RECT  1.65 0.92 1.765 1.185 ;
      RECT  1.65 1.185 2.17 1.29 ;
      RECT  2.07 0.245 2.17 1.185 ;
      RECT  1.57 1.385 2.095 1.475 ;
      RECT  1.57 1.475 1.66 1.54 ;
      RECT  2.0 1.475 2.095 1.56 ;
      RECT  0.49 0.24 0.69 0.36 ;
      RECT  0.6 0.36 0.69 1.225 ;
      RECT  0.54 1.225 1.14 1.315 ;
      RECT  1.05 1.315 1.14 1.54 ;
      RECT  0.54 1.315 0.66 1.625 ;
      RECT  1.05 1.54 1.66 1.65 ;
      RECT  2.0 1.56 2.39 1.66 ;
      LAYER M2 ;
      RECT  0.355 0.55 2.4 0.65 ;
      LAYER V1 ;
      RECT  0.4 0.55 0.5 0.65 ;
      RECT  1.315 0.55 1.415 0.65 ;
      RECT  2.26 0.55 2.36 0.65 ;
  END
END SEN_FDNQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNQ_D_2
#      Description : "D-Flip Flop, neg-edge triggered"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FDNQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.54 0.31 3.66 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.415 0.19 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.8 1.415 0.93 1.75 ;
      RECT  1.785 1.575 1.91 1.75 ;
      RECT  2.79 1.56 2.92 1.75 ;
      RECT  3.275 1.41 3.405 1.75 ;
      RECT  3.8 1.21 3.92 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  3.275 0.05 3.405 0.365 ;
      RECT  0.795 0.05 0.925 0.39 ;
      RECT  1.8 0.05 1.925 0.39 ;
      RECT  2.79 0.05 2.92 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.8 0.05 3.92 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.25 0.185 1.71 0.3 ;
      RECT  1.62 0.3 1.71 0.74 ;
      RECT  1.39 0.74 1.98 0.83 ;
      RECT  1.88 0.63 1.98 0.74 ;
      RECT  1.39 0.83 1.48 1.31 ;
      RECT  1.24 1.31 1.48 1.43 ;
      RECT  2.27 0.22 2.55 0.34 ;
      RECT  2.46 0.34 2.55 0.88 ;
      RECT  2.46 0.88 2.975 0.97 ;
      RECT  2.875 0.97 2.975 1.33 ;
      RECT  2.295 1.33 2.975 1.45 ;
      RECT  1.42 0.39 1.53 0.55 ;
      RECT  1.2 0.55 1.53 0.65 ;
      RECT  1.2 0.65 1.3 0.97 ;
      RECT  3.065 0.39 3.185 0.635 ;
      RECT  2.655 0.635 3.185 0.75 ;
      RECT  3.065 0.75 3.185 0.785 ;
      RECT  3.065 0.785 3.45 0.895 ;
      RECT  3.065 0.895 3.185 1.33 ;
      RECT  0.34 0.505 0.51 0.91 ;
      RECT  0.34 0.91 0.46 1.375 ;
      RECT  2.26 0.485 2.36 1.105 ;
      RECT  2.26 1.105 2.625 1.215 ;
      RECT  1.65 0.92 1.765 1.185 ;
      RECT  1.65 1.185 2.17 1.29 ;
      RECT  2.07 0.24 2.17 1.185 ;
      RECT  1.57 1.385 2.095 1.475 ;
      RECT  1.57 1.475 1.66 1.54 ;
      RECT  2.0 1.475 2.095 1.56 ;
      RECT  0.49 0.24 0.69 0.36 ;
      RECT  0.6 0.36 0.69 1.225 ;
      RECT  0.6 1.225 1.14 1.315 ;
      RECT  0.6 1.315 0.69 1.46 ;
      RECT  1.05 1.315 1.14 1.54 ;
      RECT  0.5 1.46 0.69 1.575 ;
      RECT  1.05 1.54 1.66 1.65 ;
      RECT  2.0 1.56 2.39 1.66 ;
      LAYER M2 ;
      RECT  0.365 0.55 2.4 0.65 ;
      LAYER V1 ;
      RECT  0.405 0.55 0.505 0.65 ;
      RECT  1.32 0.55 1.42 0.65 ;
      RECT  2.26 0.55 2.36 0.65 ;
  END
END SEN_FDNQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNQ_D_4
#      Description : "D-Flip Flop, neg-edge triggered"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FDNQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 4.26 0.69 ;
      RECT  4.15 0.69 4.26 1.105 ;
      RECT  3.55 1.105 4.26 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.8 1.415 0.93 1.75 ;
      RECT  1.785 1.575 1.91 1.75 ;
      RECT  2.8 1.54 2.93 1.75 ;
      RECT  3.34 1.21 3.46 1.75 ;
      RECT  3.875 1.41 4.005 1.75 ;
      RECT  4.4 1.21 4.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.795 0.05 0.925 0.39 ;
      RECT  1.8 0.05 1.925 0.39 ;
      RECT  2.805 0.05 2.935 0.39 ;
      RECT  3.875 0.05 4.005 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.34 0.05 3.46 0.59 ;
      RECT  4.4 0.05 4.52 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.25 0.185 1.71 0.3 ;
      RECT  1.62 0.3 1.71 0.74 ;
      RECT  1.39 0.74 1.98 0.83 ;
      RECT  1.88 0.63 1.98 0.74 ;
      RECT  1.39 0.83 1.48 1.31 ;
      RECT  1.24 1.31 1.48 1.43 ;
      RECT  2.27 0.22 2.55 0.34 ;
      RECT  2.46 0.34 2.55 0.785 ;
      RECT  2.46 0.785 3.0 0.875 ;
      RECT  2.9 0.875 3.0 1.33 ;
      RECT  2.27 1.33 3.0 1.45 ;
      RECT  1.42 0.39 1.53 0.55 ;
      RECT  1.2 0.55 1.53 0.65 ;
      RECT  1.2 0.65 1.3 1.0 ;
      RECT  3.09 0.44 3.21 0.55 ;
      RECT  2.64 0.55 3.21 0.665 ;
      RECT  3.09 0.665 3.21 0.785 ;
      RECT  3.09 0.785 4.06 0.895 ;
      RECT  3.09 0.895 3.21 1.31 ;
      RECT  0.34 0.505 0.51 0.91 ;
      RECT  0.34 0.91 0.46 1.365 ;
      RECT  2.26 0.48 2.36 1.105 ;
      RECT  2.26 1.105 2.63 1.215 ;
      RECT  1.65 0.92 1.765 1.185 ;
      RECT  1.65 1.185 2.17 1.29 ;
      RECT  2.07 0.24 2.17 1.185 ;
      RECT  1.57 1.385 2.095 1.475 ;
      RECT  1.57 1.475 1.66 1.54 ;
      RECT  2.0 1.475 2.095 1.56 ;
      RECT  0.49 0.24 0.69 0.36 ;
      RECT  0.6 0.36 0.69 1.225 ;
      RECT  0.6 1.225 1.14 1.315 ;
      RECT  0.6 1.315 0.69 1.46 ;
      RECT  1.05 1.315 1.14 1.54 ;
      RECT  0.515 1.46 0.69 1.575 ;
      RECT  1.05 1.54 1.66 1.65 ;
      RECT  2.0 1.56 2.39 1.66 ;
      LAYER M2 ;
      RECT  0.365 0.55 2.4 0.65 ;
      LAYER V1 ;
      RECT  0.405 0.55 0.505 0.65 ;
      RECT  1.325 0.55 1.425 0.65 ;
      RECT  2.26 0.55 2.36 0.65 ;
  END
END SEN_FDNQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBQ_1
#      Description : "D-Flip Flop, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBQ_1
  CLASS CORE ;
  FOREIGN SEN_FDNRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.885 ;
      RECT  0.55 0.885 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0588 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.31 5.515 0.49 ;
      RECT  5.35 0.49 5.45 1.11 ;
      RECT  5.35 1.11 5.515 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.65 0.69 ;
      RECT  4.55 0.69 4.65 0.89 ;
      RECT  2.55 0.2 2.65 0.69 ;
      RECT  1.32 0.475 1.42 0.74 ;
      RECT  1.32 0.74 1.52 0.84 ;
      LAYER M2 ;
      RECT  1.25 0.55 4.72 0.65 ;
      LAYER V1 ;
      RECT  4.55 0.55 4.65 0.65 ;
      RECT  2.55 0.55 2.65 0.65 ;
      RECT  1.32 0.55 1.42 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0684 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.615 0.48 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.83 1.615 1.0 1.75 ;
      RECT  2.405 1.615 2.575 1.75 ;
      RECT  2.76 1.615 2.93 1.75 ;
      RECT  3.28 1.615 3.45 1.75 ;
      RECT  4.56 1.61 4.73 1.75 ;
      RECT  5.13 1.44 5.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  1.38 0.05 1.51 0.385 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  2.77 0.05 2.9 0.39 ;
      RECT  4.635 0.05 4.755 0.39 ;
      RECT  3.3 0.05 3.43 0.425 ;
      RECT  5.14 0.05 5.255 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.855 0.24 2.395 0.345 ;
      RECT  1.855 0.345 2.0 0.36 ;
      RECT  2.305 0.345 2.395 0.78 ;
      RECT  1.895 0.36 2.0 1.34 ;
      RECT  2.305 0.78 3.16 0.87 ;
      RECT  2.515 0.87 3.16 0.875 ;
      RECT  2.515 0.875 2.635 1.16 ;
      RECT  0.815 0.275 1.23 0.395 ;
      RECT  1.14 0.395 1.23 0.93 ;
      RECT  1.14 0.93 1.755 1.02 ;
      RECT  1.635 0.255 1.755 0.93 ;
      RECT  1.14 1.02 1.245 1.16 ;
      RECT  1.65 1.02 1.755 1.34 ;
      RECT  3.57 0.285 3.695 0.495 ;
      RECT  3.57 0.495 3.66 0.99 ;
      RECT  3.57 0.99 3.71 1.225 ;
      RECT  3.04 0.195 3.16 0.525 ;
      RECT  3.04 0.525 3.48 0.615 ;
      RECT  3.39 0.615 3.48 1.25 ;
      RECT  2.28 0.96 2.38 1.25 ;
      RECT  2.28 1.25 3.48 1.34 ;
      RECT  0.585 0.18 0.705 0.53 ;
      RECT  0.585 0.53 0.83 0.62 ;
      RECT  0.74 0.62 0.83 1.22 ;
      RECT  0.265 0.975 0.355 1.22 ;
      RECT  0.265 1.22 0.83 1.25 ;
      RECT  0.265 1.25 1.55 1.34 ;
      RECT  1.44 1.11 1.55 1.25 ;
      RECT  3.99 0.17 4.095 0.78 ;
      RECT  3.99 0.78 4.43 0.87 ;
      RECT  4.34 0.87 4.43 1.225 ;
      RECT  3.99 1.225 4.43 1.25 ;
      RECT  3.99 1.25 5.26 1.34 ;
      RECT  5.14 0.715 5.26 1.25 ;
      RECT  3.75 0.615 3.89 0.785 ;
      RECT  3.8 0.785 3.89 1.04 ;
      RECT  3.8 1.04 4.25 1.13 ;
      RECT  4.15 0.96 4.25 1.04 ;
      RECT  3.8 1.13 3.9 1.29 ;
      RECT  4.865 0.19 4.985 0.99 ;
      RECT  4.52 0.99 4.985 1.16 ;
      RECT  2.09 0.52 2.19 1.29 ;
      RECT  0.08 0.3 0.17 1.43 ;
      RECT  0.08 1.43 3.865 1.52 ;
      RECT  3.775 1.52 3.865 1.57 ;
      RECT  1.975 1.52 2.145 1.66 ;
      RECT  3.775 1.57 4.005 1.66 ;
      RECT  4.23 1.43 5.025 1.52 ;
      LAYER M2 ;
      RECT  1.37 1.15 3.97 1.25 ;
      LAYER V1 ;
      RECT  1.445 1.15 1.545 1.25 ;
      RECT  2.09 1.15 2.19 1.25 ;
      RECT  3.8 1.15 3.9 1.25 ;
  END
END SEN_FDNRBQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBQ_2
#      Description : "D-Flip Flop, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBQ_2
  CLASS CORE ;
  FOREIGN SEN_FDNRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.885 ;
      RECT  0.55 0.885 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0492 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.425 7.075 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.06 0.51 6.36 0.69 ;
      RECT  3.25 0.2 3.35 0.69 ;
      RECT  2.15 0.49 2.25 0.67 ;
      RECT  1.58 0.67 2.25 0.78 ;
      LAYER M2 ;
      RECT  2.1 0.55 6.29 0.65 ;
      LAYER V1 ;
      RECT  6.15 0.55 6.25 0.65 ;
      RECT  3.25 0.55 3.35 0.65 ;
      RECT  2.15 0.55 2.25 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.084 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.615 0.48 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  0.83 1.615 1.0 1.75 ;
      RECT  1.37 1.615 1.54 1.75 ;
      RECT  2.75 1.615 2.92 1.75 ;
      RECT  3.43 1.615 3.6 1.75 ;
      RECT  3.97 1.61 4.14 1.75 ;
      RECT  4.505 1.615 4.675 1.75 ;
      RECT  5.99 1.61 6.16 1.75 ;
      RECT  6.69 1.44 6.82 1.75 ;
      RECT  7.215 1.215 7.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  1.6 0.05 1.77 0.325 ;
      RECT  4.47 0.05 4.595 0.365 ;
      RECT  3.95 0.05 4.08 0.37 ;
      RECT  6.115 0.05 6.245 0.385 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  3.44 0.05 3.57 0.39 ;
      RECT  6.695 0.05 6.815 0.59 ;
      RECT  7.215 0.05 7.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.795 0.14 1.485 0.24 ;
      RECT  1.365 0.24 1.485 0.415 ;
      RECT  1.365 0.415 2.055 0.535 ;
      RECT  2.07 0.22 3.085 0.325 ;
      RECT  2.59 0.325 3.085 0.34 ;
      RECT  2.995 0.34 3.085 0.78 ;
      RECT  2.59 0.34 2.68 1.06 ;
      RECT  2.995 0.78 3.695 0.87 ;
      RECT  3.2 0.87 3.29 1.16 ;
      RECT  2.175 1.06 2.68 1.15 ;
      RECT  2.175 1.15 2.295 1.315 ;
      RECT  4.685 0.22 5.955 0.34 ;
      RECT  5.865 0.34 5.955 1.22 ;
      RECT  5.39 1.22 5.955 1.25 ;
      RECT  5.39 1.25 6.8 1.34 ;
      RECT  6.69 0.72 6.8 1.25 ;
      RECT  6.375 0.24 6.57 0.36 ;
      RECT  6.48 0.36 6.57 1.015 ;
      RECT  6.075 0.8 6.185 1.015 ;
      RECT  6.075 1.015 6.57 1.135 ;
      RECT  0.585 0.215 0.705 0.53 ;
      RECT  0.585 0.53 0.83 0.62 ;
      RECT  0.74 0.62 0.83 1.2 ;
      RECT  0.265 0.975 0.355 1.2 ;
      RECT  0.265 1.2 1.83 1.29 ;
      RECT  1.72 1.11 1.83 1.2 ;
      RECT  4.165 0.455 5.165 0.56 ;
      RECT  4.575 0.56 4.665 1.0 ;
      RECT  4.21 1.0 5.085 1.105 ;
      RECT  3.695 0.27 3.815 0.595 ;
      RECT  3.695 0.595 3.875 0.685 ;
      RECT  3.785 0.685 3.875 0.795 ;
      RECT  3.785 0.795 4.485 0.885 ;
      RECT  3.785 0.885 3.875 1.25 ;
      RECT  3.01 1.17 3.11 1.25 ;
      RECT  3.01 1.25 3.875 1.34 ;
      RECT  4.915 0.68 5.265 0.79 ;
      RECT  5.175 0.79 5.265 1.02 ;
      RECT  5.175 1.02 5.775 1.13 ;
      RECT  5.175 1.13 5.265 1.2 ;
      RECT  3.965 1.11 4.065 1.2 ;
      RECT  3.965 1.2 5.265 1.29 ;
      RECT  2.41 0.435 2.5 0.87 ;
      RECT  1.54 0.87 2.5 0.96 ;
      RECT  1.54 0.96 1.63 1.005 ;
      RECT  1.93 0.96 2.035 1.31 ;
      RECT  0.92 0.33 1.25 0.42 ;
      RECT  0.92 0.42 1.01 1.005 ;
      RECT  0.92 1.005 1.63 1.11 ;
      RECT  2.8 0.485 2.9 1.31 ;
      RECT  0.08 0.43 0.17 1.43 ;
      RECT  0.08 1.43 5.1 1.52 ;
      RECT  5.01 1.52 5.1 1.57 ;
      RECT  2.345 1.52 2.455 1.65 ;
      RECT  5.01 1.57 5.44 1.66 ;
      RECT  5.66 1.43 6.6 1.52 ;
      LAYER M2 ;
      RECT  1.685 1.15 4.105 1.25 ;
      LAYER V1 ;
      RECT  1.725 1.15 1.825 1.25 ;
      RECT  2.8 1.15 2.9 1.25 ;
      RECT  3.965 1.15 4.065 1.25 ;
  END
END SEN_FDNRBQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBQ_4
#      Description : "D-Flip Flop, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBQ_4
  CLASS CORE ;
  FOREIGN SEN_FDNRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.47 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0714 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.91 ;
      RECT  1.15 0.91 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1176 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.77 0.465 8.46 0.59 ;
      RECT  8.34 0.59 8.46 1.11 ;
      RECT  7.75 1.11 8.46 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.51 7.25 0.69 ;
      RECT  7.15 0.69 7.25 0.89 ;
      RECT  3.51 0.51 3.85 0.69 ;
      RECT  2.35 0.475 2.49 0.83 ;
      LAYER M2 ;
      RECT  2.28 0.55 7.32 0.65 ;
      LAYER V1 ;
      RECT  7.15 0.55 7.25 0.65 ;
      RECT  3.55 0.55 3.65 0.65 ;
      RECT  2.35 0.55 2.45 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1056 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.59 1.575 0.72 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  1.13 1.575 1.26 1.75 ;
      RECT  1.67 1.575 1.8 1.75 ;
      RECT  3.15 1.63 3.32 1.75 ;
      RECT  3.705 1.61 3.875 1.75 ;
      RECT  4.245 1.615 4.415 1.75 ;
      RECT  4.765 1.615 4.935 1.75 ;
      RECT  5.305 1.615 5.475 1.75 ;
      RECT  6.985 1.615 7.155 1.75 ;
      RECT  7.555 1.44 7.685 1.75 ;
      RECT  8.075 1.41 8.205 1.75 ;
      RECT  8.6 1.215 8.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  4.775 0.05 4.905 0.365 ;
      RECT  5.305 0.05 5.435 0.365 ;
      RECT  8.075 0.05 8.205 0.37 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.58 0.05 0.705 0.39 ;
      RECT  7.055 0.05 7.185 0.39 ;
      RECT  3.635 0.05 3.765 0.4 ;
      RECT  1.9 0.05 2.01 0.405 ;
      RECT  7.56 0.05 7.68 0.59 ;
      RECT  8.6 0.05 8.72 0.59 ;
      RECT  4.26 0.05 4.38 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.12 0.15 1.67 0.24 ;
      RECT  1.57 0.24 1.67 0.29 ;
      RECT  1.12 0.24 1.225 0.43 ;
      RECT  1.57 0.29 1.81 0.41 ;
      RECT  1.72 0.41 1.81 0.495 ;
      RECT  1.72 0.495 2.26 0.585 ;
      RECT  2.145 0.36 2.26 0.495 ;
      RECT  2.43 0.18 2.975 0.255 ;
      RECT  2.43 0.255 3.38 0.27 ;
      RECT  2.885 0.27 3.38 0.375 ;
      RECT  2.43 0.27 2.55 0.385 ;
      RECT  3.29 0.375 3.38 0.79 ;
      RECT  2.885 0.375 2.975 1.235 ;
      RECT  3.29 0.79 3.97 0.895 ;
      RECT  3.46 0.895 3.97 0.9 ;
      RECT  3.46 0.9 3.58 1.16 ;
      RECT  2.05 1.155 2.145 1.235 ;
      RECT  2.05 1.235 2.975 1.34 ;
      RECT  0.795 0.24 1.03 0.36 ;
      RECT  0.94 0.36 1.03 1.185 ;
      RECT  0.355 0.8 0.445 1.185 ;
      RECT  0.355 1.185 1.03 1.215 ;
      RECT  0.355 1.215 1.96 1.305 ;
      RECT  1.86 1.0 1.96 1.215 ;
      RECT  7.305 0.215 7.435 0.385 ;
      RECT  7.345 0.385 7.435 1.015 ;
      RECT  6.945 0.885 7.055 1.015 ;
      RECT  6.945 1.015 7.435 1.135 ;
      RECT  3.955 0.315 4.15 0.435 ;
      RECT  4.06 0.435 4.15 0.79 ;
      RECT  4.06 0.79 5.045 0.9 ;
      RECT  4.06 0.9 4.15 1.25 ;
      RECT  3.255 1.005 3.36 1.25 ;
      RECT  3.255 1.25 4.15 1.34 ;
      RECT  4.47 0.455 6.045 0.575 ;
      RECT  5.135 0.575 5.225 1.015 ;
      RECT  4.47 1.015 6.245 1.12 ;
      RECT  6.14 0.935 6.245 1.015 ;
      RECT  0.325 0.305 0.445 0.6 ;
      RECT  0.175 0.6 0.445 0.69 ;
      RECT  0.175 0.69 0.265 1.395 ;
      RECT  0.175 1.395 1.975 1.45 ;
      RECT  0.175 1.45 5.655 1.485 ;
      RECT  3.065 1.43 5.655 1.45 ;
      RECT  1.885 1.485 5.655 1.52 ;
      RECT  1.885 1.52 3.155 1.54 ;
      RECT  5.565 1.52 5.655 1.57 ;
      RECT  2.715 1.54 2.825 1.65 ;
      RECT  5.565 1.57 6.32 1.66 ;
      RECT  1.315 0.5 1.63 0.62 ;
      RECT  1.54 0.62 1.63 0.82 ;
      RECT  1.54 0.82 2.22 0.91 ;
      RECT  2.13 0.91 2.22 0.92 ;
      RECT  1.54 0.91 1.63 1.02 ;
      RECT  2.13 0.92 2.795 1.01 ;
      RECT  2.69 0.36 2.795 0.92 ;
      RECT  2.285 1.01 2.455 1.14 ;
      RECT  1.355 1.02 1.63 1.125 ;
      RECT  5.815 0.745 6.425 0.845 ;
      RECT  6.335 0.845 6.425 1.055 ;
      RECT  6.335 1.055 6.655 1.145 ;
      RECT  6.545 0.905 6.655 1.055 ;
      RECT  6.335 1.145 6.425 1.21 ;
      RECT  4.24 1.09 4.34 1.21 ;
      RECT  4.24 1.21 6.425 1.3 ;
      RECT  7.555 0.785 8.24 0.895 ;
      RECT  7.555 0.895 7.645 1.235 ;
      RECT  5.57 0.255 6.605 0.365 ;
      RECT  6.515 0.365 6.605 0.63 ;
      RECT  6.515 0.63 6.855 0.72 ;
      RECT  6.765 0.72 6.855 1.235 ;
      RECT  6.515 1.235 7.645 1.325 ;
      RECT  6.515 1.325 6.605 1.39 ;
      RECT  5.82 1.39 6.605 1.48 ;
      RECT  3.065 0.68 3.165 1.29 ;
      RECT  6.695 1.415 7.465 1.52 ;
      LAYER M2 ;
      RECT  1.79 1.15 4.41 1.25 ;
      LAYER V1 ;
      RECT  1.86 1.15 1.96 1.25 ;
      RECT  3.065 1.15 3.165 1.25 ;
      RECT  4.24 1.15 4.34 1.25 ;
  END
END SEN_FDNRBQ_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBQ_D_1
#      Description : "D-Flip Flop, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FDNRBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.31 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.178 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.665 0.9 ;
      RECT  2.115 0.655 2.285 0.98 ;
      LAYER M2 ;
      RECT  2.145 0.75 3.69 0.85 ;
      LAYER V1 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  2.185 0.75 2.285 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.042 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.81 1.495 0.98 1.75 ;
      RECT  1.81 1.63 1.98 1.75 ;
      RECT  2.26 1.63 2.47 1.75 ;
      RECT  3.445 1.28 3.575 1.75 ;
      RECT  4.015 1.41 4.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  3.34 0.05 3.51 0.17 ;
      RECT  0.82 0.05 0.99 0.2 ;
      RECT  2.305 0.05 2.475 0.205 ;
      RECT  4.07 0.05 4.2 0.375 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.155 0.16 2.165 0.25 ;
      RECT  2.075 0.25 2.165 0.295 ;
      RECT  1.155 0.25 1.245 0.3 ;
      RECT  2.075 0.295 3.105 0.385 ;
      RECT  3.005 0.16 3.105 0.295 ;
      RECT  0.575 0.3 1.245 0.39 ;
      RECT  0.575 0.39 0.72 0.485 ;
      RECT  0.63 0.485 0.72 1.0 ;
      RECT  0.575 1.0 0.72 1.2 ;
      RECT  1.48 0.34 1.985 0.445 ;
      RECT  1.895 0.445 1.985 0.475 ;
      RECT  1.895 0.475 2.495 0.565 ;
      RECT  2.39 0.565 2.495 0.84 ;
      RECT  1.895 0.565 1.985 0.875 ;
      RECT  1.41 0.875 1.985 0.965 ;
      RECT  1.41 0.965 1.5 1.235 ;
      RECT  1.32 1.235 1.5 1.355 ;
      RECT  3.235 0.26 3.345 0.495 ;
      RECT  3.235 0.495 4.26 0.615 ;
      RECT  4.145 0.615 4.26 1.175 ;
      RECT  3.71 1.175 4.26 1.265 ;
      RECT  3.71 1.265 3.83 1.5 ;
      RECT  2.585 0.48 2.755 0.6 ;
      RECT  2.585 0.6 2.675 1.07 ;
      RECT  1.78 1.07 2.705 1.16 ;
      RECT  2.6 1.16 2.705 1.33 ;
      RECT  2.845 0.48 3.085 0.6 ;
      RECT  2.98 0.6 3.085 0.995 ;
      RECT  2.98 0.995 3.92 1.085 ;
      RECT  3.81 0.895 3.92 0.995 ;
      RECT  2.98 1.085 3.1 1.46 ;
      RECT  2.765 0.69 2.885 0.87 ;
      RECT  2.795 0.87 2.885 1.45 ;
      RECT  1.695 0.58 1.805 0.695 ;
      RECT  1.14 0.695 1.805 0.785 ;
      RECT  1.14 0.785 1.295 0.935 ;
      RECT  1.14 0.935 1.23 1.31 ;
      RECT  0.34 0.45 0.445 0.725 ;
      RECT  0.34 0.725 0.54 0.905 ;
      RECT  0.34 0.905 0.445 1.31 ;
      RECT  0.34 1.31 1.23 1.4 ;
      RECT  1.14 1.4 1.23 1.45 ;
      RECT  1.14 1.45 2.885 1.54 ;
      RECT  2.795 1.54 2.885 1.55 ;
      RECT  2.795 1.55 3.25 1.64 ;
      RECT  1.59 1.25 2.25 1.355 ;
  END
END SEN_FDNRBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBQ_D_2
#      Description : "D-Flip Flop, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FDNRBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.31 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.665 0.9 ;
      RECT  2.115 0.655 2.285 0.98 ;
      LAYER M2 ;
      RECT  2.145 0.75 3.69 0.85 ;
      LAYER V1 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  2.185 0.75 2.285 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.81 1.495 0.98 1.75 ;
      RECT  1.81 1.63 1.98 1.75 ;
      RECT  2.26 1.63 2.47 1.75 ;
      RECT  3.445 1.28 3.575 1.75 ;
      RECT  4.015 1.4 4.145 1.75 ;
      RECT  4.6 1.21 4.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  3.34 0.05 3.51 0.17 ;
      RECT  0.82 0.05 0.99 0.2 ;
      RECT  2.305 0.05 2.475 0.205 ;
      RECT  4.075 0.05 4.205 0.375 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  4.6 0.05 4.72 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.155 0.16 2.165 0.25 ;
      RECT  2.075 0.25 2.165 0.295 ;
      RECT  1.155 0.25 1.245 0.3 ;
      RECT  2.075 0.295 3.105 0.385 ;
      RECT  3.005 0.16 3.105 0.295 ;
      RECT  0.575 0.3 1.245 0.39 ;
      RECT  0.575 0.39 0.72 0.485 ;
      RECT  0.63 0.485 0.72 1.0 ;
      RECT  0.575 1.0 0.72 1.2 ;
      RECT  1.48 0.34 1.985 0.445 ;
      RECT  1.895 0.445 1.985 0.475 ;
      RECT  1.895 0.475 2.495 0.565 ;
      RECT  2.39 0.565 2.495 0.82 ;
      RECT  1.895 0.565 1.985 0.875 ;
      RECT  1.41 0.875 1.985 0.965 ;
      RECT  1.41 0.965 1.5 1.235 ;
      RECT  1.32 1.235 1.5 1.355 ;
      RECT  3.235 0.26 3.345 0.495 ;
      RECT  3.235 0.495 4.26 0.615 ;
      RECT  4.145 0.615 4.26 1.175 ;
      RECT  3.71 1.175 4.26 1.265 ;
      RECT  3.71 1.265 3.83 1.5 ;
      RECT  2.585 0.48 2.755 0.6 ;
      RECT  2.585 0.6 2.675 1.07 ;
      RECT  1.77 1.07 2.705 1.16 ;
      RECT  2.6 1.16 2.705 1.33 ;
      RECT  2.845 0.48 3.085 0.6 ;
      RECT  2.98 0.6 3.085 0.995 ;
      RECT  2.98 0.995 3.92 1.085 ;
      RECT  3.81 0.745 3.92 0.995 ;
      RECT  2.98 1.085 3.1 1.46 ;
      RECT  2.765 0.69 2.885 0.87 ;
      RECT  2.795 0.87 2.885 1.45 ;
      RECT  1.695 0.58 1.805 0.695 ;
      RECT  1.14 0.695 1.805 0.785 ;
      RECT  1.14 0.785 1.295 0.935 ;
      RECT  1.14 0.935 1.23 1.31 ;
      RECT  0.34 0.45 0.445 0.725 ;
      RECT  0.34 0.725 0.54 0.905 ;
      RECT  0.34 0.905 0.445 1.31 ;
      RECT  0.34 1.31 1.23 1.4 ;
      RECT  1.14 1.4 1.23 1.45 ;
      RECT  1.14 1.45 2.885 1.54 ;
      RECT  2.795 1.54 2.885 1.55 ;
      RECT  2.795 1.55 3.25 1.64 ;
      RECT  1.59 1.25 2.25 1.355 ;
  END
END SEN_FDNRBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBQ_D_4
#      Description : "D-Flip Flop, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FDNRBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.3 0.51 5.05 0.69 ;
      RECT  4.95 0.69 5.05 1.11 ;
      RECT  4.35 1.11 5.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.665 0.9 ;
      RECT  2.115 0.655 2.285 0.98 ;
      LAYER M2 ;
      RECT  2.145 0.75 3.69 0.85 ;
      LAYER V1 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  2.185 0.75 2.285 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  0.79 1.495 1.0 1.75 ;
      RECT  1.81 1.63 1.98 1.75 ;
      RECT  2.26 1.63 2.47 1.75 ;
      RECT  3.445 1.28 3.575 1.75 ;
      RECT  4.02 1.41 4.15 1.75 ;
      RECT  4.595 1.41 4.725 1.75 ;
      RECT  5.15 1.21 5.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  3.34 0.05 3.51 0.17 ;
      RECT  0.82 0.05 0.99 0.2 ;
      RECT  2.305 0.05 2.475 0.205 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  4.075 0.05 4.205 0.39 ;
      RECT  4.595 0.05 4.725 0.39 ;
      RECT  5.15 0.05 5.27 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.155 0.16 2.165 0.25 ;
      RECT  2.075 0.25 2.165 0.295 ;
      RECT  1.155 0.25 1.245 0.3 ;
      RECT  2.075 0.295 3.105 0.385 ;
      RECT  3.005 0.16 3.105 0.295 ;
      RECT  0.575 0.3 1.245 0.39 ;
      RECT  0.575 0.39 0.72 0.485 ;
      RECT  0.63 0.485 0.72 1.0 ;
      RECT  0.575 1.0 0.72 1.2 ;
      RECT  1.48 0.34 1.985 0.445 ;
      RECT  1.895 0.445 1.985 0.475 ;
      RECT  1.895 0.475 2.495 0.565 ;
      RECT  2.39 0.565 2.495 0.84 ;
      RECT  1.895 0.565 1.985 0.875 ;
      RECT  1.41 0.875 1.985 0.965 ;
      RECT  1.41 0.965 1.5 1.235 ;
      RECT  1.32 1.235 1.5 1.355 ;
      RECT  3.235 0.26 3.345 0.495 ;
      RECT  3.235 0.495 4.14 0.615 ;
      RECT  4.05 0.615 4.14 0.785 ;
      RECT  4.05 0.785 4.86 0.895 ;
      RECT  4.05 0.895 4.14 1.175 ;
      RECT  3.71 1.175 4.14 1.265 ;
      RECT  3.71 1.265 3.83 1.5 ;
      RECT  2.585 0.48 2.755 0.6 ;
      RECT  2.585 0.6 2.675 1.07 ;
      RECT  1.78 1.07 2.705 1.16 ;
      RECT  2.6 1.16 2.705 1.33 ;
      RECT  2.845 0.48 3.085 0.6 ;
      RECT  2.98 0.6 3.085 0.995 ;
      RECT  2.98 0.995 3.925 1.085 ;
      RECT  3.815 0.74 3.925 0.995 ;
      RECT  2.98 1.085 3.1 1.46 ;
      RECT  2.765 0.69 2.885 0.87 ;
      RECT  2.795 0.87 2.885 1.45 ;
      RECT  1.695 0.58 1.805 0.695 ;
      RECT  1.14 0.695 1.805 0.785 ;
      RECT  1.14 0.785 1.295 0.935 ;
      RECT  1.14 0.935 1.23 1.31 ;
      RECT  0.34 0.4 0.445 0.725 ;
      RECT  0.34 0.725 0.54 0.905 ;
      RECT  0.34 0.905 0.445 1.31 ;
      RECT  0.34 1.31 1.23 1.4 ;
      RECT  1.14 1.4 1.23 1.45 ;
      RECT  1.14 1.45 2.885 1.54 ;
      RECT  2.795 1.54 2.885 1.55 ;
      RECT  2.795 1.55 3.25 1.64 ;
      RECT  1.59 1.25 2.25 1.355 ;
  END
END SEN_FDNRBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBSBQ_1
#      Description : "D-Flip Flop neg-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBSBQ_1
  CLASS CORE ;
  FOREIGN SEN_FDNRBSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.48 4.85 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0885 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.275 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0387 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.31 5.935 0.49 ;
      RECT  5.75 0.49 5.85 0.995 ;
      RECT  5.75 0.995 5.935 1.18 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.915 0.51 4.05 0.97 ;
      RECT  2.845 0.745 3.145 0.915 ;
      LAYER M2 ;
      RECT  2.965 0.75 4.09 0.85 ;
      LAYER V1 ;
      RECT  3.915 0.75 4.015 0.85 ;
      RECT  3.005 0.75 3.105 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.51 5.51 0.6 ;
      RECT  5.15 0.6 5.25 1.025 ;
      RECT  5.15 1.025 5.39 1.12 ;
      RECT  1.815 0.91 2.08 1.09 ;
      LAYER M2 ;
      RECT  1.79 0.95 5.32 1.05 ;
      LAYER V1 ;
      RECT  5.15 0.95 5.25 1.05 ;
      RECT  1.86 0.95 1.96 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0561 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  3.735 1.24 4.42 1.335 ;
      RECT  3.735 1.335 3.855 1.75 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  1.97 1.44 2.08 1.75 ;
      RECT  2.72 1.39 2.85 1.75 ;
      RECT  5.035 1.41 5.155 1.75 ;
      RECT  5.555 1.4 5.675 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  2.94 0.05 3.07 0.225 ;
      RECT  0.365 0.05 0.495 0.39 ;
      RECT  4.0 0.05 4.13 0.39 ;
      RECT  5.49 0.05 5.62 0.41 ;
      RECT  1.69 0.05 1.82 0.455 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.735 0.21 4.855 0.3 ;
      RECT  4.53 0.3 4.855 0.39 ;
      RECT  4.53 0.39 4.63 1.22 ;
      RECT  4.51 1.22 4.63 1.39 ;
      RECT  0.62 0.265 0.85 0.385 ;
      RECT  0.76 0.385 0.85 1.025 ;
      RECT  0.55 1.025 0.85 1.145 ;
      RECT  1.42 0.225 1.58 0.395 ;
      RECT  1.42 0.395 1.52 1.015 ;
      RECT  1.325 1.015 1.52 1.13 ;
      RECT  4.97 0.22 5.085 0.395 ;
      RECT  4.97 0.395 5.06 1.21 ;
      RECT  4.97 1.21 5.415 1.3 ;
      RECT  5.295 1.3 5.415 1.57 ;
      RECT  2.425 0.315 3.57 0.405 ;
      RECT  2.425 0.405 2.755 0.435 ;
      RECT  3.465 0.405 3.57 0.58 ;
      RECT  2.655 0.435 2.755 1.165 ;
      RECT  2.425 1.165 2.755 1.18 ;
      RECT  2.425 1.18 3.105 1.285 ;
      RECT  2.985 1.285 3.105 1.62 ;
      RECT  3.68 0.24 3.88 0.41 ;
      RECT  3.68 0.41 3.78 0.75 ;
      RECT  3.415 0.75 3.78 0.84 ;
      RECT  3.415 0.84 3.6 0.92 ;
      RECT  3.49 0.92 3.6 1.06 ;
      RECT  3.49 1.06 4.44 1.15 ;
      RECT  4.35 0.95 4.44 1.06 ;
      RECT  3.49 1.15 3.595 1.585 ;
      RECT  0.065 0.26 0.185 0.505 ;
      RECT  0.065 0.505 0.455 0.595 ;
      RECT  0.365 0.595 0.455 1.235 ;
      RECT  0.065 1.235 0.455 1.26 ;
      RECT  0.065 1.26 1.03 1.35 ;
      RECT  0.94 0.22 1.03 1.26 ;
      RECT  0.065 1.35 0.185 1.48 ;
      RECT  3.2 0.495 3.325 0.665 ;
      RECT  3.235 0.665 3.325 1.05 ;
      RECT  3.235 1.05 3.4 1.29 ;
      RECT  2.05 0.62 2.14 0.73 ;
      RECT  1.61 0.73 2.14 0.82 ;
      RECT  1.61 0.82 1.7 1.3 ;
      RECT  1.12 0.225 1.32 0.395 ;
      RECT  1.12 0.395 1.225 1.3 ;
      RECT  1.12 1.3 1.7 1.39 ;
      RECT  2.23 0.3 2.335 0.765 ;
      RECT  2.23 0.765 2.565 0.855 ;
      RECT  2.465 0.855 2.565 0.995 ;
      RECT  2.23 0.855 2.335 1.25 ;
      RECT  1.79 1.25 2.335 1.34 ;
      RECT  1.79 1.34 1.88 1.48 ;
      RECT  1.645 1.48 1.88 1.585 ;
      RECT  0.545 0.51 0.67 0.875 ;
      RECT  5.515 0.75 5.615 1.29 ;
      RECT  4.755 1.215 4.87 1.48 ;
      RECT  3.95 1.48 4.87 1.595 ;
      LAYER M2 ;
      RECT  0.5 0.55 3.85 0.65 ;
      RECT  1.35 0.75 2.795 0.85 ;
      RECT  3.23 1.15 5.69 1.25 ;
      LAYER V1 ;
      RECT  0.57 0.55 0.67 0.65 ;
      RECT  3.68 0.55 3.78 0.65 ;
      RECT  1.42 0.75 1.52 0.85 ;
      RECT  2.655 0.75 2.755 0.85 ;
      RECT  3.3 1.15 3.4 1.25 ;
      RECT  4.53 1.15 4.63 1.25 ;
      RECT  5.515 1.15 5.615 1.25 ;
  END
END SEN_FDNRBSBQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBSBQ_2
#      Description : "D-Flip Flop neg-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBSBQ_2
  CLASS CORE ;
  FOREIGN SEN_FDNRBSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.47 0.51 5.65 0.745 ;
      RECT  5.55 0.745 5.65 0.955 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1131 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.68 0.27 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.3 6.675 0.52 ;
      RECT  6.55 0.52 6.65 1.115 ;
      RECT  6.55 1.115 6.675 1.31 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.695 4.85 0.915 ;
      RECT  2.89 0.69 3.175 0.87 ;
      LAYER M2 ;
      RECT  2.995 0.75 4.82 0.85 ;
      LAYER V1 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  3.035 0.75 3.135 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0822 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.465 6.25 0.555 ;
      RECT  6.15 0.555 6.25 0.69 ;
      RECT  5.95 0.555 6.05 1.13 ;
      RECT  1.825 0.91 2.03 1.145 ;
      LAYER M2 ;
      RECT  1.89 0.95 6.09 1.05 ;
      LAYER V1 ;
      RECT  5.95 0.95 6.05 1.05 ;
      RECT  1.93 0.95 2.03 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0645 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.47 1.285 5.145 1.375 ;
      RECT  4.47 1.375 4.56 1.75 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  1.98 1.44 2.09 1.75 ;
      RECT  2.48 1.41 2.61 1.75 ;
      RECT  3.07 1.435 3.21 1.75 ;
      RECT  5.775 1.4 5.89 1.75 ;
      RECT  6.295 1.39 6.415 1.75 ;
      RECT  6.815 1.21 6.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  2.795 0.05 2.965 0.2 ;
      RECT  0.35 0.05 0.52 0.33 ;
      RECT  6.295 0.05 6.42 0.385 ;
      RECT  4.74 0.05 4.87 0.455 ;
      RECT  1.705 0.05 1.825 0.59 ;
      RECT  6.815 0.05 6.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.16 0.23 3.8 0.29 ;
      RECT  2.49 0.29 3.8 0.325 ;
      RECT  2.49 0.325 3.28 0.38 ;
      RECT  0.625 0.215 0.85 0.335 ;
      RECT  0.76 0.335 0.85 1.025 ;
      RECT  0.545 1.025 0.85 1.145 ;
      RECT  5.74 0.255 5.975 0.365 ;
      RECT  5.74 0.365 5.83 1.04 ;
      RECT  5.7 1.04 5.83 1.22 ;
      RECT  5.7 1.22 6.155 1.31 ;
      RECT  6.035 1.31 6.155 1.61 ;
      RECT  1.4 0.225 1.59 0.395 ;
      RECT  1.4 0.395 1.505 1.16 ;
      RECT  5.28 0.285 5.645 0.405 ;
      RECT  5.28 0.405 5.38 1.255 ;
      RECT  5.235 1.255 5.38 1.43 ;
      RECT  3.89 0.275 4.01 0.415 ;
      RECT  3.695 0.415 4.01 0.505 ;
      RECT  3.695 0.505 3.795 1.43 ;
      RECT  0.065 0.29 0.185 0.42 ;
      RECT  0.065 0.42 0.45 0.51 ;
      RECT  0.36 0.51 0.45 1.26 ;
      RECT  0.065 1.26 1.03 1.35 ;
      RECT  0.94 0.28 1.03 1.26 ;
      RECT  0.065 1.35 0.185 1.49 ;
      RECT  4.485 0.25 4.605 0.425 ;
      RECT  4.345 0.425 4.605 0.515 ;
      RECT  4.345 0.515 4.445 0.78 ;
      RECT  4.095 0.78 4.445 0.87 ;
      RECT  4.095 0.87 4.23 0.95 ;
      RECT  4.14 0.95 4.23 1.085 ;
      RECT  4.14 1.085 5.18 1.175 ;
      RECT  5.01 1.055 5.18 1.085 ;
      RECT  4.15 0.45 4.255 0.595 ;
      RECT  3.915 0.595 4.255 0.685 ;
      RECT  3.915 0.685 4.005 1.2 ;
      RECT  3.915 1.2 4.05 1.52 ;
      RECT  2.48 0.47 3.575 0.56 ;
      RECT  2.48 0.56 2.58 0.89 ;
      RECT  3.485 0.56 3.575 1.225 ;
      RECT  2.695 1.225 3.575 1.345 ;
      RECT  3.42 1.345 3.575 1.52 ;
      RECT  3.42 1.52 4.05 1.61 ;
      RECT  0.54 0.425 0.67 0.79 ;
      RECT  1.62 0.73 2.21 0.82 ;
      RECT  2.12 0.82 2.21 1.17 ;
      RECT  1.62 0.82 1.71 1.315 ;
      RECT  1.12 0.225 1.31 0.395 ;
      RECT  1.12 0.395 1.225 1.315 ;
      RECT  1.12 1.315 1.71 1.405 ;
      RECT  6.225 0.79 6.415 0.89 ;
      RECT  6.315 0.89 6.415 1.29 ;
      RECT  2.3 0.435 2.39 0.995 ;
      RECT  2.3 0.995 3.395 1.085 ;
      RECT  3.305 0.69 3.395 0.995 ;
      RECT  2.3 1.085 2.39 1.26 ;
      RECT  1.8 1.26 2.39 1.35 ;
      RECT  1.8 1.35 1.89 1.495 ;
      RECT  2.225 1.35 2.39 1.53 ;
      RECT  1.63 1.495 1.89 1.6 ;
      RECT  4.69 1.48 4.86 1.52 ;
      RECT  4.69 1.52 5.6 1.61 ;
      RECT  5.495 1.22 5.6 1.52 ;
      LAYER M2 ;
      RECT  0.53 0.55 4.485 0.65 ;
      RECT  1.365 0.75 2.62 0.85 ;
      RECT  3.655 1.15 6.455 1.25 ;
      LAYER V1 ;
      RECT  0.57 0.55 0.67 0.65 ;
      RECT  4.345 0.55 4.445 0.65 ;
      RECT  1.405 0.75 1.505 0.85 ;
      RECT  2.48 0.75 2.58 0.85 ;
      RECT  3.695 1.15 3.795 1.25 ;
      RECT  5.28 1.15 5.38 1.25 ;
      RECT  6.315 1.15 6.415 1.25 ;
  END
END SEN_FDNRBSBQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDNRBSBQ_4
#      Description : "D-Flip Flop neg-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDNRBSBQ_4
  CLASS CORE ;
  FOREIGN SEN_FDNRBSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.495 0.35 6.675 0.72 ;
      RECT  5.485 0.24 5.585 0.66 ;
      LAYER M2 ;
      RECT  5.445 0.35 6.675 0.45 ;
      LAYER V1 ;
      RECT  6.535 0.35 6.635 0.45 ;
      RECT  5.485 0.35 5.585 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1506 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.255 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.56 0.47 8.25 0.59 ;
      RECT  8.15 0.59 8.25 1.11 ;
      RECT  7.59 1.025 7.94 1.11 ;
      RECT  7.59 1.11 8.25 1.145 ;
      RECT  7.85 1.145 8.25 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.635 6.13 0.95 ;
      RECT  5.495 0.75 5.675 1.14 ;
      RECT  3.15 0.75 3.66 0.925 ;
      LAYER M2 ;
      RECT  3.255 0.75 6.14 0.85 ;
      LAYER V1 ;
      RECT  6.0 0.75 6.1 0.85 ;
      RECT  5.535 0.75 5.635 0.85 ;
      RECT  3.295 0.75 3.395 0.85 ;
      RECT  3.52 0.75 3.62 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1143 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.215 0.47 7.305 0.89 ;
      RECT  6.97 0.89 7.305 0.98 ;
      RECT  6.97 0.98 7.075 1.145 ;
      RECT  1.895 0.81 2.31 0.9 ;
      RECT  2.21 0.9 2.31 1.16 ;
      LAYER M2 ;
      RECT  2.17 0.95 7.11 1.05 ;
      LAYER V1 ;
      RECT  6.97 0.95 7.07 1.05 ;
      RECT  2.21 0.95 2.31 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0762 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  5.465 1.27 6.15 1.385 ;
      RECT  5.465 1.385 5.555 1.75 ;
      RECT  0.3 1.475 0.47 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  2.055 1.45 2.175 1.75 ;
      RECT  2.58 1.45 2.71 1.75 ;
      RECT  3.115 1.45 3.245 1.75 ;
      RECT  3.635 1.45 3.765 1.75 ;
      RECT  4.945 1.19 5.055 1.75 ;
      RECT  6.795 1.44 6.925 1.75 ;
      RECT  7.335 1.43 7.465 1.75 ;
      RECT  7.87 1.415 8.0 1.75 ;
      RECT  8.41 1.21 8.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  3.625 0.05 3.755 0.225 ;
      RECT  5.895 0.05 6.065 0.34 ;
      RECT  0.32 0.05 0.43 0.36 ;
      RECT  1.975 0.05 2.105 0.36 ;
      RECT  7.35 0.05 7.48 0.38 ;
      RECT  7.87 0.05 8.0 0.38 ;
      RECT  3.095 0.05 3.22 0.41 ;
      RECT  8.41 0.05 8.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.525 0.14 1.57 0.23 ;
      RECT  0.525 0.23 0.625 0.925 ;
      RECT  6.26 0.14 6.76 0.26 ;
      RECT  6.26 0.26 6.35 1.21 ;
      RECT  6.26 1.21 6.44 1.45 ;
      RECT  2.27 0.2 3.0 0.305 ;
      RECT  2.27 0.305 2.395 0.45 ;
      RECT  1.72 0.3 1.84 0.45 ;
      RECT  1.72 0.45 2.395 0.54 ;
      RECT  4.725 0.19 5.39 0.305 ;
      RECT  5.27 0.305 5.39 0.41 ;
      RECT  4.725 0.305 4.825 0.515 ;
      RECT  2.805 0.515 4.825 0.635 ;
      RECT  2.805 0.635 2.905 0.9 ;
      RECT  4.585 0.635 4.675 1.07 ;
      RECT  3.93 1.07 4.675 1.16 ;
      RECT  3.93 1.16 4.02 1.25 ;
      RECT  2.805 1.25 4.02 1.36 ;
      RECT  3.9 1.36 4.02 1.48 ;
      RECT  3.9 1.48 4.59 1.595 ;
      RECT  3.31 0.315 4.635 0.42 ;
      RECT  0.065 0.32 0.185 0.45 ;
      RECT  0.065 0.45 0.435 0.54 ;
      RECT  0.345 0.54 0.435 1.295 ;
      RECT  0.065 1.295 1.065 1.385 ;
      RECT  0.965 0.41 1.065 1.295 ;
      RECT  0.065 1.385 0.185 1.52 ;
      RECT  0.715 0.33 0.845 0.5 ;
      RECT  0.755 0.5 0.845 1.09 ;
      RECT  0.57 1.09 0.845 1.205 ;
      RECT  4.95 0.415 5.155 0.535 ;
      RECT  4.95 0.535 5.04 0.85 ;
      RECT  4.765 0.85 5.04 0.94 ;
      RECT  4.765 0.94 4.855 1.25 ;
      RECT  4.13 1.25 4.855 1.365 ;
      RECT  4.675 1.365 4.855 1.45 ;
      RECT  1.47 0.34 1.605 0.54 ;
      RECT  1.505 0.54 1.605 1.225 ;
      RECT  5.675 0.235 5.765 0.55 ;
      RECT  5.675 0.55 5.855 0.65 ;
      RECT  5.765 0.65 5.855 1.04 ;
      RECT  5.765 1.04 6.17 1.15 ;
      RECT  6.865 0.2 6.985 0.55 ;
      RECT  6.765 0.55 6.985 0.64 ;
      RECT  6.765 0.64 6.865 0.81 ;
      RECT  6.55 0.81 6.865 0.915 ;
      RECT  6.76 0.915 6.865 1.26 ;
      RECT  6.76 1.26 7.18 1.35 ;
      RECT  7.06 1.35 7.18 1.61 ;
      RECT  5.245 0.51 5.345 0.65 ;
      RECT  5.13 0.65 5.345 0.82 ;
      RECT  5.255 0.82 5.345 1.315 ;
      RECT  5.205 1.315 5.345 1.485 ;
      RECT  1.695 0.63 2.49 0.72 ;
      RECT  2.4 0.72 2.49 1.145 ;
      RECT  1.695 0.72 1.785 1.315 ;
      RECT  1.205 0.35 1.315 1.315 ;
      RECT  1.205 1.315 1.785 1.405 ;
      RECT  3.75 0.75 4.495 0.86 ;
      RECT  3.75 0.86 3.84 1.015 ;
      RECT  2.515 0.415 2.715 0.535 ;
      RECT  2.625 0.535 2.715 1.015 ;
      RECT  2.625 1.015 3.84 1.115 ;
      RECT  2.625 1.115 2.715 1.26 ;
      RECT  1.875 1.26 2.715 1.36 ;
      RECT  1.875 1.36 1.965 1.495 ;
      RECT  1.74 1.495 1.965 1.6 ;
      RECT  7.41 0.785 8.02 0.895 ;
      RECT  7.41 0.895 7.5 1.235 ;
      RECT  7.41 1.235 7.69 1.325 ;
      RECT  7.59 1.325 7.69 1.49 ;
      RECT  5.685 1.49 5.855 1.54 ;
      RECT  5.685 1.54 6.64 1.645 ;
      RECT  6.53 1.21 6.64 1.54 ;
      LAYER M2 ;
      RECT  0.485 0.55 5.855 0.65 ;
      RECT  1.465 0.75 2.945 0.85 ;
      RECT  4.675 1.35 7.73 1.45 ;
      LAYER V1 ;
      RECT  0.525 0.55 0.625 0.65 ;
      RECT  5.245 0.55 5.345 0.65 ;
      RECT  5.715 0.55 5.815 0.65 ;
      RECT  1.505 0.75 1.605 0.85 ;
      RECT  2.805 0.75 2.905 0.85 ;
      RECT  4.715 1.35 4.815 1.45 ;
      RECT  6.3 1.35 6.4 1.45 ;
      RECT  7.59 1.35 7.69 1.45 ;
  END
END SEN_FDNRBSBQ_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPCBQ_1
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&RS)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPCBQ_1
  CLASS CORE ;
  FOREIGN SEN_FDPCBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 5.135 0.69 ;
      RECT  4.75 0.69 4.85 1.11 ;
      RECT  4.75 1.11 5.135 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.065 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END RS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.845 1.63 1.015 1.75 ;
      RECT  1.415 1.63 1.585 1.75 ;
      RECT  2.565 1.63 2.735 1.75 ;
      RECT  3.095 1.63 3.265 1.75 ;
      RECT  4.495 1.41 4.62 1.75 ;
      RECT  4.75 1.41 4.89 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  4.22 0.05 4.35 0.38 ;
      RECT  3.205 0.05 3.335 0.385 ;
      RECT  0.1 0.05 0.23 0.39 ;
      RECT  0.915 0.05 1.045 0.39 ;
      RECT  4.75 0.05 4.88 0.39 ;
      RECT  2.655 0.05 2.785 0.42 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.085 0.21 2.56 0.3 ;
      RECT  2.47 0.3 2.56 0.745 ;
      RECT  2.085 0.3 2.195 1.18 ;
      RECT  2.47 0.745 3.005 0.855 ;
      RECT  1.155 0.24 1.925 0.36 ;
      RECT  1.155 0.36 1.275 1.165 ;
      RECT  1.805 0.36 1.925 1.18 ;
      RECT  3.67 0.24 4.1 0.36 ;
      RECT  4.01 0.36 4.1 0.715 ;
      RECT  4.01 0.715 4.445 0.805 ;
      RECT  4.315 0.805 4.445 0.885 ;
      RECT  4.315 0.885 4.405 1.465 ;
      RECT  3.9 1.465 4.405 1.585 ;
      RECT  4.495 0.18 4.625 0.5 ;
      RECT  4.19 0.5 4.625 0.61 ;
      RECT  4.535 0.61 4.625 0.99 ;
      RECT  4.495 0.99 4.625 1.185 ;
      RECT  2.88 0.475 3.185 0.58 ;
      RECT  3.095 0.58 3.185 0.745 ;
      RECT  3.095 0.745 3.36 0.855 ;
      RECT  3.095 0.855 3.185 1.015 ;
      RECT  2.465 1.015 3.185 1.135 ;
      RECT  0.375 0.285 0.495 0.71 ;
      RECT  0.375 0.71 0.65 0.82 ;
      RECT  0.375 0.82 0.465 1.45 ;
      RECT  0.375 1.45 2.145 1.46 ;
      RECT  0.3 1.46 2.145 1.52 ;
      RECT  0.3 1.52 3.68 1.54 ;
      RECT  2.385 1.45 3.68 1.52 ;
      RECT  0.3 1.54 0.47 1.58 ;
      RECT  2.055 1.54 2.475 1.63 ;
      RECT  3.57 1.54 3.68 1.66 ;
      RECT  3.47 0.395 3.585 1.18 ;
      RECT  3.675 0.67 3.765 1.255 ;
      RECT  3.675 1.255 4.225 1.27 ;
      RECT  4.115 1.145 4.225 1.255 ;
      RECT  0.625 0.185 0.745 0.455 ;
      RECT  0.625 0.455 0.845 0.545 ;
      RECT  0.755 0.545 0.845 1.24 ;
      RECT  0.555 1.24 0.845 1.27 ;
      RECT  0.555 1.27 4.225 1.36 ;
      RECT  2.285 0.41 2.375 1.27 ;
  END
END SEN_FDPCBQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPCBQ_1P5
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&RS)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPCBQ_1P5
  CLASS CORE ;
  FOREIGN SEN_FDPCBQ_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0354 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.465 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.3 5.85 1.315 ;
      RECT  5.75 1.315 5.87 1.5 ;
    END
    ANTENNADIFFAREA 0.164 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END RS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.825 1.615 0.995 1.75 ;
      RECT  1.385 1.615 1.555 1.75 ;
      RECT  2.63 1.615 2.8 1.75 ;
      RECT  3.645 1.615 3.815 1.75 ;
      RECT  5.21 1.41 5.335 1.75 ;
      RECT  5.49 1.21 5.61 1.75 ;
      RECT  6.01 1.21 6.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  3.7 0.05 3.825 0.385 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.845 0.05 0.975 0.39 ;
      RECT  2.64 0.05 2.77 0.39 ;
      RECT  3.18 0.05 3.31 0.39 ;
      RECT  4.96 0.05 5.09 0.39 ;
      RECT  5.475 0.05 5.605 0.39 ;
      RECT  6.01 0.05 6.13 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.02 0.21 2.53 0.3 ;
      RECT  2.44 0.3 2.53 0.745 ;
      RECT  2.02 0.3 2.125 1.16 ;
      RECT  2.44 0.745 3.085 0.855 ;
      RECT  1.14 0.24 1.88 0.36 ;
      RECT  1.14 0.36 1.26 1.16 ;
      RECT  1.76 0.36 1.88 1.16 ;
      RECT  3.915 0.24 4.785 0.36 ;
      RECT  4.695 0.36 4.785 0.745 ;
      RECT  4.695 0.745 5.475 0.855 ;
      RECT  5.025 0.855 5.115 1.455 ;
      RECT  4.62 1.455 5.115 1.575 ;
      RECT  3.445 0.285 3.565 0.49 ;
      RECT  3.445 0.49 4.405 0.58 ;
      RECT  3.99 0.58 4.08 1.025 ;
      RECT  3.375 1.025 4.08 1.04 ;
      RECT  3.375 1.04 4.425 1.145 ;
      RECT  5.22 0.19 5.34 0.525 ;
      RECT  4.875 0.525 5.655 0.615 ;
      RECT  5.565 0.615 5.655 1.005 ;
      RECT  5.22 1.005 5.655 1.095 ;
      RECT  5.22 1.095 5.34 1.225 ;
      RECT  2.86 0.49 3.275 0.61 ;
      RECT  3.185 0.61 3.275 0.755 ;
      RECT  3.185 0.755 3.9 0.845 ;
      RECT  3.185 0.845 3.275 1.02 ;
      RECT  2.465 1.02 3.275 1.14 ;
      RECT  0.34 0.37 0.45 0.73 ;
      RECT  0.34 0.73 0.505 0.9 ;
      RECT  0.34 0.9 0.43 1.435 ;
      RECT  0.34 1.435 4.21 1.525 ;
      RECT  0.34 1.525 0.445 1.615 ;
      RECT  4.12 1.525 4.21 1.64 ;
      RECT  2.235 1.525 2.345 1.66 ;
      RECT  4.25 0.68 4.605 0.79 ;
      RECT  4.515 0.79 4.605 1.255 ;
      RECT  0.595 0.195 0.7 1.255 ;
      RECT  0.595 1.255 4.935 1.345 ;
      RECT  2.215 0.405 2.305 1.255 ;
      RECT  4.835 1.12 4.935 1.255 ;
  END
END SEN_FDPCBQ_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPCBQ_2
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&RS)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPCBQ_2
  CLASS CORE ;
  FOREIGN SEN_FDPCBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0414 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  1.91 0.71 2.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0657 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.31 6.27 0.51 ;
      RECT  6.15 0.51 6.45 0.69 ;
      RECT  6.35 0.69 6.45 1.0 ;
      RECT  6.15 1.0 6.45 1.09 ;
      RECT  6.15 1.09 6.27 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  0.95 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0657 ;
  END RS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.57 0.46 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.87 1.57 1.0 1.75 ;
      RECT  1.41 1.57 1.54 1.75 ;
      RECT  1.95 1.57 2.08 1.75 ;
      RECT  3.135 1.575 3.265 1.75 ;
      RECT  3.95 1.57 4.08 1.75 ;
      RECT  5.63 1.44 5.755 1.75 ;
      RECT  5.885 1.44 6.015 1.75 ;
      RECT  6.415 1.21 6.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.41 0.05 1.54 0.24 ;
      RECT  4.2 0.05 4.325 0.36 ;
      RECT  5.49 0.05 5.62 0.375 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  3.18 0.05 3.29 0.39 ;
      RECT  3.68 0.05 3.81 0.39 ;
      RECT  6.41 0.05 6.54 0.39 ;
      RECT  0.86 0.05 0.99 0.41 ;
      RECT  5.89 0.05 6.01 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.6 0.14 3.065 0.23 ;
      RECT  2.975 0.23 3.065 0.62 ;
      RECT  2.6 0.23 2.69 1.03 ;
      RECT  2.975 0.62 3.375 0.71 ;
      RECT  3.265 0.71 3.375 0.86 ;
      RECT  2.55 1.03 2.72 1.12 ;
      RECT  2.215 0.24 2.45 0.36 ;
      RECT  2.36 0.36 2.45 1.03 ;
      RECT  1.665 0.51 1.785 1.03 ;
      RECT  1.09 1.03 2.45 1.12 ;
      RECT  3.425 0.215 3.555 0.385 ;
      RECT  3.465 0.385 3.555 0.755 ;
      RECT  3.465 0.755 4.12 0.865 ;
      RECT  3.465 0.865 3.555 1.03 ;
      RECT  3.025 0.8 3.115 1.03 ;
      RECT  3.025 1.03 3.555 1.12 ;
      RECT  1.12 0.33 2.11 0.42 ;
      RECT  3.895 0.455 4.895 0.56 ;
      RECT  3.895 0.56 4.445 0.575 ;
      RECT  4.355 0.575 4.445 1.0 ;
      RECT  3.66 1.0 4.445 1.01 ;
      RECT  3.66 1.01 4.955 1.12 ;
      RECT  0.355 0.415 0.445 0.71 ;
      RECT  0.355 0.71 0.515 0.895 ;
      RECT  0.355 0.895 0.445 1.39 ;
      RECT  0.065 1.31 0.185 1.39 ;
      RECT  0.065 1.39 4.39 1.48 ;
      RECT  0.065 1.48 0.185 1.53 ;
      RECT  4.3 1.48 4.39 1.57 ;
      RECT  2.755 1.48 2.865 1.65 ;
      RECT  4.3 1.57 4.89 1.66 ;
      RECT  5.62 0.485 5.745 0.72 ;
      RECT  5.415 0.72 5.745 0.83 ;
      RECT  5.635 0.83 5.745 1.16 ;
      RECT  4.68 0.715 5.135 0.825 ;
      RECT  5.045 0.825 5.135 1.21 ;
      RECT  2.795 0.39 2.885 0.875 ;
      RECT  2.795 0.875 2.935 0.965 ;
      RECT  2.845 0.965 2.935 1.21 ;
      RECT  0.605 0.25 0.725 1.21 ;
      RECT  0.605 1.21 5.36 1.3 ;
      RECT  5.27 1.13 5.36 1.21 ;
      RECT  5.835 0.785 6.235 0.895 ;
      RECT  5.835 0.895 5.925 1.26 ;
      RECT  4.415 0.225 5.315 0.345 ;
      RECT  5.225 0.345 5.315 0.92 ;
      RECT  5.225 0.92 5.54 1.01 ;
      RECT  5.45 1.01 5.54 1.26 ;
      RECT  5.45 1.26 5.925 1.35 ;
      RECT  5.45 1.35 5.54 1.52 ;
      RECT  4.49 1.39 5.21 1.48 ;
      RECT  5.09 1.48 5.21 1.52 ;
      RECT  5.09 1.52 5.54 1.61 ;
  END
END SEN_FDPCBQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPCBQ_3
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&RS)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPCBQ_3
  CLASS CORE ;
  FOREIGN SEN_FDPCBQ_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.575 2.25 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.14 0.31 7.25 0.475 ;
      RECT  6.565 0.475 7.25 0.59 ;
      RECT  7.15 0.59 7.25 1.11 ;
      RECT  6.605 1.11 7.25 1.29 ;
    END
    ANTENNADIFFAREA 0.4 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0804 ;
  END RS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.615 0.545 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  0.915 1.615 1.085 1.75 ;
      RECT  1.475 1.615 1.645 1.75 ;
      RECT  2.04 1.615 2.21 1.75 ;
      RECT  3.235 1.615 3.405 1.75 ;
      RECT  3.775 1.615 3.945 1.75 ;
      RECT  4.315 1.615 4.485 1.75 ;
      RECT  5.995 1.44 6.12 1.75 ;
      RECT  6.345 1.415 6.475 1.75 ;
      RECT  6.865 1.415 6.995 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  3.785 0.05 3.915 0.36 ;
      RECT  1.31 0.05 1.48 0.365 ;
      RECT  4.305 0.05 4.435 0.365 ;
      RECT  6.865 0.05 6.995 0.385 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  5.82 0.05 5.95 0.39 ;
      RECT  0.58 0.05 0.71 0.395 ;
      RECT  3.27 0.05 3.39 0.585 ;
      RECT  6.35 0.05 6.47 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.59 0.2 2.3 0.305 ;
      RECT  1.59 0.305 1.715 0.455 ;
      RECT  1.075 0.3 1.195 0.455 ;
      RECT  1.075 0.455 1.715 0.545 ;
      RECT  2.69 0.215 3.18 0.305 ;
      RECT  3.09 0.305 3.18 0.745 ;
      RECT  2.69 0.305 2.78 1.075 ;
      RECT  3.09 0.745 3.65 0.855 ;
      RECT  2.65 1.075 2.82 1.165 ;
      RECT  1.835 0.395 2.56 0.485 ;
      RECT  1.835 0.485 1.93 1.06 ;
      RECT  2.47 0.485 2.56 1.075 ;
      RECT  1.175 1.06 1.93 1.165 ;
      RECT  2.39 1.075 2.56 1.165 ;
      RECT  4.0 0.455 5.265 0.555 ;
      RECT  4.0 0.555 4.755 0.575 ;
      RECT  4.665 0.575 4.755 1.03 ;
      RECT  4.02 1.03 5.255 1.12 ;
      RECT  5.165 0.89 5.255 1.03 ;
      RECT  3.505 0.45 3.83 0.565 ;
      RECT  3.74 0.565 3.83 0.745 ;
      RECT  3.74 0.745 4.45 0.855 ;
      RECT  3.74 0.855 3.83 1.0 ;
      RECT  3.13 0.95 3.24 1.0 ;
      RECT  3.13 1.0 3.83 1.12 ;
      RECT  6.08 0.215 6.2 0.71 ;
      RECT  6.08 0.71 6.245 0.74 ;
      RECT  5.725 0.74 6.245 0.85 ;
      RECT  6.155 0.85 6.245 1.015 ;
      RECT  6.03 1.015 6.245 1.135 ;
      RECT  5.04 0.645 5.435 0.755 ;
      RECT  5.345 0.755 5.435 1.21 ;
      RECT  2.91 0.415 3.0 1.21 ;
      RECT  2.91 1.21 5.7 1.255 ;
      RECT  0.845 0.31 0.965 0.49 ;
      RECT  0.77 0.49 0.965 0.58 ;
      RECT  0.77 0.58 0.86 1.225 ;
      RECT  0.62 1.225 0.86 1.255 ;
      RECT  0.62 1.255 5.7 1.3 ;
      RECT  0.62 1.3 3.0 1.345 ;
      RECT  5.59 1.3 5.7 1.39 ;
      RECT  6.37 0.785 6.865 0.895 ;
      RECT  6.37 0.895 6.48 1.225 ;
      RECT  4.78 0.225 5.615 0.345 ;
      RECT  5.525 0.345 5.615 0.95 ;
      RECT  5.525 0.95 5.905 1.04 ;
      RECT  5.815 1.04 5.905 1.225 ;
      RECT  5.815 1.225 6.48 1.315 ;
      RECT  5.815 1.315 5.905 1.48 ;
      RECT  4.83 1.39 5.48 1.48 ;
      RECT  5.38 1.48 5.905 1.585 ;
      RECT  0.34 0.26 0.43 0.955 ;
      RECT  0.34 0.955 0.68 1.045 ;
      RECT  0.34 1.045 0.43 1.425 ;
      RECT  0.085 1.425 0.43 1.435 ;
      RECT  0.085 1.435 4.74 1.525 ;
      RECT  4.65 1.525 4.74 1.57 ;
      RECT  2.865 1.525 2.955 1.66 ;
      RECT  4.65 1.57 5.23 1.66 ;
  END
END SEN_FDPCBQ_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPCBQ_4
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&RS)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPCBQ_4
  CLASS CORE ;
  FOREIGN SEN_FDPCBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0585 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.17 0.51 7.86 0.69 ;
      RECT  7.75 0.69 7.86 1.11 ;
      RECT  7.15 1.11 7.86 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END RS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.485 1.57 0.615 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  1.025 1.57 1.155 1.75 ;
      RECT  1.585 1.57 1.715 1.75 ;
      RECT  2.145 1.57 2.275 1.75 ;
      RECT  3.46 1.575 3.59 1.75 ;
      RECT  4.005 1.575 4.135 1.75 ;
      RECT  4.525 1.57 4.655 1.75 ;
      RECT  5.065 1.57 5.195 1.75 ;
      RECT  6.705 1.44 6.835 1.75 ;
      RECT  6.955 1.44 7.085 1.75 ;
      RECT  7.475 1.41 7.605 1.75 ;
      RECT  8.0 1.21 8.12 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  1.365 0.05 1.535 0.185 ;
      RECT  4.495 0.05 4.625 0.385 ;
      RECT  5.015 0.05 5.145 0.385 ;
      RECT  3.465 0.05 3.58 0.39 ;
      RECT  6.375 0.05 6.505 0.39 ;
      RECT  7.475 0.05 7.605 0.39 ;
      RECT  0.08 0.05 0.2 0.59 ;
      RECT  0.61 0.05 0.73 0.59 ;
      RECT  6.96 0.05 7.08 0.59 ;
      RECT  8.0 0.05 8.12 0.59 ;
      RECT  3.985 0.05 4.095 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.43 0.215 3.375 0.305 ;
      RECT  2.895 0.305 3.375 0.335 ;
      RECT  2.43 0.305 2.55 0.385 ;
      RECT  3.285 0.335 3.375 0.735 ;
      RECT  2.895 0.335 2.985 1.015 ;
      RECT  3.285 0.735 3.705 0.845 ;
      RECT  2.68 1.015 2.985 1.12 ;
      RECT  1.08 0.275 2.325 0.38 ;
      RECT  2.7 0.395 2.805 0.475 ;
      RECT  1.655 0.475 2.805 0.575 ;
      RECT  1.655 0.575 1.745 1.015 ;
      RECT  2.42 0.575 2.51 1.015 ;
      RECT  1.26 1.015 2.035 1.12 ;
      RECT  2.42 1.015 2.59 1.12 ;
      RECT  3.66 0.44 3.895 0.56 ;
      RECT  3.805 0.56 3.895 0.745 ;
      RECT  3.805 0.745 5.01 0.855 ;
      RECT  3.805 0.855 3.895 0.975 ;
      RECT  3.3 0.975 3.895 1.095 ;
      RECT  4.185 0.475 5.8 0.59 ;
      RECT  4.185 0.59 5.485 0.595 ;
      RECT  5.395 0.595 5.485 0.97 ;
      RECT  5.395 0.97 5.925 0.99 ;
      RECT  4.21 0.99 5.925 1.11 ;
      RECT  6.69 0.19 6.81 0.695 ;
      RECT  6.38 0.695 6.81 0.805 ;
      RECT  6.69 0.805 6.81 1.16 ;
      RECT  5.62 0.73 6.105 0.84 ;
      RECT  6.015 0.84 6.105 1.21 ;
      RECT  0.87 0.31 0.99 1.18 ;
      RECT  0.71 1.18 0.99 1.21 ;
      RECT  0.71 1.21 6.375 1.3 ;
      RECT  3.08 0.72 3.19 1.21 ;
      RECT  6.9 0.785 7.66 0.895 ;
      RECT  6.9 0.895 6.99 1.25 ;
      RECT  5.32 0.24 6.285 0.36 ;
      RECT  6.195 0.36 6.285 0.925 ;
      RECT  6.195 0.925 6.6 1.035 ;
      RECT  6.51 1.035 6.6 1.25 ;
      RECT  6.51 1.25 6.99 1.35 ;
      RECT  6.51 1.35 6.6 1.39 ;
      RECT  5.505 1.39 6.6 1.48 ;
      RECT  6.075 1.48 6.195 1.63 ;
      RECT  0.345 0.3 0.46 0.945 ;
      RECT  0.345 0.945 0.73 1.055 ;
      RECT  0.345 1.055 0.445 1.39 ;
      RECT  0.17 1.39 5.375 1.48 ;
      RECT  5.285 1.48 5.375 1.57 ;
      RECT  2.84 1.48 2.95 1.66 ;
      RECT  5.285 1.57 5.93 1.66 ;
  END
END SEN_FDPCBQ_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPCBQ_D_1
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&RS)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPCBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FDPCBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.31 4.135 0.49 ;
      RECT  3.95 0.49 4.05 1.11 ;
      RECT  3.95 1.11 4.135 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0297 ;
  END RS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.045 1.595 1.215 1.75 ;
      RECT  2.195 1.605 2.365 1.75 ;
      RECT  3.225 1.455 3.395 1.75 ;
      RECT  3.74 1.21 3.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.53 0.05 0.66 0.22 ;
      RECT  1.035 0.05 1.165 0.22 ;
      RECT  2.25 0.05 2.38 0.39 ;
      RECT  3.235 0.05 3.365 0.39 ;
      RECT  3.74 0.05 3.86 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.065 0.19 0.185 0.32 ;
      RECT  0.065 0.32 1.65 0.41 ;
      RECT  1.53 0.19 1.65 0.32 ;
      RECT  1.765 0.215 2.01 0.335 ;
      RECT  1.92 0.335 2.01 0.535 ;
      RECT  1.92 0.535 2.435 0.625 ;
      RECT  2.335 0.625 2.435 0.84 ;
      RECT  1.92 0.625 2.01 1.215 ;
      RECT  1.765 1.215 2.01 1.335 ;
      RECT  2.72 0.215 2.995 0.335 ;
      RECT  2.905 0.335 2.995 0.865 ;
      RECT  2.905 0.865 3.425 0.965 ;
      RECT  3.325 0.965 3.425 1.275 ;
      RECT  2.775 1.275 3.425 1.365 ;
      RECT  2.775 1.365 2.895 1.47 ;
      RECT  3.51 0.29 3.63 0.665 ;
      RECT  3.11 0.665 3.63 0.755 ;
      RECT  3.11 0.755 3.855 0.77 ;
      RECT  3.515 0.77 3.855 0.925 ;
      RECT  3.515 0.925 3.63 1.47 ;
      RECT  1.72 0.51 1.83 0.975 ;
      RECT  2.715 0.51 2.815 1.085 ;
      RECT  2.715 1.085 3.08 1.185 ;
      RECT  2.135 0.855 2.235 1.14 ;
      RECT  2.135 1.14 2.625 1.26 ;
      RECT  2.525 0.27 2.625 1.14 ;
      RECT  0.74 0.51 0.84 1.17 ;
      RECT  0.325 1.26 0.945 1.35 ;
      RECT  0.855 1.35 0.945 1.41 ;
      RECT  0.325 1.35 0.445 1.63 ;
      RECT  0.855 1.41 1.495 1.5 ;
      RECT  1.325 1.5 1.495 1.66 ;
      RECT  2.005 1.425 2.62 1.515 ;
      RECT  2.005 1.515 2.095 1.55 ;
      RECT  2.53 1.515 2.62 1.56 ;
      RECT  0.93 0.51 1.46 0.6 ;
      RECT  1.34 0.6 1.46 0.755 ;
      RECT  0.93 0.6 1.025 0.955 ;
      RECT  1.34 0.755 1.53 0.925 ;
      RECT  1.34 0.925 1.46 1.15 ;
      RECT  1.34 1.15 1.675 1.24 ;
      RECT  1.585 1.24 1.675 1.55 ;
      RECT  1.585 1.55 2.095 1.65 ;
      RECT  2.53 1.56 2.845 1.66 ;
      LAYER M2 ;
      RECT  0.7 0.55 2.855 0.65 ;
      LAYER V1 ;
      RECT  0.74 0.55 0.84 0.65 ;
      RECT  1.725 0.55 1.825 0.65 ;
      RECT  2.715 0.55 2.815 0.65 ;
  END
END SEN_FDPCBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPCBQ_D_2
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&RS)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPCBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FDPCBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.31 4.085 0.49 ;
      RECT  3.95 0.49 4.05 1.31 ;
      RECT  3.95 1.31 4.085 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0297 ;
  END RS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.045 1.595 1.215 1.75 ;
      RECT  2.195 1.605 2.365 1.75 ;
      RECT  3.225 1.455 3.395 1.75 ;
      RECT  3.7 1.41 3.83 1.75 ;
      RECT  4.22 1.41 4.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.53 0.05 0.66 0.22 ;
      RECT  1.035 0.05 1.165 0.22 ;
      RECT  3.7 0.05 3.83 0.37 ;
      RECT  2.25 0.05 2.38 0.39 ;
      RECT  4.22 0.05 4.345 0.39 ;
      RECT  3.25 0.05 3.37 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.065 0.19 0.185 0.32 ;
      RECT  0.065 0.32 1.65 0.41 ;
      RECT  1.53 0.19 1.65 0.32 ;
      RECT  1.765 0.215 2.01 0.335 ;
      RECT  1.92 0.335 2.01 0.535 ;
      RECT  1.92 0.535 2.435 0.625 ;
      RECT  2.335 0.625 2.435 0.84 ;
      RECT  1.92 0.625 2.01 1.215 ;
      RECT  1.765 1.215 2.01 1.335 ;
      RECT  2.725 0.215 2.995 0.335 ;
      RECT  2.905 0.335 2.995 0.865 ;
      RECT  2.905 0.865 3.425 0.965 ;
      RECT  3.325 0.965 3.425 1.275 ;
      RECT  2.775 1.275 3.425 1.365 ;
      RECT  2.775 1.365 2.895 1.47 ;
      RECT  3.52 0.465 3.64 0.665 ;
      RECT  3.11 0.665 3.64 0.77 ;
      RECT  3.515 0.77 3.64 0.785 ;
      RECT  3.515 0.785 3.86 0.895 ;
      RECT  3.515 0.895 3.63 1.35 ;
      RECT  1.72 0.51 1.83 0.975 ;
      RECT  2.715 0.51 2.815 1.085 ;
      RECT  2.715 1.085 3.08 1.185 ;
      RECT  2.135 0.855 2.235 1.14 ;
      RECT  2.135 1.14 2.625 1.26 ;
      RECT  2.525 0.21 2.625 1.14 ;
      RECT  0.74 0.51 0.84 1.17 ;
      RECT  0.325 1.26 0.945 1.35 ;
      RECT  0.855 1.35 0.945 1.41 ;
      RECT  0.325 1.35 0.445 1.63 ;
      RECT  0.855 1.41 1.495 1.5 ;
      RECT  1.325 1.5 1.495 1.66 ;
      RECT  2.005 1.425 2.62 1.515 ;
      RECT  2.005 1.515 2.095 1.55 ;
      RECT  2.53 1.515 2.62 1.56 ;
      RECT  0.93 0.51 1.46 0.6 ;
      RECT  1.34 0.6 1.46 0.755 ;
      RECT  0.93 0.6 1.025 0.955 ;
      RECT  1.34 0.755 1.53 0.925 ;
      RECT  1.34 0.925 1.46 1.15 ;
      RECT  1.34 1.15 1.675 1.24 ;
      RECT  1.585 1.24 1.675 1.55 ;
      RECT  1.585 1.55 2.095 1.65 ;
      RECT  2.53 1.56 2.845 1.66 ;
      LAYER M2 ;
      RECT  0.7 0.55 2.855 0.65 ;
      LAYER V1 ;
      RECT  0.74 0.55 0.84 0.65 ;
      RECT  1.725 0.55 1.825 0.65 ;
      RECT  2.715 0.55 2.815 0.65 ;
  END
END SEN_FDPCBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPCBQ_D_4
#      Description : "D-Flip Flop, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&RS)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPCBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FDPCBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.02 0.51 4.65 0.69 ;
      RECT  4.55 0.69 4.65 1.11 ;
      RECT  4.02 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0297 ;
  END RS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.045 1.595 1.215 1.75 ;
      RECT  2.195 1.605 2.365 1.75 ;
      RECT  3.225 1.455 3.395 1.75 ;
      RECT  3.76 1.21 3.88 1.75 ;
      RECT  4.275 1.41 4.405 1.75 ;
      RECT  4.8 1.21 4.92 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.53 0.05 0.66 0.22 ;
      RECT  1.035 0.05 1.165 0.22 ;
      RECT  2.25 0.05 2.38 0.385 ;
      RECT  3.245 0.05 3.375 0.39 ;
      RECT  4.275 0.05 4.405 0.39 ;
      RECT  3.76 0.05 3.88 0.59 ;
      RECT  4.8 0.05 4.92 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.065 0.19 0.185 0.32 ;
      RECT  0.065 0.32 1.65 0.41 ;
      RECT  1.53 0.19 1.65 0.32 ;
      RECT  1.765 0.215 2.01 0.335 ;
      RECT  1.92 0.335 2.01 0.535 ;
      RECT  1.92 0.535 2.435 0.625 ;
      RECT  2.335 0.625 2.435 0.84 ;
      RECT  1.92 0.625 2.01 1.215 ;
      RECT  1.765 1.215 2.01 1.335 ;
      RECT  2.73 0.215 2.995 0.335 ;
      RECT  2.905 0.335 2.995 0.78 ;
      RECT  2.905 0.78 3.425 0.88 ;
      RECT  3.325 0.88 3.425 1.275 ;
      RECT  2.775 1.275 3.425 1.365 ;
      RECT  2.775 1.365 2.895 1.47 ;
      RECT  3.115 0.5 3.63 0.605 ;
      RECT  3.115 0.605 3.225 0.69 ;
      RECT  3.515 0.605 3.63 0.785 ;
      RECT  3.515 0.785 4.45 0.895 ;
      RECT  3.515 0.895 3.63 1.26 ;
      RECT  1.72 0.51 1.83 0.975 ;
      RECT  2.715 0.51 2.815 1.085 ;
      RECT  2.715 1.085 3.08 1.185 ;
      RECT  2.135 0.855 2.235 1.14 ;
      RECT  2.135 1.14 2.625 1.26 ;
      RECT  2.525 0.21 2.625 1.14 ;
      RECT  0.74 0.51 0.84 1.17 ;
      RECT  0.325 1.26 0.945 1.35 ;
      RECT  0.855 1.35 0.945 1.41 ;
      RECT  0.325 1.35 0.445 1.62 ;
      RECT  0.855 1.41 1.495 1.5 ;
      RECT  1.325 1.5 1.495 1.66 ;
      RECT  2.005 1.425 2.62 1.515 ;
      RECT  2.005 1.515 2.095 1.55 ;
      RECT  2.53 1.515 2.62 1.56 ;
      RECT  0.93 0.51 1.46 0.6 ;
      RECT  1.34 0.6 1.46 0.755 ;
      RECT  0.93 0.6 1.025 0.955 ;
      RECT  1.34 0.755 1.53 0.925 ;
      RECT  1.34 0.925 1.46 1.15 ;
      RECT  1.34 1.15 1.675 1.24 ;
      RECT  1.585 1.24 1.675 1.55 ;
      RECT  1.585 1.55 2.095 1.65 ;
      RECT  2.53 1.56 2.845 1.66 ;
      LAYER M2 ;
      RECT  0.7 0.55 2.855 0.65 ;
      LAYER V1 ;
      RECT  0.74 0.55 0.84 0.65 ;
      RECT  1.725 0.55 1.825 0.65 ;
      RECT  2.715 0.55 2.815 0.65 ;
  END
END SEN_FDPCBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPHQ_D_2
#      Description : "D-Flip Flop, pos-edge triggered, sync hold, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D&!EN)|(iq&EN)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPHQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FDPHQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.645 0.51 1.85 0.865 ;
      RECT  1.55 0.865 1.85 0.92 ;
      RECT  1.55 0.92 1.735 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0498 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.6 0.85 0.725 ;
      RECT  0.75 0.725 0.9 1.065 ;
      RECT  0.75 1.065 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.4 1.125 0.49 ;
      RECT  0.35 0.49 0.45 0.715 ;
      RECT  1.035 0.49 1.125 0.795 ;
      RECT  0.265 0.715 0.45 0.955 ;
      RECT  0.35 0.955 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0747 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.31 5.475 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.58 0.495 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  1.665 1.61 1.835 1.75 ;
      RECT  1.925 1.61 2.095 1.75 ;
      RECT  3.42 1.6 3.59 1.75 ;
      RECT  4.655 1.16 4.765 1.75 ;
      RECT  5.095 1.41 5.215 1.75 ;
      RECT  5.615 1.21 5.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  2.095 0.05 2.215 0.245 ;
      RECT  0.325 0.05 0.495 0.31 ;
      RECT  5.09 0.05 5.22 0.36 ;
      RECT  1.645 0.05 1.775 0.39 ;
      RECT  4.645 0.05 4.775 0.39 ;
      RECT  3.36 0.05 3.49 0.56 ;
      RECT  5.615 0.05 5.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.95 0.235 4.315 0.335 ;
      RECT  4.225 0.335 4.315 0.8 ;
      RECT  4.09 0.8 4.315 0.9 ;
      RECT  4.09 0.9 4.19 1.54 ;
      RECT  4.09 1.54 4.315 1.65 ;
      RECT  2.575 0.18 2.695 0.34 ;
      RECT  2.24 0.34 2.695 0.43 ;
      RECT  2.24 0.43 2.33 1.4 ;
      RECT  0.84 0.205 1.32 0.31 ;
      RECT  1.23 0.31 1.32 1.175 ;
      RECT  0.99 1.175 1.45 1.285 ;
      RECT  1.36 1.285 1.45 1.4 ;
      RECT  1.36 1.4 2.33 1.49 ;
      RECT  2.24 1.49 2.64 1.58 ;
      RECT  2.55 1.58 2.64 1.66 ;
      RECT  2.845 0.215 3.02 0.39 ;
      RECT  2.93 0.39 3.02 0.74 ;
      RECT  2.93 0.74 3.585 0.84 ;
      RECT  3.475 0.84 3.585 0.99 ;
      RECT  2.93 0.84 3.02 1.47 ;
      RECT  4.405 0.175 4.535 0.535 ;
      RECT  4.405 0.535 4.495 1.095 ;
      RECT  4.335 1.095 4.495 1.28 ;
      RECT  3.635 0.405 3.82 0.595 ;
      RECT  3.71 0.595 3.82 1.11 ;
      RECT  3.205 1.11 3.82 1.2 ;
      RECT  3.715 1.2 3.82 1.29 ;
      RECT  3.91 0.435 4.135 0.645 ;
      RECT  3.91 0.645 4.0 1.4 ;
      RECT  3.13 1.4 4.0 1.49 ;
      RECT  3.13 1.49 3.225 1.57 ;
      RECT  3.83 1.49 4.0 1.64 ;
      RECT  2.7 0.535 2.82 0.745 ;
      RECT  2.73 0.745 2.82 1.57 ;
      RECT  2.73 1.57 3.225 1.66 ;
      RECT  1.94 0.45 2.13 0.66 ;
      RECT  2.025 0.66 2.13 1.02 ;
      RECT  1.915 1.02 2.13 1.215 ;
      RECT  4.915 0.44 5.02 0.725 ;
      RECT  4.585 0.725 5.02 0.785 ;
      RECT  4.585 0.785 5.26 0.83 ;
      RECT  4.92 0.83 5.26 0.895 ;
      RECT  4.585 0.83 4.69 0.9 ;
      RECT  4.92 0.895 5.04 1.33 ;
      RECT  1.435 0.2 1.535 0.77 ;
      RECT  2.435 0.525 2.58 1.265 ;
      RECT  0.065 0.165 0.17 1.4 ;
      RECT  0.065 1.4 0.98 1.49 ;
      RECT  0.54 0.6 0.63 1.4 ;
      RECT  0.89 1.49 0.98 1.57 ;
      RECT  0.065 1.49 0.185 1.62 ;
      RECT  0.89 1.57 1.3 1.66 ;
      LAYER M2 ;
      RECT  1.34 0.35 4.64 0.45 ;
      LAYER V1 ;
      RECT  1.435 0.35 1.535 0.45 ;
      RECT  4.42 0.35 4.52 0.45 ;
  END
END SEN_FDPHQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPHRBSBQ_2
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear/set, sync hold, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(iq&EN)|(!EN&D),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPHRBSBQ_2
  CLASS CORE ;
  FOREIGN SEN_FDPHRBSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.085 0.91 6.25 1.265 ;
      RECT  5.15 0.71 5.45 0.89 ;
      RECT  5.35 0.89 5.45 1.09 ;
      LAYER M2 ;
      RECT  5.31 0.95 6.225 1.05 ;
      LAYER V1 ;
      RECT  6.085 0.95 6.185 1.05 ;
      RECT  5.35 0.95 5.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1011 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.26 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1029 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.31 7.875 0.53 ;
      RECT  7.75 0.53 7.85 1.065 ;
      RECT  7.75 1.065 7.875 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.545 0.87 6.645 1.29 ;
      RECT  3.565 1.125 3.915 1.25 ;
      LAYER M2 ;
      RECT  3.735 1.15 6.685 1.25 ;
      LAYER V1 ;
      RECT  6.545 1.15 6.645 1.25 ;
      RECT  3.775 1.15 3.875 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0786 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.505 7.05 0.865 ;
      RECT  6.915 0.865 7.05 1.035 ;
      RECT  3.855 0.51 4.065 0.855 ;
      LAYER M2 ;
      RECT  3.925 0.55 7.09 0.65 ;
      LAYER V1 ;
      RECT  6.95 0.55 7.05 0.65 ;
      RECT  3.965 0.55 4.065 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.57 1.425 0.68 1.75 ;
      RECT  1.63 1.21 1.72 1.75 ;
      RECT  3.24 1.535 3.37 1.75 ;
      RECT  3.78 1.535 3.91 1.75 ;
      RECT  4.31 1.48 4.48 1.75 ;
      RECT  5.15 1.455 5.275 1.75 ;
      RECT  6.43 1.605 6.6 1.75 ;
      RECT  6.965 1.415 7.09 1.75 ;
      RECT  7.495 1.21 7.615 1.75 ;
      RECT  8.015 1.21 8.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  6.73 0.05 6.86 0.235 ;
      RECT  3.25 0.05 3.38 0.36 ;
      RECT  3.785 0.05 3.915 0.36 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  4.88 0.05 5.01 0.39 ;
      RECT  1.35 0.05 1.48 0.41 ;
      RECT  7.495 0.05 7.615 0.59 ;
      RECT  8.015 0.05 8.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.575 0.17 1.16 0.26 ;
      RECT  0.575 0.26 0.695 0.36 ;
      RECT  1.07 0.26 1.16 0.515 ;
      RECT  1.07 0.515 1.72 0.605 ;
      RECT  1.615 0.38 1.72 0.515 ;
      RECT  7.05 0.175 7.35 0.285 ;
      RECT  7.05 0.285 7.14 0.325 ;
      RECT  5.405 0.14 6.535 0.23 ;
      RECT  6.445 0.23 6.535 0.325 ;
      RECT  5.905 0.23 6.045 0.42 ;
      RECT  5.405 0.23 5.525 0.47 ;
      RECT  6.445 0.325 7.14 0.415 ;
      RECT  5.905 0.42 5.995 1.365 ;
      RECT  5.905 1.365 6.045 1.465 ;
      RECT  5.365 1.465 6.045 1.585 ;
      RECT  0.325 0.2 0.46 0.39 ;
      RECT  0.36 0.39 0.46 1.285 ;
      RECT  0.325 1.285 0.46 1.515 ;
      RECT  4.57 0.235 4.745 0.405 ;
      RECT  4.57 0.405 4.67 1.04 ;
      RECT  4.57 1.04 4.71 1.21 ;
      RECT  6.135 0.32 6.355 0.435 ;
      RECT  6.135 0.435 6.225 0.73 ;
      RECT  6.135 0.73 6.43 0.82 ;
      RECT  6.34 0.82 6.43 1.405 ;
      RECT  6.135 1.405 6.875 1.515 ;
      RECT  0.8 0.35 0.98 0.465 ;
      RECT  0.57 0.465 0.98 0.585 ;
      RECT  0.57 0.585 0.66 1.215 ;
      RECT  0.57 1.215 0.86 1.305 ;
      RECT  0.77 1.305 0.86 1.44 ;
      RECT  0.77 1.44 1.265 1.56 ;
      RECT  1.81 0.31 2.015 0.49 ;
      RECT  1.81 0.49 1.9 1.4 ;
      RECT  1.81 1.4 2.61 1.49 ;
      RECT  5.145 0.37 5.265 0.5 ;
      RECT  4.9 0.5 5.265 0.59 ;
      RECT  4.9 0.59 5.005 0.71 ;
      RECT  4.76 0.71 5.005 0.955 ;
      RECT  4.885 0.955 5.005 1.175 ;
      RECT  2.685 0.45 3.68 0.54 ;
      RECT  6.315 0.55 6.825 0.64 ;
      RECT  6.735 0.64 6.825 1.125 ;
      RECT  6.735 1.125 7.33 1.215 ;
      RECT  7.23 0.435 7.33 1.125 ;
      RECT  7.23 1.215 7.33 1.61 ;
      RECT  4.155 0.265 4.255 0.73 ;
      RECT  4.155 0.73 4.285 0.8 ;
      RECT  4.195 0.8 4.285 0.94 ;
      RECT  1.14 0.71 1.305 0.925 ;
      RECT  1.14 0.925 1.235 1.07 ;
      RECT  3.145 0.8 3.235 0.945 ;
      RECT  3.145 0.945 4.095 1.035 ;
      RECT  4.005 1.035 4.095 1.065 ;
      RECT  4.005 1.065 4.48 1.185 ;
      RECT  4.39 0.215 4.48 1.065 ;
      RECT  2.615 0.85 2.86 1.09 ;
      RECT  1.99 0.69 2.09 1.13 ;
      RECT  2.18 0.2 2.28 1.185 ;
      RECT  2.18 1.185 2.85 1.275 ;
      RECT  5.665 0.34 5.785 1.275 ;
      RECT  4.88 1.275 5.785 1.3 ;
      RECT  4.01 1.3 5.785 1.34 ;
      RECT  2.41 0.215 3.16 0.335 ;
      RECT  2.41 0.335 2.5 0.67 ;
      RECT  2.41 0.67 3.04 0.76 ;
      RECT  2.95 0.76 3.04 1.34 ;
      RECT  2.95 1.34 5.785 1.365 ;
      RECT  2.95 1.365 4.945 1.39 ;
      RECT  2.95 1.39 4.085 1.43 ;
      RECT  2.95 1.43 3.62 1.445 ;
      RECT  3.53 1.445 3.62 1.55 ;
      RECT  1.44 0.72 1.54 1.51 ;
      LAYER M2 ;
      RECT  0.8 0.35 1.95 0.45 ;
      RECT  2.14 0.35 4.295 0.45 ;
      RECT  0.32 0.75 1.28 0.85 ;
      RECT  1.95 0.75 4.9 0.85 ;
      RECT  2.72 0.95 4.71 1.05 ;
      RECT  1.4 1.35 7.37 1.45 ;
      LAYER V1 ;
      RECT  0.84 0.35 0.94 0.45 ;
      RECT  1.81 0.35 1.91 0.45 ;
      RECT  2.18 0.35 2.28 0.45 ;
      RECT  4.155 0.35 4.255 0.45 ;
      RECT  0.36 0.75 0.46 0.85 ;
      RECT  1.14 0.75 1.24 0.85 ;
      RECT  1.99 0.75 2.09 0.85 ;
      RECT  4.76 0.75 4.86 0.85 ;
      RECT  2.76 0.95 2.86 1.05 ;
      RECT  4.57 0.95 4.67 1.05 ;
      RECT  1.44 1.35 1.54 1.45 ;
      RECT  7.23 1.35 7.33 1.45 ;
  END
END SEN_FDPHRBSBQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPMQ_D_1
#      Description : "D-Flip Flop, pos-edge triggered, 2-to-1 muxed data inputs, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D0&!S)|(D1&S)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPMQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FDPMQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.585 0.7 2.05 0.9 ;
      RECT  1.55 0.9 2.05 0.935 ;
      RECT  1.55 0.935 1.69 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.1 ;
      RECT  0.55 1.1 0.85 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.12 0.5 1.25 0.9 ;
      RECT  1.12 0.9 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.31 5.335 0.485 ;
      RECT  5.15 0.485 5.25 1.115 ;
      RECT  5.15 1.115 5.335 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.71 0.16 1.29 0.25 ;
      RECT  0.71 0.25 0.8 0.3 ;
      RECT  1.2 0.25 1.29 0.3 ;
      RECT  0.55 0.3 0.8 0.39 ;
      RECT  1.2 0.3 1.465 0.39 ;
      RECT  0.55 0.39 0.65 0.89 ;
      RECT  1.35 0.39 1.465 0.79 ;
      RECT  0.275 0.89 0.65 0.99 ;
      RECT  0.275 0.99 0.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0747 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.61 0.48 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  1.93 1.6 2.14 1.75 ;
      RECT  3.285 1.51 3.455 1.75 ;
      RECT  4.395 1.565 4.565 1.75 ;
      RECT  4.955 1.21 5.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  1.445 0.05 1.615 0.19 ;
      RECT  3.32 0.05 3.49 0.33 ;
      RECT  0.33 0.05 0.46 0.39 ;
      RECT  1.975 0.05 2.105 0.39 ;
      RECT  4.405 0.05 4.535 0.39 ;
      RECT  4.925 0.05 5.045 0.565 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.575 0.22 2.69 0.41 ;
      RECT  2.6 0.41 2.69 1.175 ;
      RECT  2.57 1.175 2.69 1.295 ;
      RECT  0.94 0.36 1.03 1.295 ;
      RECT  0.94 1.295 2.69 1.385 ;
      RECT  2.78 0.205 2.945 0.44 ;
      RECT  2.78 0.44 3.525 0.53 ;
      RECT  3.435 0.53 3.525 0.81 ;
      RECT  2.78 0.53 2.87 1.13 ;
      RECT  2.78 1.13 2.93 1.305 ;
      RECT  1.725 0.37 1.845 0.5 ;
      RECT  1.725 0.5 2.24 0.59 ;
      RECT  2.15 0.59 2.24 1.1 ;
      RECT  1.78 1.03 1.885 1.1 ;
      RECT  1.78 1.1 2.24 1.2 ;
      RECT  0.065 0.18 0.185 0.63 ;
      RECT  0.065 0.63 0.45 0.74 ;
      RECT  0.065 0.74 0.165 1.41 ;
      RECT  0.065 1.41 0.85 1.495 ;
      RECT  0.065 1.495 1.83 1.5 ;
      RECT  0.75 1.5 1.83 1.6 ;
      RECT  0.065 1.5 0.185 1.62 ;
      RECT  4.675 0.26 4.795 0.63 ;
      RECT  4.34 0.63 4.855 0.72 ;
      RECT  4.765 0.72 4.855 0.795 ;
      RECT  4.34 0.72 4.43 0.885 ;
      RECT  4.765 0.795 5.06 0.885 ;
      RECT  4.765 0.885 4.855 1.41 ;
      RECT  4.71 1.41 4.855 1.6 ;
      RECT  2.33 0.42 2.42 0.755 ;
      RECT  2.33 0.755 2.51 0.925 ;
      RECT  2.33 0.925 2.42 1.185 ;
      RECT  2.96 0.665 3.11 0.84 ;
      RECT  3.02 0.84 3.11 1.31 ;
      RECT  3.02 1.31 3.89 1.4 ;
      RECT  3.8 0.535 3.89 1.31 ;
      RECT  3.75 1.4 3.89 1.565 ;
      RECT  3.75 1.565 4.245 1.66 ;
      RECT  4.53 0.855 4.675 1.025 ;
      RECT  4.53 1.025 4.62 1.365 ;
      RECT  3.84 0.23 4.07 0.35 ;
      RECT  3.98 0.35 4.07 1.365 ;
      RECT  3.98 1.365 4.62 1.455 ;
      RECT  3.2 0.64 3.3 1.09 ;
      RECT  3.2 1.09 3.71 1.19 ;
      RECT  3.62 0.2 3.71 1.09 ;
      RECT  4.16 0.2 4.25 1.11 ;
      RECT  4.16 1.11 4.38 1.23 ;
  END
END SEN_FDPMQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQ_1
#      Description : "D-Flip Flop, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQ_1
  CLASS CORE ;
  FOREIGN SEN_FDPQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.425 0.825 3.525 1.35 ;
      RECT  2.805 0.765 2.945 1.105 ;
      RECT  0.535 0.85 0.625 0.95 ;
      RECT  0.44 0.95 0.625 0.99 ;
      RECT  0.305 0.99 0.625 1.08 ;
      LAYER M2 ;
      RECT  0.44 0.95 3.565 1.05 ;
      LAYER V1 ;
      RECT  3.425 0.95 3.525 1.05 ;
      RECT  2.83 0.95 2.93 1.05 ;
      RECT  0.48 0.95 0.58 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0756 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.92 0.51 1.05 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.31 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.57 0.2 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.765 1.59 0.94 1.75 ;
      RECT  1.805 1.45 1.975 1.75 ;
      RECT  2.305 1.44 2.475 1.75 ;
      RECT  3.795 1.405 3.9 1.75 ;
      RECT  4.065 1.185 4.185 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.475 0.05 2.645 0.355 ;
      RECT  0.8 0.05 0.935 0.36 ;
      RECT  3.475 0.05 3.61 0.36 ;
      RECT  2.0 0.05 2.14 0.47 ;
      RECT  0.31 0.05 0.485 0.58 ;
      RECT  4.065 0.05 4.185 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.98 0.215 3.335 0.335 ;
      RECT  3.245 0.335 3.335 0.47 ;
      RECT  3.245 0.47 3.705 0.56 ;
      RECT  3.615 0.56 3.705 0.73 ;
      RECT  3.615 0.73 3.795 0.9 ;
      RECT  3.615 0.9 3.705 1.465 ;
      RECT  3.24 1.465 3.705 1.585 ;
      RECT  1.035 0.225 1.23 0.345 ;
      RECT  1.14 0.345 1.23 0.99 ;
      RECT  1.015 0.99 1.23 1.105 ;
      RECT  3.7 0.21 3.885 0.38 ;
      RECT  3.795 0.38 3.885 0.42 ;
      RECT  3.795 0.42 3.975 0.59 ;
      RECT  3.885 0.59 3.975 0.99 ;
      RECT  3.795 0.99 3.975 1.16 ;
      RECT  1.32 0.31 1.87 0.43 ;
      RECT  1.78 0.43 1.87 0.625 ;
      RECT  1.32 0.43 1.41 0.96 ;
      RECT  1.78 0.625 2.28 0.715 ;
      RECT  2.17 0.715 2.28 0.855 ;
      RECT  1.32 0.96 1.44 1.14 ;
      RECT  2.27 0.28 2.385 0.445 ;
      RECT  2.27 0.445 2.505 0.535 ;
      RECT  2.405 0.535 2.505 1.03 ;
      RECT  1.79 1.03 2.505 1.145 ;
      RECT  2.595 0.445 3.135 0.56 ;
      RECT  3.035 0.56 3.135 1.16 ;
      RECT  2.595 0.56 2.715 1.17 ;
      RECT  1.5 0.57 1.65 0.74 ;
      RECT  1.56 0.74 1.65 1.23 ;
      RECT  0.595 0.445 0.715 0.67 ;
      RECT  0.275 0.67 0.805 0.76 ;
      RECT  0.275 0.76 0.365 0.9 ;
      RECT  0.715 0.76 0.805 1.17 ;
      RECT  0.465 1.17 0.805 1.23 ;
      RECT  0.465 1.23 1.65 1.26 ;
      RECT  0.465 1.26 3.325 1.28 ;
      RECT  3.225 0.67 3.325 1.26 ;
      RECT  0.72 1.28 3.325 1.32 ;
      RECT  1.495 1.32 3.325 1.35 ;
      RECT  1.495 1.35 1.595 1.66 ;
      RECT  0.075 0.45 0.18 1.37 ;
      RECT  0.075 1.37 0.455 1.41 ;
      RECT  0.075 1.41 1.145 1.46 ;
      RECT  0.335 1.46 1.145 1.5 ;
      RECT  1.055 1.5 1.145 1.57 ;
      RECT  0.335 1.5 0.455 1.605 ;
      RECT  1.055 1.57 1.385 1.66 ;
  END
END SEN_FDPQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQ_2
#      Description : "D-Flip Flop, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQ_2
  CLASS CORE ;
  FOREIGN SEN_FDPQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.855 0.84 3.955 1.35 ;
      RECT  3.25 0.765 3.375 1.12 ;
      RECT  0.455 0.74 0.595 0.95 ;
      RECT  0.275 0.95 0.56 1.05 ;
      LAYER M2 ;
      RECT  0.38 0.95 4.0 1.05 ;
      LAYER V1 ;
      RECT  3.855 0.95 3.955 1.05 ;
      RECT  3.25 0.95 3.35 1.05 ;
      RECT  0.42 0.95 0.52 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0885 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.92 0.51 1.05 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0552 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.31 4.865 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.495 0.47 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.775 1.555 0.895 1.75 ;
      RECT  1.85 1.44 1.99 1.75 ;
      RECT  2.385 1.44 2.555 1.75 ;
      RECT  2.915 1.44 3.07 1.75 ;
      RECT  4.225 1.38 4.325 1.75 ;
      RECT  4.495 1.185 4.615 1.75 ;
      RECT  5.015 1.185 5.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.02 0.05 2.19 0.31 ;
      RECT  2.815 0.05 2.985 0.34 ;
      RECT  0.79 0.05 0.935 0.36 ;
      RECT  3.905 0.05 4.04 0.36 ;
      RECT  0.31 0.05 0.455 0.385 ;
      RECT  4.495 0.05 4.615 0.585 ;
      RECT  5.015 0.05 5.135 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.41 0.215 3.765 0.335 ;
      RECT  3.675 0.335 3.765 0.47 ;
      RECT  3.675 0.47 4.135 0.56 ;
      RECT  4.045 0.56 4.135 0.73 ;
      RECT  4.045 0.73 4.225 0.9 ;
      RECT  4.045 0.9 4.135 1.465 ;
      RECT  3.165 1.465 4.135 1.585 ;
      RECT  1.125 0.2 1.23 0.37 ;
      RECT  1.14 0.37 1.23 0.99 ;
      RECT  1.015 0.99 1.23 1.105 ;
      RECT  4.13 0.21 4.315 0.38 ;
      RECT  4.225 0.38 4.315 0.42 ;
      RECT  4.225 0.42 4.405 0.59 ;
      RECT  4.315 0.59 4.405 1.02 ;
      RECT  4.225 1.02 4.405 1.19 ;
      RECT  1.51 0.25 1.63 0.4 ;
      RECT  1.34 0.4 2.235 0.49 ;
      RECT  2.145 0.49 2.235 0.8 ;
      RECT  1.34 0.49 1.44 1.16 ;
      RECT  2.145 0.8 2.39 0.9 ;
      RECT  0.045 0.24 0.185 0.43 ;
      RECT  0.045 0.43 0.135 1.315 ;
      RECT  0.045 1.315 0.655 1.375 ;
      RECT  0.045 1.375 1.075 1.405 ;
      RECT  0.565 1.405 1.075 1.465 ;
      RECT  0.045 1.405 0.185 1.61 ;
      RECT  0.985 1.465 1.075 1.57 ;
      RECT  0.985 1.57 1.375 1.66 ;
      RECT  2.58 0.35 2.7 0.44 ;
      RECT  2.58 0.44 3.57 0.53 ;
      RECT  2.675 0.53 3.57 0.555 ;
      RECT  3.47 0.555 3.57 1.16 ;
      RECT  2.675 0.555 2.795 1.17 ;
      RECT  2.35 0.215 2.465 0.62 ;
      RECT  2.35 0.62 2.585 0.71 ;
      RECT  2.485 0.71 2.585 1.025 ;
      RECT  1.76 0.58 2.03 0.68 ;
      RECT  1.76 0.68 1.85 1.025 ;
      RECT  1.76 1.025 2.585 1.145 ;
      RECT  0.225 0.53 0.83 0.65 ;
      RECT  0.225 0.65 0.315 0.86 ;
      RECT  0.74 0.65 0.83 1.135 ;
      RECT  0.59 1.135 0.83 1.195 ;
      RECT  0.59 1.195 1.255 1.225 ;
      RECT  0.74 1.225 1.255 1.26 ;
      RECT  0.74 1.26 3.765 1.285 ;
      RECT  3.665 0.7 3.765 1.26 ;
      RECT  1.165 1.285 3.765 1.35 ;
      RECT  1.47 1.35 1.57 1.59 ;
  END
END SEN_FDPQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQ_4
#      Description : "D-Flip Flop, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQ_4
  CLASS CORE ;
  FOREIGN SEN_FDPQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.745 0.805 4.845 1.35 ;
      RECT  4.015 0.74 4.22 0.85 ;
      RECT  4.015 0.85 4.115 1.14 ;
      RECT  0.59 0.74 0.68 0.95 ;
      RECT  0.59 0.95 0.87 1.05 ;
      LAYER M2 ;
      RECT  0.62 0.95 4.95 1.05 ;
      LAYER V1 ;
      RECT  4.745 0.95 4.845 1.05 ;
      RECT  4.015 0.95 4.115 1.05 ;
      RECT  0.66 0.95 0.76 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1263 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  0.95 0.71 1.25 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0714 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.64 0.415 5.765 0.91 ;
      RECT  5.64 0.91 6.275 1.09 ;
      RECT  6.15 0.31 6.275 0.91 ;
      RECT  5.64 1.09 5.765 1.235 ;
      RECT  6.15 1.09 6.275 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.595 0.48 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.05 1.6 1.225 1.75 ;
      RECT  2.135 1.44 2.255 1.75 ;
      RECT  2.39 1.44 2.56 1.75 ;
      RECT  2.93 1.44 3.08 1.75 ;
      RECT  3.45 1.44 3.6 1.75 ;
      RECT  5.115 1.38 5.225 1.75 ;
      RECT  5.385 1.185 5.505 1.75 ;
      RECT  5.905 1.215 6.025 1.75 ;
      RECT  6.415 1.415 6.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.275 0.05 1.45 0.24 ;
      RECT  2.315 0.05 2.485 0.31 ;
      RECT  4.795 0.05 4.93 0.36 ;
      RECT  5.375 0.05 5.515 0.36 ;
      RECT  6.415 0.05 6.545 0.385 ;
      RECT  3.37 0.05 3.52 0.39 ;
      RECT  2.855 0.05 2.99 0.43 ;
      RECT  0.31 0.05 0.455 0.45 ;
      RECT  0.835 0.05 0.95 0.62 ;
      RECT  5.905 0.05 6.025 0.68 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.04 0.18 1.15 0.33 ;
      RECT  1.04 0.33 1.69 0.42 ;
      RECT  1.57 0.21 1.69 0.33 ;
      RECT  1.365 0.42 1.455 1.145 ;
      RECT  3.775 0.215 4.655 0.335 ;
      RECT  4.565 0.335 4.655 0.47 ;
      RECT  4.565 0.47 5.025 0.56 ;
      RECT  4.935 0.56 5.025 0.76 ;
      RECT  4.935 0.76 5.37 0.87 ;
      RECT  4.935 0.87 5.025 1.465 ;
      RECT  4.0 1.465 5.025 1.585 ;
      RECT  5.02 0.21 5.22 0.38 ;
      RECT  5.115 0.38 5.22 0.5 ;
      RECT  5.115 0.5 5.55 0.59 ;
      RECT  5.46 0.59 5.55 0.99 ;
      RECT  5.115 0.99 5.55 1.08 ;
      RECT  5.115 1.08 5.215 1.19 ;
      RECT  1.83 0.225 1.95 0.4 ;
      RECT  1.83 0.4 2.53 0.49 ;
      RECT  1.83 0.49 1.92 0.57 ;
      RECT  2.44 0.49 2.53 0.745 ;
      RECT  1.555 0.57 1.92 0.66 ;
      RECT  1.555 0.66 1.645 1.025 ;
      RECT  2.44 0.745 2.675 0.845 ;
      RECT  1.555 1.025 1.76 1.13 ;
      RECT  4.065 0.43 4.235 0.44 ;
      RECT  3.8 0.44 4.455 0.53 ;
      RECT  3.07 0.53 4.455 0.555 ;
      RECT  3.07 0.555 3.89 0.65 ;
      RECT  4.335 0.555 4.455 1.16 ;
      RECT  3.8 0.65 3.89 1.05 ;
      RECT  3.155 1.05 3.89 1.17 ;
      RECT  2.62 0.215 2.725 0.565 ;
      RECT  2.62 0.565 2.92 0.655 ;
      RECT  2.825 0.655 2.92 0.77 ;
      RECT  2.825 0.77 3.52 0.88 ;
      RECT  2.825 0.88 2.92 1.025 ;
      RECT  2.05 0.58 2.35 0.67 ;
      RECT  2.05 0.67 2.14 1.025 ;
      RECT  2.05 1.025 2.92 1.145 ;
      RECT  1.74 0.76 1.94 0.93 ;
      RECT  1.85 0.93 1.94 1.235 ;
      RECT  0.585 0.38 0.695 0.56 ;
      RECT  0.265 0.56 0.695 0.65 ;
      RECT  0.265 0.65 0.355 1.235 ;
      RECT  0.265 1.235 1.94 1.26 ;
      RECT  0.265 1.26 4.655 1.325 ;
      RECT  4.55 0.65 4.655 1.26 ;
      RECT  1.85 1.325 4.655 1.35 ;
      RECT  0.065 0.35 0.17 1.415 ;
      RECT  0.065 1.415 1.7 1.505 ;
      RECT  1.61 1.505 1.7 1.57 ;
      RECT  1.61 1.57 1.925 1.66 ;
  END
END SEN_FDPQ_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQ_D_1
#      Description : "D-Flip Flop, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FDPQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.5 1.05 0.94 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.34 0.31 3.46 1.29 ;
    END
    ANTENNADIFFAREA 0.2 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.8 1.44 0.93 1.75 ;
      RECT  1.785 1.575 1.91 1.75 ;
      RECT  2.79 1.54 2.92 1.75 ;
      RECT  3.6 1.21 3.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.795 0.05 0.925 0.39 ;
      RECT  1.8 0.05 1.925 0.39 ;
      RECT  2.79 0.05 2.92 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.6 0.05 3.72 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.25 0.185 1.71 0.3 ;
      RECT  1.62 0.3 1.71 0.74 ;
      RECT  1.39 0.74 1.98 0.83 ;
      RECT  1.88 0.63 1.98 0.74 ;
      RECT  1.39 0.83 1.48 1.31 ;
      RECT  1.24 1.31 1.48 1.43 ;
      RECT  2.27 0.22 2.55 0.34 ;
      RECT  2.46 0.34 2.55 0.88 ;
      RECT  2.46 0.88 2.975 0.97 ;
      RECT  2.875 0.97 2.975 1.33 ;
      RECT  2.27 1.33 2.975 1.45 ;
      RECT  1.42 0.39 1.53 0.55 ;
      RECT  1.2 0.55 1.53 0.65 ;
      RECT  1.2 0.65 1.3 1.08 ;
      RECT  0.49 0.24 0.69 0.36 ;
      RECT  0.6 0.36 0.69 1.0 ;
      RECT  0.54 1.0 0.69 1.08 ;
      RECT  0.54 1.08 1.3 1.17 ;
      RECT  3.065 0.26 3.185 0.59 ;
      RECT  2.655 0.59 3.185 0.705 ;
      RECT  3.065 0.705 3.185 0.755 ;
      RECT  3.065 0.755 3.25 0.925 ;
      RECT  3.065 0.925 3.185 1.46 ;
      RECT  2.26 0.51 2.36 1.105 ;
      RECT  2.26 1.105 2.625 1.215 ;
      RECT  1.65 0.92 1.765 1.185 ;
      RECT  1.65 1.185 2.17 1.29 ;
      RECT  2.07 0.24 2.17 1.185 ;
      RECT  1.57 1.385 2.095 1.475 ;
      RECT  1.57 1.475 1.66 1.54 ;
      RECT  2.0 1.475 2.095 1.56 ;
      RECT  0.34 0.47 0.46 0.74 ;
      RECT  0.34 0.74 0.51 0.91 ;
      RECT  0.34 0.91 0.43 1.26 ;
      RECT  0.34 1.26 1.14 1.35 ;
      RECT  1.05 1.35 1.14 1.54 ;
      RECT  0.34 1.35 0.46 1.61 ;
      RECT  1.05 1.54 1.66 1.65 ;
      RECT  2.0 1.56 2.39 1.66 ;
      LAYER M2 ;
      RECT  1.35 0.55 2.4 0.65 ;
      LAYER V1 ;
      RECT  1.39 0.55 1.49 0.65 ;
      RECT  2.26 0.55 2.36 0.65 ;
  END
END SEN_FDPQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQ_D_1P5
#      Description : "D-Flip Flop, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQ_D_1P5
  CLASS CORE ;
  FOREIGN SEN_FDPQ_D_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.925 0.51 1.25 0.69 ;
      RECT  0.925 0.69 1.05 0.97 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.31 3.85 1.385 ;
    END
    ANTENNADIFFAREA 0.172 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.44 0.195 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.775 1.455 0.905 1.75 ;
      RECT  1.815 1.615 1.985 1.75 ;
      RECT  2.96 1.215 3.08 1.75 ;
      RECT  3.475 1.215 3.595 1.75 ;
      RECT  4.01 1.215 4.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.065 0.05 0.195 0.385 ;
      RECT  0.805 0.05 0.945 0.41 ;
      RECT  2.95 0.05 3.09 0.415 ;
      RECT  1.865 0.05 1.98 0.42 ;
      RECT  3.475 0.05 3.595 0.56 ;
      RECT  4.01 0.05 4.13 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.3 0.24 1.775 0.36 ;
      RECT  1.685 0.36 1.775 0.715 ;
      RECT  1.555 0.715 2.035 0.805 ;
      RECT  1.945 0.805 2.035 0.915 ;
      RECT  1.555 0.805 1.645 0.99 ;
      RECT  1.36 0.99 1.645 1.08 ;
      RECT  1.36 1.08 1.48 1.16 ;
      RECT  2.125 0.24 2.345 0.36 ;
      RECT  2.125 0.36 2.215 1.07 ;
      RECT  1.735 0.99 1.825 1.07 ;
      RECT  1.735 1.07 2.215 1.16 ;
      RECT  3.22 0.31 3.34 0.58 ;
      RECT  2.75 0.58 3.34 0.67 ;
      RECT  3.23 0.67 3.34 0.78 ;
      RECT  3.23 0.78 3.655 0.89 ;
      RECT  3.23 0.89 3.34 1.4 ;
      RECT  1.375 0.48 1.595 0.59 ;
      RECT  1.375 0.59 1.465 0.81 ;
      RECT  1.175 0.81 1.465 0.9 ;
      RECT  1.175 0.9 1.265 1.08 ;
      RECT  0.555 0.19 0.69 0.36 ;
      RECT  0.6 0.36 0.69 1.0 ;
      RECT  0.52 1.0 0.69 1.08 ;
      RECT  0.52 1.08 1.265 1.17 ;
      RECT  1.175 1.17 1.265 1.25 ;
      RECT  1.175 1.25 2.7 1.34 ;
      RECT  2.305 0.56 2.395 1.25 ;
      RECT  2.61 1.34 2.7 1.66 ;
      RECT  0.34 0.21 0.43 0.73 ;
      RECT  0.34 0.73 0.505 0.9 ;
      RECT  0.34 0.9 0.43 1.26 ;
      RECT  0.34 1.26 1.085 1.35 ;
      RECT  0.995 1.35 1.085 1.43 ;
      RECT  0.34 1.35 0.445 1.61 ;
      RECT  0.995 1.43 2.41 1.52 ;
      RECT  2.3 1.52 2.41 1.64 ;
      RECT  1.48 1.52 1.59 1.66 ;
      RECT  2.485 0.19 2.59 0.785 ;
      RECT  2.485 0.785 3.135 0.875 ;
      RECT  3.03 0.875 3.135 0.995 ;
      RECT  2.485 0.875 2.59 1.16 ;
  END
END SEN_FDPQ_D_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQ_D_2
#      Description : "D-Flip Flop, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FDPQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.5 1.05 0.94 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.54 0.31 3.66 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.8 1.44 0.93 1.75 ;
      RECT  1.785 1.575 1.91 1.75 ;
      RECT  2.79 1.56 2.92 1.75 ;
      RECT  3.275 1.41 3.405 1.75 ;
      RECT  3.8 1.21 3.92 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.795 0.05 0.925 0.39 ;
      RECT  1.8 0.05 1.925 0.39 ;
      RECT  2.79 0.05 2.92 0.39 ;
      RECT  3.275 0.05 3.405 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.8 0.05 3.92 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.25 0.185 1.71 0.3 ;
      RECT  1.62 0.3 1.71 0.74 ;
      RECT  1.39 0.74 1.98 0.83 ;
      RECT  1.88 0.66 1.98 0.74 ;
      RECT  1.39 0.83 1.48 1.31 ;
      RECT  1.24 1.31 1.48 1.43 ;
      RECT  2.27 0.22 2.55 0.34 ;
      RECT  2.46 0.34 2.55 0.88 ;
      RECT  2.46 0.88 2.975 0.97 ;
      RECT  2.875 0.97 2.975 1.33 ;
      RECT  2.27 1.33 2.975 1.45 ;
      RECT  1.42 0.39 1.53 0.55 ;
      RECT  1.2 0.55 1.53 0.65 ;
      RECT  1.2 0.65 1.3 1.08 ;
      RECT  0.49 0.24 0.69 0.36 ;
      RECT  0.6 0.36 0.69 1.0 ;
      RECT  0.54 1.0 0.69 1.08 ;
      RECT  0.54 1.08 1.3 1.17 ;
      RECT  3.065 0.39 3.185 0.635 ;
      RECT  2.655 0.635 3.185 0.75 ;
      RECT  3.065 0.75 3.185 0.785 ;
      RECT  3.065 0.785 3.45 0.895 ;
      RECT  3.065 0.895 3.185 1.33 ;
      RECT  2.26 0.485 2.36 1.105 ;
      RECT  2.26 1.105 2.625 1.215 ;
      RECT  1.65 0.92 1.765 1.185 ;
      RECT  1.65 1.185 2.17 1.29 ;
      RECT  2.07 0.24 2.17 1.185 ;
      RECT  1.57 1.385 2.095 1.475 ;
      RECT  1.57 1.475 1.66 1.54 ;
      RECT  2.0 1.475 2.095 1.56 ;
      RECT  0.34 0.47 0.46 0.74 ;
      RECT  0.34 0.74 0.51 0.91 ;
      RECT  0.34 0.91 0.43 1.26 ;
      RECT  0.34 1.26 1.14 1.35 ;
      RECT  1.05 1.35 1.14 1.54 ;
      RECT  0.34 1.35 0.46 1.61 ;
      RECT  1.05 1.54 1.66 1.65 ;
      RECT  2.0 1.56 2.39 1.66 ;
      LAYER M2 ;
      RECT  1.35 0.55 2.4 0.65 ;
      LAYER V1 ;
      RECT  1.39 0.55 1.49 0.65 ;
      RECT  2.26 0.55 2.36 0.65 ;
  END
END SEN_FDPQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQ_D_3
#      Description : "D-Flip Flop, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQ_D_3
  CLASS CORE ;
  FOREIGN SEN_FDPQ_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.25 0.69 ;
      RECT  0.95 0.69 1.05 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.31 4.45 0.47 ;
      RECT  3.77 0.47 4.45 0.59 ;
      RECT  4.35 0.59 4.45 1.11 ;
      RECT  3.8 1.11 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.415 0.195 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.825 1.44 0.945 1.75 ;
      RECT  1.89 1.615 2.06 1.75 ;
      RECT  3.035 1.19 3.155 1.75 ;
      RECT  3.56 1.215 3.68 1.75 ;
      RECT  4.07 1.415 4.21 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  4.07 0.05 4.21 0.37 ;
      RECT  0.065 0.05 0.195 0.385 ;
      RECT  3.03 0.05 3.17 0.41 ;
      RECT  0.825 0.05 0.965 0.415 ;
      RECT  1.925 0.05 2.055 0.42 ;
      RECT  3.56 0.05 3.68 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.36 0.24 1.835 0.36 ;
      RECT  1.745 0.36 1.835 0.71 ;
      RECT  1.62 0.71 2.095 0.8 ;
      RECT  1.985 0.58 2.095 0.71 ;
      RECT  1.62 0.8 1.71 0.99 ;
      RECT  1.43 0.99 1.71 1.08 ;
      RECT  1.43 1.08 1.55 1.16 ;
      RECT  3.325 0.39 3.415 0.545 ;
      RECT  2.86 0.545 3.415 0.655 ;
      RECT  3.325 0.655 3.415 0.785 ;
      RECT  3.325 0.785 4.24 0.895 ;
      RECT  3.325 0.895 3.43 1.29 ;
      RECT  1.44 0.455 1.65 0.565 ;
      RECT  1.44 0.565 1.53 0.81 ;
      RECT  1.215 0.81 1.53 0.9 ;
      RECT  1.215 0.9 1.315 1.08 ;
      RECT  0.575 0.215 0.695 0.435 ;
      RECT  0.595 0.435 0.695 1.0 ;
      RECT  0.59 1.0 0.695 1.08 ;
      RECT  0.59 1.08 1.315 1.17 ;
      RECT  1.215 1.17 1.315 1.25 ;
      RECT  1.215 1.25 2.79 1.34 ;
      RECT  2.39 0.53 2.48 1.25 ;
      RECT  2.675 1.34 2.79 1.66 ;
      RECT  0.34 0.445 0.445 0.77 ;
      RECT  0.34 0.77 0.505 0.94 ;
      RECT  0.34 0.94 0.43 1.26 ;
      RECT  0.34 1.26 1.125 1.35 ;
      RECT  1.035 1.35 1.125 1.435 ;
      RECT  0.34 1.35 0.445 1.575 ;
      RECT  1.035 1.435 2.515 1.525 ;
      RECT  1.55 1.525 1.66 1.66 ;
      RECT  2.405 1.525 2.515 1.66 ;
      RECT  2.57 0.19 2.675 0.88 ;
      RECT  2.57 0.88 3.215 0.97 ;
      RECT  3.105 0.765 3.215 0.88 ;
      RECT  2.57 0.97 2.675 1.16 ;
      RECT  1.8 0.915 1.91 1.055 ;
      RECT  1.8 1.055 2.3 1.145 ;
      RECT  2.195 0.255 2.3 1.055 ;
  END
END SEN_FDPQ_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQ_D_4
#      Description : "D-Flip Flop, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FDPQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.5 1.05 0.94 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 4.26 0.69 ;
      RECT  4.15 0.69 4.26 1.105 ;
      RECT  3.55 1.105 4.26 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.8 1.44 0.93 1.75 ;
      RECT  1.785 1.575 1.91 1.75 ;
      RECT  2.8 1.56 2.93 1.75 ;
      RECT  3.34 1.21 3.46 1.75 ;
      RECT  3.875 1.415 4.005 1.75 ;
      RECT  4.4 1.21 4.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.795 0.05 0.925 0.39 ;
      RECT  1.8 0.05 1.925 0.39 ;
      RECT  2.805 0.05 2.935 0.39 ;
      RECT  3.875 0.05 4.005 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.34 0.05 3.46 0.59 ;
      RECT  4.4 0.05 4.52 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.25 0.185 1.71 0.3 ;
      RECT  1.62 0.3 1.71 0.74 ;
      RECT  1.39 0.74 1.98 0.83 ;
      RECT  1.88 0.63 1.98 0.74 ;
      RECT  1.39 0.83 1.48 1.31 ;
      RECT  1.24 1.31 1.48 1.43 ;
      RECT  2.27 0.22 2.55 0.34 ;
      RECT  2.46 0.34 2.55 0.785 ;
      RECT  2.46 0.785 3.0 0.875 ;
      RECT  2.9 0.875 3.0 1.33 ;
      RECT  2.27 1.33 3.0 1.45 ;
      RECT  1.42 0.39 1.53 0.55 ;
      RECT  1.2 0.55 1.53 0.65 ;
      RECT  1.2 0.65 1.3 1.08 ;
      RECT  0.49 0.24 0.69 0.36 ;
      RECT  0.6 0.36 0.69 1.0 ;
      RECT  0.54 1.0 0.69 1.08 ;
      RECT  0.54 1.08 1.3 1.17 ;
      RECT  3.09 0.42 3.21 0.55 ;
      RECT  2.64 0.55 3.21 0.665 ;
      RECT  3.09 0.665 3.21 0.785 ;
      RECT  3.09 0.785 4.06 0.895 ;
      RECT  3.09 0.895 3.21 1.24 ;
      RECT  2.26 0.485 2.36 1.105 ;
      RECT  2.26 1.105 2.625 1.215 ;
      RECT  1.65 0.92 1.765 1.185 ;
      RECT  1.65 1.185 2.17 1.29 ;
      RECT  2.07 0.24 2.17 1.185 ;
      RECT  1.57 1.385 2.095 1.475 ;
      RECT  1.57 1.475 1.66 1.54 ;
      RECT  2.0 1.475 2.095 1.56 ;
      RECT  0.34 0.47 0.46 0.74 ;
      RECT  0.34 0.74 0.51 0.91 ;
      RECT  0.34 0.91 0.43 1.26 ;
      RECT  0.34 1.26 1.14 1.35 ;
      RECT  1.05 1.35 1.14 1.54 ;
      RECT  0.34 1.35 0.46 1.61 ;
      RECT  1.05 1.54 1.66 1.65 ;
      RECT  2.0 1.56 2.39 1.66 ;
      LAYER M2 ;
      RECT  1.35 0.55 2.4 0.65 ;
      LAYER V1 ;
      RECT  1.39 0.55 1.49 0.65 ;
      RECT  2.26 0.55 2.36 0.65 ;
  END
END SEN_FDPQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQB_1
#      Description : "D-Flip Flop, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQB_1
  CLASS CORE ;
  FOREIGN SEN_FDPQB_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0453 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.31 4.335 0.485 ;
      RECT  4.15 0.485 4.25 1.0 ;
      RECT  4.15 1.0 4.335 1.09 ;
      RECT  4.215 1.09 4.335 1.24 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.095 1.415 0.225 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.855 1.63 1.025 1.75 ;
      RECT  2.23 1.63 2.4 1.75 ;
      RECT  3.655 1.44 3.795 1.75 ;
      RECT  3.955 1.215 4.075 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.985 0.05 1.125 0.225 ;
      RECT  0.095 0.05 0.235 0.365 ;
      RECT  3.405 0.05 3.545 0.38 ;
      RECT  2.36 0.05 2.5 0.42 ;
      RECT  3.93 0.05 4.06 0.425 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.515 0.21 1.635 0.34 ;
      RECT  0.925 0.34 1.635 0.46 ;
      RECT  0.925 0.46 1.015 1.025 ;
      RECT  0.925 1.025 1.365 1.12 ;
      RECT  1.75 0.235 2.255 0.355 ;
      RECT  2.165 0.355 2.255 0.725 ;
      RECT  1.75 0.355 1.87 1.16 ;
      RECT  2.165 0.725 2.485 0.815 ;
      RECT  2.395 0.815 2.485 0.95 ;
      RECT  2.845 0.235 3.255 0.355 ;
      RECT  3.165 0.355 3.255 0.725 ;
      RECT  3.165 0.725 3.665 0.825 ;
      RECT  3.46 0.825 3.665 0.895 ;
      RECT  3.46 0.895 3.55 1.465 ;
      RECT  3.06 1.465 3.55 1.585 ;
      RECT  2.62 0.21 2.755 0.38 ;
      RECT  2.62 0.38 2.71 1.06 ;
      RECT  2.165 0.92 2.265 1.06 ;
      RECT  2.165 1.06 2.71 1.18 ;
      RECT  3.68 0.18 3.785 0.475 ;
      RECT  3.345 0.475 3.785 0.48 ;
      RECT  3.345 0.48 3.845 0.58 ;
      RECT  3.755 0.58 3.845 0.99 ;
      RECT  3.7 0.99 3.845 1.16 ;
      RECT  0.34 0.3 0.48 0.63 ;
      RECT  0.34 0.63 0.645 0.8 ;
      RECT  0.34 0.8 0.43 1.45 ;
      RECT  0.34 1.45 1.425 1.52 ;
      RECT  0.34 1.52 2.83 1.54 ;
      RECT  1.99 1.45 2.83 1.52 ;
      RECT  1.335 1.54 2.095 1.63 ;
      RECT  2.72 1.54 2.83 1.66 ;
      RECT  2.8 0.585 2.89 1.265 ;
      RECT  2.8 1.265 3.37 1.27 ;
      RECT  3.28 1.16 3.37 1.265 ;
      RECT  0.735 0.185 0.835 1.24 ;
      RECT  0.545 1.24 0.835 1.25 ;
      RECT  0.545 1.25 2.075 1.27 ;
      RECT  1.985 0.47 2.075 1.25 ;
      RECT  0.545 1.27 3.37 1.36 ;
  END
END SEN_FDPQB_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQB_2
#      Description : "D-Flip Flop, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQB_2
  CLASS CORE ;
  FOREIGN SEN_FDPQB_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0414 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.71 ;
      RECT  1.55 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.715 0.31 5.85 0.545 ;
      RECT  5.75 0.545 5.85 1.25 ;
      RECT  5.715 1.25 5.85 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.61 0.48 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.85 1.61 1.02 1.75 ;
      RECT  1.41 1.61 1.58 1.75 ;
      RECT  2.925 1.575 3.065 1.75 ;
      RECT  3.425 1.575 3.565 1.75 ;
      RECT  5.165 1.44 5.3 1.75 ;
      RECT  5.45 1.44 5.58 1.75 ;
      RECT  5.995 1.215 6.115 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  1.105 0.05 1.275 0.225 ;
      RECT  3.55 0.05 3.69 0.36 ;
      RECT  3.015 0.05 3.145 0.39 ;
      RECT  0.16 0.05 0.3 0.4 ;
      RECT  4.92 0.05 5.06 0.405 ;
      RECT  1.66 0.05 1.78 0.46 ;
      RECT  5.455 0.05 5.575 0.585 ;
      RECT  5.995 0.05 6.115 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.875 0.215 2.925 0.335 ;
      RECT  2.835 0.335 2.925 0.785 ;
      RECT  2.455 0.335 2.555 1.09 ;
      RECT  2.835 0.785 3.515 0.895 ;
      RECT  3.87 0.215 4.75 0.335 ;
      RECT  4.66 0.335 4.75 0.995 ;
      RECT  4.66 0.995 5.05 1.085 ;
      RECT  4.96 1.085 5.05 1.25 ;
      RECT  4.96 1.25 5.59 1.34 ;
      RECT  5.49 0.715 5.59 1.25 ;
      RECT  4.96 1.34 5.05 1.465 ;
      RECT  3.92 1.39 4.67 1.465 ;
      RECT  3.92 1.465 5.05 1.48 ;
      RECT  4.56 1.48 5.05 1.585 ;
      RECT  1.155 0.34 1.57 0.46 ;
      RECT  1.155 0.46 1.26 0.98 ;
      RECT  1.155 0.98 2.31 1.07 ;
      RECT  2.19 0.43 2.31 0.98 ;
      RECT  1.155 1.07 1.275 1.16 ;
      RECT  3.215 0.475 4.36 0.595 ;
      RECT  3.215 0.595 3.85 0.6 ;
      RECT  3.76 0.6 3.85 1.0 ;
      RECT  2.835 1.0 4.39 1.12 ;
      RECT  5.185 0.165 5.305 0.78 ;
      RECT  4.86 0.78 5.305 0.89 ;
      RECT  5.185 0.89 5.305 1.16 ;
      RECT  4.15 0.74 4.57 0.85 ;
      RECT  4.48 0.85 4.57 1.18 ;
      RECT  4.48 1.18 4.87 1.21 ;
      RECT  1.66 1.17 1.75 1.18 ;
      RECT  1.545 1.18 2.745 1.21 ;
      RECT  2.655 0.45 2.745 1.18 ;
      RECT  1.545 1.21 4.87 1.25 ;
      RECT  0.655 0.25 0.85 0.37 ;
      RECT  0.75 0.37 0.85 1.17 ;
      RECT  0.62 1.17 0.85 1.25 ;
      RECT  0.62 1.25 4.87 1.27 ;
      RECT  2.655 1.27 4.87 1.3 ;
      RECT  0.62 1.27 1.76 1.34 ;
      RECT  4.78 1.3 4.87 1.35 ;
      RECT  1.85 1.36 2.56 1.46 ;
      RECT  2.71 1.395 3.83 1.485 ;
      RECT  2.71 1.485 2.8 1.57 ;
      RECT  3.74 1.485 3.83 1.57 ;
      RECT  0.44 0.46 0.575 0.91 ;
      RECT  0.44 0.91 0.635 1.08 ;
      RECT  0.44 1.08 0.53 1.43 ;
      RECT  0.065 1.305 0.185 1.43 ;
      RECT  0.065 1.43 1.76 1.52 ;
      RECT  1.67 1.52 1.76 1.57 ;
      RECT  1.67 1.57 2.8 1.66 ;
      RECT  3.74 1.57 4.32 1.66 ;
  END
END SEN_FDPQB_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQB_3
#      Description : "D-Flip Flop, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQB_3
  CLASS CORE ;
  FOREIGN SEN_FDPQB_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.71 ;
      RECT  1.55 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0786 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.615 0.315 6.735 0.45 ;
      RECT  6.045 0.45 6.735 0.54 ;
      RECT  6.045 0.54 6.45 0.57 ;
      RECT  6.35 0.57 6.45 1.11 ;
      RECT  6.095 1.11 6.72 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.46 1.595 0.63 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.0 1.595 1.17 1.75 ;
      RECT  1.575 1.575 1.705 1.75 ;
      RECT  3.04 1.575 3.21 1.75 ;
      RECT  3.3 1.575 3.47 1.75 ;
      RECT  3.84 1.575 4.01 1.75 ;
      RECT  5.515 1.43 5.655 1.75 ;
      RECT  5.825 1.43 5.965 1.75 ;
      RECT  6.345 1.415 6.485 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  1.18 0.05 1.32 0.235 ;
      RECT  6.345 0.05 6.485 0.345 ;
      RECT  3.665 0.05 3.805 0.36 ;
      RECT  3.145 0.05 3.285 0.39 ;
      RECT  5.275 0.05 5.415 0.39 ;
      RECT  0.07 0.05 0.205 0.395 ;
      RECT  1.78 0.05 1.91 0.4 ;
      RECT  0.595 0.05 0.735 0.44 ;
      RECT  5.835 0.05 5.955 0.595 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.01 0.215 3.04 0.335 ;
      RECT  2.95 0.335 3.04 0.785 ;
      RECT  2.59 0.335 2.68 1.07 ;
      RECT  2.95 0.785 4.085 0.895 ;
      RECT  3.365 0.475 4.625 0.595 ;
      RECT  4.19 0.595 4.625 0.61 ;
      RECT  4.19 0.61 4.28 1.005 ;
      RECT  2.95 1.005 4.28 1.015 ;
      RECT  2.95 1.015 4.835 1.12 ;
      RECT  2.345 0.43 2.5 0.6 ;
      RECT  2.41 0.6 2.5 0.98 ;
      RECT  1.28 0.34 1.68 0.46 ;
      RECT  1.28 0.46 1.37 0.98 ;
      RECT  1.28 0.98 2.5 1.09 ;
      RECT  1.28 1.09 1.45 1.125 ;
      RECT  5.565 0.17 5.71 0.735 ;
      RECT  5.29 0.735 5.71 0.845 ;
      RECT  5.61 0.845 5.71 1.015 ;
      RECT  5.52 1.015 5.71 1.135 ;
      RECT  4.555 0.7 4.645 0.83 ;
      RECT  4.555 0.83 5.015 0.925 ;
      RECT  4.925 0.925 5.015 1.18 ;
      RECT  4.925 1.18 5.23 1.21 ;
      RECT  2.77 0.45 2.86 1.18 ;
      RECT  1.575 1.18 2.86 1.21 ;
      RECT  1.575 1.21 5.23 1.215 ;
      RECT  0.855 0.3 0.965 0.525 ;
      RECT  0.875 0.525 0.965 1.17 ;
      RECT  0.73 1.17 0.965 1.215 ;
      RECT  0.73 1.215 5.23 1.27 ;
      RECT  2.775 1.27 5.23 1.3 ;
      RECT  0.73 1.27 1.665 1.305 ;
      RECT  5.14 1.3 5.23 1.35 ;
      RECT  5.835 0.785 6.26 0.895 ;
      RECT  5.835 0.895 5.93 1.225 ;
      RECT  4.135 0.215 5.0 0.335 ;
      RECT  4.91 0.335 5.0 0.65 ;
      RECT  4.91 0.65 5.195 0.74 ;
      RECT  5.105 0.74 5.195 0.96 ;
      RECT  5.105 0.96 5.41 1.07 ;
      RECT  5.32 1.07 5.41 1.225 ;
      RECT  5.32 1.225 5.93 1.315 ;
      RECT  5.32 1.315 5.41 1.465 ;
      RECT  4.37 1.39 5.055 1.465 ;
      RECT  4.37 1.465 5.41 1.48 ;
      RECT  4.945 1.48 5.41 1.585 ;
      RECT  1.975 1.365 2.71 1.475 ;
      RECT  2.8 1.395 4.28 1.485 ;
      RECT  2.8 1.485 2.89 1.57 ;
      RECT  4.19 1.485 4.28 1.57 ;
      RECT  0.34 0.22 0.465 0.83 ;
      RECT  0.34 0.83 0.785 1.0 ;
      RECT  0.34 1.0 0.43 1.395 ;
      RECT  0.215 1.395 1.885 1.485 ;
      RECT  1.795 1.485 1.885 1.57 ;
      RECT  0.215 1.485 0.335 1.615 ;
      RECT  1.795 1.57 2.89 1.66 ;
      RECT  4.19 1.57 4.765 1.66 ;
  END
END SEN_FDPQB_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQB_4
#      Description : "D-Flip Flop, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQB_4
  CLASS CORE ;
  FOREIGN SEN_FDPQB_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0585 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.71 ;
      RECT  1.55 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0906 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.92 0.31 7.05 0.445 ;
      RECT  6.35 0.445 7.05 0.56 ;
      RECT  6.95 0.56 7.05 1.11 ;
      RECT  6.35 1.11 7.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.48 1.6 0.65 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  1.02 1.6 1.19 1.75 ;
      RECT  1.595 1.575 1.725 1.75 ;
      RECT  3.06 1.6 3.23 1.75 ;
      RECT  3.58 1.6 3.75 1.75 ;
      RECT  4.12 1.6 4.29 1.75 ;
      RECT  5.805 1.405 5.945 1.75 ;
      RECT  6.13 1.405 6.27 1.75 ;
      RECT  6.65 1.415 6.79 1.75 ;
      RECT  7.2 1.21 7.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  1.205 0.05 1.375 0.24 ;
      RECT  6.65 0.05 6.79 0.345 ;
      RECT  3.745 0.05 3.885 0.385 ;
      RECT  4.265 0.05 4.395 0.385 ;
      RECT  0.085 0.05 0.225 0.39 ;
      RECT  1.825 0.05 1.995 0.395 ;
      RECT  3.225 0.05 3.365 0.395 ;
      RECT  5.56 0.05 5.7 0.4 ;
      RECT  0.615 0.05 0.745 0.45 ;
      RECT  6.14 0.05 6.26 0.59 ;
      RECT  7.2 0.05 7.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.085 0.215 3.12 0.32 ;
      RECT  2.62 0.32 3.12 0.335 ;
      RECT  3.03 0.335 3.12 0.785 ;
      RECT  2.62 0.335 2.71 1.05 ;
      RECT  3.03 0.785 4.07 0.89 ;
      RECT  4.775 0.41 4.97 0.48 ;
      RECT  3.44 0.48 4.97 0.58 ;
      RECT  3.44 0.58 4.56 0.6 ;
      RECT  4.47 0.6 4.56 0.98 ;
      RECT  3.06 0.98 4.56 1.03 ;
      RECT  3.06 1.03 5.075 1.12 ;
      RECT  4.97 0.93 5.075 1.03 ;
      RECT  3.06 1.12 3.48 1.15 ;
      RECT  2.32 0.415 2.53 0.535 ;
      RECT  2.44 0.535 2.53 0.98 ;
      RECT  1.3 0.33 1.705 0.5 ;
      RECT  1.3 0.5 1.39 0.98 ;
      RECT  1.3 0.98 2.53 1.07 ;
      RECT  1.3 1.07 1.47 1.12 ;
      RECT  5.87 0.18 6.015 0.79 ;
      RECT  5.54 0.79 6.015 0.89 ;
      RECT  5.925 0.89 6.015 1.015 ;
      RECT  5.815 1.015 6.015 1.135 ;
      RECT  4.755 0.71 5.255 0.82 ;
      RECT  5.165 0.82 5.255 1.18 ;
      RECT  5.165 1.18 5.51 1.21 ;
      RECT  4.47 1.21 5.51 1.24 ;
      RECT  2.85 0.45 2.94 1.16 ;
      RECT  1.84 1.16 2.94 1.215 ;
      RECT  0.835 0.34 1.03 0.46 ;
      RECT  0.935 0.46 1.03 1.185 ;
      RECT  0.72 1.185 1.03 1.215 ;
      RECT  0.72 1.215 2.94 1.24 ;
      RECT  0.72 1.24 5.51 1.25 ;
      RECT  2.85 1.25 5.51 1.3 ;
      RECT  0.72 1.25 1.925 1.305 ;
      RECT  2.85 1.3 4.56 1.33 ;
      RECT  5.42 1.3 5.51 1.35 ;
      RECT  6.12 0.785 6.84 0.895 ;
      RECT  6.12 0.895 6.21 1.225 ;
      RECT  4.49 0.2 5.435 0.32 ;
      RECT  5.345 0.32 5.435 0.98 ;
      RECT  5.345 0.98 5.69 1.09 ;
      RECT  5.6 1.09 5.69 1.225 ;
      RECT  5.6 1.225 6.21 1.315 ;
      RECT  5.6 1.315 5.69 1.465 ;
      RECT  4.65 1.39 5.31 1.465 ;
      RECT  4.65 1.465 5.69 1.48 ;
      RECT  5.2 1.48 5.69 1.585 ;
      RECT  2.01 1.34 2.76 1.455 ;
      RECT  2.88 1.42 4.56 1.51 ;
      RECT  2.88 1.51 2.97 1.57 ;
      RECT  4.47 1.51 4.56 1.57 ;
      RECT  0.365 0.285 0.485 0.88 ;
      RECT  0.365 0.88 0.845 0.99 ;
      RECT  0.365 0.99 0.475 1.355 ;
      RECT  0.235 1.355 0.475 1.395 ;
      RECT  0.235 1.395 1.905 1.485 ;
      RECT  1.815 1.485 1.905 1.57 ;
      RECT  0.235 1.485 0.36 1.58 ;
      RECT  1.815 1.57 2.97 1.66 ;
      RECT  4.47 1.57 5.045 1.66 ;
  END
END SEN_FDPQB_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQB_D_1
#      Description : "D-Flip Flop, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQB_D_1
  CLASS CORE ;
  FOREIGN SEN_FDPQB_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0375 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.48 1.05 0.995 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.51 3.945 0.68 ;
      RECT  3.75 0.68 3.85 0.99 ;
      RECT  3.75 0.99 3.945 1.09 ;
      RECT  3.825 1.09 3.945 1.2 ;
    END
    ANTENNADIFFAREA 0.142 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.815 1.48 0.985 1.75 ;
      RECT  1.955 1.575 2.095 1.75 ;
      RECT  3.055 1.05 3.18 1.75 ;
      RECT  3.565 1.225 3.685 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  0.85 0.05 0.97 0.39 ;
      RECT  3.55 0.05 3.69 0.39 ;
      RECT  2.99 0.05 3.13 0.395 ;
      RECT  1.895 0.05 2.035 0.405 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.315 0.215 1.79 0.335 ;
      RECT  1.7 0.335 1.79 0.75 ;
      RECT  1.47 0.75 2.095 0.84 ;
      RECT  1.995 0.645 2.095 0.75 ;
      RECT  1.47 0.84 1.575 1.125 ;
      RECT  2.39 0.235 2.7 0.355 ;
      RECT  2.61 0.355 2.7 0.785 ;
      RECT  2.61 0.785 3.44 0.895 ;
      RECT  2.61 0.895 2.715 1.24 ;
      RECT  3.28 0.185 3.4 0.58 ;
      RECT  2.82 0.58 3.4 0.59 ;
      RECT  2.82 0.59 3.65 0.69 ;
      RECT  3.55 0.69 3.65 1.015 ;
      RECT  3.27 1.015 3.65 1.135 ;
      RECT  0.34 0.38 0.47 0.685 ;
      RECT  0.34 0.685 0.58 0.86 ;
      RECT  0.34 0.86 0.43 1.3 ;
      RECT  0.34 1.3 1.2 1.39 ;
      RECT  1.11 1.39 1.2 1.395 ;
      RECT  0.34 1.39 0.445 1.61 ;
      RECT  1.11 1.395 2.34 1.485 ;
      RECT  2.25 1.485 2.34 1.545 ;
      RECT  2.25 1.545 2.6 1.645 ;
      RECT  2.365 0.625 2.52 0.795 ;
      RECT  2.43 0.795 2.52 1.215 ;
      RECT  1.22 0.45 1.61 0.62 ;
      RECT  1.22 0.62 1.31 1.085 ;
      RECT  1.22 1.085 1.38 1.105 ;
      RECT  0.585 0.19 0.76 0.36 ;
      RECT  0.67 0.36 0.76 1.105 ;
      RECT  0.53 1.105 1.38 1.21 ;
      RECT  1.29 1.21 1.38 1.215 ;
      RECT  1.29 1.215 2.52 1.305 ;
      RECT  2.43 1.305 2.52 1.33 ;
      RECT  2.43 1.33 2.815 1.42 ;
      RECT  2.725 1.42 2.815 1.65 ;
      RECT  2.185 0.32 2.275 0.93 ;
      RECT  1.805 0.93 2.275 0.955 ;
      RECT  1.805 0.955 2.34 1.125 ;
  END
END SEN_FDPQB_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQB_D_2
#      Description : "D-Flip Flop, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQB_D_2
  CLASS CORE ;
  FOREIGN SEN_FDPQB_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0375 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.48 1.05 0.995 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.31 3.87 0.535 ;
      RECT  3.75 0.535 3.85 1.26 ;
      RECT  3.75 1.26 3.87 1.49 ;
    END
    ANTENNADIFFAREA 0.218 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.825 1.48 0.995 1.75 ;
      RECT  1.965 1.575 2.105 1.75 ;
      RECT  3.075 1.24 3.2 1.75 ;
      RECT  3.495 1.225 3.615 1.75 ;
      RECT  4.015 1.215 4.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  2.91 0.05 3.05 0.375 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  0.85 0.05 0.98 0.39 ;
      RECT  1.91 0.05 2.04 0.405 ;
      RECT  3.48 0.05 3.62 0.41 ;
      RECT  4.015 0.05 4.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.335 0.215 1.8 0.335 ;
      RECT  1.71 0.335 1.8 0.75 ;
      RECT  1.48 0.75 2.105 0.84 ;
      RECT  2.005 0.645 2.105 0.75 ;
      RECT  1.48 0.84 1.57 1.125 ;
      RECT  2.39 0.235 2.71 0.355 ;
      RECT  2.62 0.355 2.71 0.745 ;
      RECT  2.62 0.745 3.46 0.855 ;
      RECT  2.62 0.855 2.725 1.24 ;
      RECT  2.84 0.485 2.95 0.565 ;
      RECT  2.84 0.565 3.66 0.655 ;
      RECT  3.21 0.185 3.33 0.565 ;
      RECT  3.57 0.655 3.66 1.015 ;
      RECT  3.175 1.015 3.66 1.135 ;
      RECT  0.34 0.385 0.46 0.755 ;
      RECT  0.34 0.755 0.58 0.925 ;
      RECT  0.34 0.925 0.43 1.3 ;
      RECT  0.34 1.3 1.21 1.39 ;
      RECT  1.12 1.39 1.21 1.395 ;
      RECT  0.34 1.39 0.445 1.61 ;
      RECT  1.12 1.395 2.35 1.485 ;
      RECT  2.26 1.485 2.35 1.545 ;
      RECT  2.26 1.545 2.61 1.645 ;
      RECT  2.375 0.625 2.53 0.795 ;
      RECT  2.44 0.795 2.53 1.215 ;
      RECT  1.23 0.45 1.62 0.62 ;
      RECT  1.23 0.62 1.32 1.085 ;
      RECT  1.23 1.085 1.39 1.105 ;
      RECT  0.59 0.19 0.76 0.36 ;
      RECT  0.67 0.36 0.76 1.105 ;
      RECT  0.54 1.105 1.39 1.21 ;
      RECT  1.3 1.21 1.39 1.215 ;
      RECT  1.3 1.215 2.53 1.305 ;
      RECT  2.44 1.305 2.53 1.33 ;
      RECT  2.44 1.33 2.825 1.42 ;
      RECT  2.73 1.42 2.825 1.65 ;
      RECT  2.195 0.32 2.285 0.955 ;
      RECT  2.195 0.955 2.35 0.96 ;
      RECT  1.77 0.96 2.35 1.125 ;
  END
END SEN_FDPQB_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQB_D_3
#      Description : "D-Flip Flop, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQB_D_3
  CLASS CORE ;
  FOREIGN SEN_FDPQB_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0375 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.48 1.05 0.98 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.21 0.42 4.335 0.475 ;
      RECT  3.64 0.475 4.335 0.59 ;
      RECT  3.95 0.59 4.05 1.11 ;
      RECT  3.695 1.11 4.335 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.825 1.48 0.995 1.75 ;
      RECT  1.965 1.575 2.105 1.75 ;
      RECT  3.075 1.43 3.215 1.75 ;
      RECT  3.425 1.425 3.565 1.75 ;
      RECT  3.945 1.41 4.085 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  3.94 0.05 4.08 0.385 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  0.85 0.05 0.98 0.39 ;
      RECT  3.42 0.05 3.56 0.39 ;
      RECT  2.89 0.05 3.03 0.405 ;
      RECT  1.905 0.05 2.045 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.335 0.215 1.8 0.335 ;
      RECT  1.71 0.335 1.8 0.75 ;
      RECT  1.48 0.75 2.105 0.84 ;
      RECT  2.015 0.64 2.105 0.75 ;
      RECT  1.48 0.84 1.585 1.125 ;
      RECT  3.165 0.18 3.285 0.745 ;
      RECT  2.82 0.745 3.285 0.755 ;
      RECT  2.82 0.755 3.31 0.855 ;
      RECT  3.22 0.855 3.31 1.015 ;
      RECT  3.125 1.015 3.31 1.135 ;
      RECT  0.34 0.39 0.48 0.755 ;
      RECT  0.34 0.755 0.58 0.925 ;
      RECT  0.34 0.925 0.43 1.3 ;
      RECT  0.34 1.3 1.21 1.39 ;
      RECT  1.12 1.39 1.21 1.395 ;
      RECT  0.34 1.39 0.445 1.61 ;
      RECT  1.12 1.395 2.35 1.485 ;
      RECT  2.26 1.485 2.35 1.545 ;
      RECT  2.26 1.545 2.61 1.645 ;
      RECT  2.375 0.625 2.53 0.795 ;
      RECT  2.44 0.795 2.53 1.215 ;
      RECT  1.23 0.45 1.62 0.62 ;
      RECT  1.23 0.62 1.32 1.105 ;
      RECT  0.605 0.19 0.76 0.36 ;
      RECT  0.67 0.36 0.76 1.105 ;
      RECT  0.54 1.105 1.39 1.21 ;
      RECT  1.3 1.21 1.39 1.215 ;
      RECT  1.3 1.215 2.53 1.305 ;
      RECT  2.44 1.305 2.53 1.33 ;
      RECT  2.44 1.33 2.825 1.42 ;
      RECT  2.735 1.42 2.825 1.65 ;
      RECT  3.405 0.785 3.835 0.895 ;
      RECT  3.405 0.895 3.495 1.245 ;
      RECT  2.39 0.235 2.71 0.355 ;
      RECT  2.62 0.355 2.71 1.15 ;
      RECT  2.62 1.15 3.035 1.24 ;
      RECT  2.945 1.24 3.035 1.245 ;
      RECT  2.945 1.245 3.495 1.335 ;
      RECT  2.195 0.32 2.285 0.93 ;
      RECT  1.825 0.93 2.285 0.955 ;
      RECT  1.825 0.955 2.35 1.125 ;
  END
END SEN_FDPQB_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPQB_D_4
#      Description : "D-Flip Flop, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPQB_D_4
  CLASS CORE ;
  FOREIGN SEN_FDPQB_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0375 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.48 1.05 0.915 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.58 0.44 4.305 0.56 ;
      RECT  4.15 0.56 4.25 1.11 ;
      RECT  3.55 1.11 4.3 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.44 0.185 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.825 1.48 0.995 1.75 ;
      RECT  1.975 1.575 2.095 1.75 ;
      RECT  3.085 1.47 3.205 1.75 ;
      RECT  3.35 1.45 3.52 1.75 ;
      RECT  3.895 1.415 4.015 1.75 ;
      RECT  4.415 1.215 4.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  3.9 0.05 4.02 0.35 ;
      RECT  0.85 0.05 0.97 0.36 ;
      RECT  1.91 0.05 2.03 0.38 ;
      RECT  2.89 0.05 3.01 0.38 ;
      RECT  0.065 0.05 0.185 0.385 ;
      RECT  3.38 0.05 3.5 0.385 ;
      RECT  4.415 0.05 4.535 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.36 0.215 1.8 0.335 ;
      RECT  1.71 0.335 1.8 0.75 ;
      RECT  1.48 0.75 2.105 0.84 ;
      RECT  2.015 0.67 2.105 0.75 ;
      RECT  1.48 0.84 1.57 1.125 ;
      RECT  2.185 0.21 2.285 0.38 ;
      RECT  2.195 0.38 2.285 0.93 ;
      RECT  1.825 0.93 2.285 0.955 ;
      RECT  1.825 0.955 2.35 1.125 ;
      RECT  3.15 0.21 3.27 0.385 ;
      RECT  3.15 0.385 3.25 0.785 ;
      RECT  2.82 0.785 3.25 0.905 ;
      RECT  3.12 0.905 3.21 1.16 ;
      RECT  0.34 0.19 0.46 0.47 ;
      RECT  0.34 0.47 0.58 0.64 ;
      RECT  0.34 0.64 0.43 1.3 ;
      RECT  0.34 1.3 1.21 1.39 ;
      RECT  1.12 1.39 1.21 1.395 ;
      RECT  0.34 1.39 0.43 1.61 ;
      RECT  1.12 1.395 2.35 1.485 ;
      RECT  2.26 1.485 2.35 1.545 ;
      RECT  2.26 1.545 2.58 1.645 ;
      RECT  2.375 0.625 2.53 0.795 ;
      RECT  2.44 0.795 2.53 1.215 ;
      RECT  1.23 0.45 1.62 0.62 ;
      RECT  1.23 0.62 1.32 1.085 ;
      RECT  1.23 1.085 1.39 1.105 ;
      RECT  0.605 0.19 0.76 0.36 ;
      RECT  0.67 0.36 0.76 1.105 ;
      RECT  0.565 1.105 1.39 1.21 ;
      RECT  1.3 1.21 1.39 1.215 ;
      RECT  1.3 1.215 2.53 1.305 ;
      RECT  2.44 1.305 2.53 1.33 ;
      RECT  2.44 1.33 2.825 1.42 ;
      RECT  2.735 1.42 2.825 1.645 ;
      RECT  3.34 0.745 4.01 0.855 ;
      RECT  3.34 0.855 3.43 1.27 ;
      RECT  2.405 0.235 2.71 0.355 ;
      RECT  2.62 0.355 2.71 1.15 ;
      RECT  2.62 1.15 3.005 1.24 ;
      RECT  2.915 1.24 3.005 1.27 ;
      RECT  2.915 1.27 3.43 1.36 ;
  END
END SEN_FDPQB_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBQ_1
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBQ_1
  CLASS CORE ;
  FOREIGN SEN_FDPRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.405 0.755 3.505 1.205 ;
      RECT  3.405 1.205 4.135 1.235 ;
      RECT  2.875 0.71 3.05 0.925 ;
      RECT  2.95 0.925 3.05 1.235 ;
      RECT  2.95 1.235 4.135 1.305 ;
      RECT  2.95 1.305 3.505 1.335 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.072 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.73 0.89 0.87 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.31 5.325 0.49 ;
      RECT  5.15 0.49 5.25 1.11 ;
      RECT  5.15 1.11 5.325 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.155 0.51 4.55 0.69 ;
      RECT  1.865 0.55 2.05 0.65 ;
      RECT  1.935 0.65 2.05 0.98 ;
      RECT  0.75 0.51 0.85 0.69 ;
      RECT  0.505 0.69 0.85 0.78 ;
      RECT  0.505 0.78 0.63 0.96 ;
      LAYER M2 ;
      RECT  0.68 0.55 4.495 0.65 ;
      LAYER V1 ;
      RECT  4.355 0.55 4.455 0.65 ;
      RECT  1.905 0.55 2.005 0.65 ;
      RECT  0.75 0.55 0.85 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0753 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.45 0.46 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  1.88 1.47 2.0 1.75 ;
      RECT  2.145 1.45 2.265 1.75 ;
      RECT  2.945 1.44 3.065 1.75 ;
      RECT  4.31 1.61 4.48 1.75 ;
      RECT  4.945 1.415 5.065 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  2.085 0.05 2.255 0.28 ;
      RECT  2.91 0.05 3.08 0.305 ;
      RECT  4.425 0.05 4.545 0.385 ;
      RECT  0.35 0.05 0.46 0.39 ;
      RECT  4.95 0.05 5.06 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.55 0.14 1.325 0.23 ;
      RECT  0.55 0.23 0.64 0.51 ;
      RECT  1.21 0.23 1.325 1.08 ;
      RECT  0.245 0.51 0.64 0.6 ;
      RECT  0.245 0.6 0.345 0.99 ;
      RECT  1.21 1.08 2.23 1.18 ;
      RECT  3.33 0.19 3.89 0.29 ;
      RECT  3.33 0.29 3.43 0.395 ;
      RECT  2.615 0.365 2.825 0.395 ;
      RECT  2.615 0.395 3.43 0.485 ;
      RECT  2.615 0.485 2.715 1.055 ;
      RECT  2.615 1.055 2.81 1.175 ;
      RECT  0.83 0.32 1.12 0.42 ;
      RECT  1.03 0.42 1.12 1.38 ;
      RECT  0.83 1.38 1.12 1.48 ;
      RECT  1.415 0.37 2.525 0.46 ;
      RECT  1.415 0.46 1.515 0.99 ;
      RECT  2.425 0.46 2.525 1.17 ;
      RECT  3.18 0.575 3.35 0.665 ;
      RECT  3.18 0.665 3.315 1.145 ;
      RECT  4.675 0.235 4.795 0.785 ;
      RECT  4.11 0.785 4.795 0.895 ;
      RECT  4.675 0.895 4.795 1.145 ;
      RECT  3.595 0.44 3.7 1.01 ;
      RECT  3.595 1.01 4.45 1.11 ;
      RECT  4.36 1.11 4.45 1.235 ;
      RECT  4.36 1.235 5.05 1.325 ;
      RECT  4.95 0.755 5.05 1.235 ;
      RECT  1.21 1.27 2.705 1.36 ;
      RECT  1.685 1.36 1.79 1.56 ;
      RECT  1.21 1.36 1.3 1.57 ;
      RECT  2.605 1.36 2.705 1.66 ;
      RECT  0.09 0.21 0.19 0.34 ;
      RECT  0.055 0.34 0.19 0.43 ;
      RECT  0.055 0.43 0.155 1.27 ;
      RECT  0.055 1.27 0.64 1.36 ;
      RECT  0.55 1.36 0.64 1.57 ;
      RECT  0.55 1.57 1.3 1.66 ;
      RECT  4.04 1.415 4.75 1.52 ;
  END
END SEN_FDPRBQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBQ_2
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBQ_2
  CLASS CORE ;
  FOREIGN SEN_FDPRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.85 0.89 ;
      RECT  3.95 0.89 4.05 1.05 ;
      RECT  4.75 0.89 4.85 1.09 ;
      RECT  3.83 1.05 4.05 1.15 ;
      RECT  3.83 1.15 3.93 1.25 ;
      RECT  3.15 0.51 3.25 0.71 ;
      RECT  3.15 0.71 3.305 0.95 ;
      RECT  3.215 0.95 3.305 1.25 ;
      RECT  3.215 1.25 3.93 1.34 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.087 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.045 ;
      RECT  0.28 1.045 0.45 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0555 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.31 6.275 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.51 5.25 0.71 ;
      RECT  5.15 0.71 5.45 0.89 ;
      RECT  2.065 0.51 2.165 0.71 ;
      RECT  2.065 0.71 2.25 0.925 ;
      RECT  0.15 0.51 0.25 0.93 ;
      LAYER M2 ;
      RECT  0.11 0.55 5.29 0.65 ;
      LAYER V1 ;
      RECT  5.15 0.55 5.25 0.65 ;
      RECT  2.065 0.55 2.165 0.65 ;
      RECT  0.15 0.55 0.25 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.078 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.385 0.185 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.615 1.43 0.735 1.75 ;
      RECT  2.065 1.47 2.195 1.75 ;
      RECT  2.43 1.47 2.56 1.75 ;
      RECT  3.24 1.43 3.41 1.75 ;
      RECT  3.785 1.62 3.955 1.75 ;
      RECT  5.11 1.615 5.28 1.75 ;
      RECT  5.895 1.44 6.015 1.75 ;
      RECT  6.415 1.21 6.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  3.785 0.05 3.955 0.185 ;
      RECT  3.225 0.05 3.395 0.2 ;
      RECT  1.045 0.05 1.215 0.28 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  2.435 0.05 2.545 0.43 ;
      RECT  6.415 0.05 6.535 0.59 ;
      RECT  5.375 0.05 5.495 0.62 ;
      RECT  5.895 0.05 6.015 0.65 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.635 0.14 3.05 0.29 ;
      RECT  2.635 0.29 4.665 0.295 ;
      RECT  4.155 0.195 4.665 0.29 ;
      RECT  2.635 0.295 4.245 0.31 ;
      RECT  2.94 0.31 4.245 0.4 ;
      RECT  2.94 0.4 3.05 1.065 ;
      RECT  2.94 1.065 3.125 1.185 ;
      RECT  1.815 0.33 2.345 0.42 ;
      RECT  2.255 0.42 2.345 0.52 ;
      RECT  1.815 0.42 1.905 0.795 ;
      RECT  2.255 0.52 2.85 0.61 ;
      RECT  2.73 0.61 2.85 1.2 ;
      RECT  1.67 0.795 1.905 0.965 ;
      RECT  0.54 0.37 1.49 0.47 ;
      RECT  0.54 0.47 0.65 1.225 ;
      RECT  0.54 1.225 1.295 1.245 ;
      RECT  0.325 1.245 1.295 1.34 ;
      RECT  0.325 1.34 0.445 1.595 ;
      RECT  4.31 0.5 5.03 0.59 ;
      RECT  4.94 0.59 5.03 1.24 ;
      RECT  4.02 1.24 6.05 1.34 ;
      RECT  5.95 0.745 6.05 1.24 ;
      RECT  3.485 0.495 4.22 0.615 ;
      RECT  3.485 0.615 3.575 1.05 ;
      RECT  3.485 1.05 3.695 1.16 ;
      RECT  0.755 0.56 0.96 0.68 ;
      RECT  0.755 0.68 0.845 1.025 ;
      RECT  0.755 1.025 1.07 1.135 ;
      RECT  1.415 0.56 1.725 0.68 ;
      RECT  1.415 0.68 1.515 0.785 ;
      RECT  0.935 0.785 1.515 0.895 ;
      RECT  1.415 0.895 1.515 1.055 ;
      RECT  1.415 1.055 2.415 1.175 ;
      RECT  1.415 1.175 1.525 1.365 ;
      RECT  5.625 0.44 5.745 1.035 ;
      RECT  5.12 1.035 5.745 1.145 ;
      RECT  1.85 1.29 2.845 1.38 ;
      RECT  1.85 1.38 1.96 1.455 ;
      RECT  2.755 1.38 2.845 1.52 ;
      RECT  0.855 1.455 1.96 1.57 ;
      RECT  2.755 1.52 3.06 1.63 ;
      RECT  4.815 1.43 5.68 1.525 ;
      RECT  3.5 1.43 4.51 1.53 ;
  END
END SEN_FDPRBQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBQ_4
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBQ_4
  CLASS CORE ;
  FOREIGN SEN_FDPRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.125 0.63 5.325 0.74 ;
      RECT  5.235 0.74 5.325 1.255 ;
      RECT  3.615 0.805 3.725 1.035 ;
      RECT  3.615 1.035 3.85 1.125 ;
      RECT  3.75 1.125 3.85 1.255 ;
      RECT  3.75 1.255 5.325 1.345 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1197 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0792 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.51 7.45 0.69 ;
      RECT  7.15 0.69 7.25 1.11 ;
      RECT  6.75 1.11 7.475 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.465 6.05 0.89 ;
      RECT  1.95 0.71 2.125 0.965 ;
      RECT  0.735 0.71 0.865 1.22 ;
      LAYER M2 ;
      RECT  0.71 0.75 6.09 0.85 ;
      LAYER V1 ;
      RECT  5.95 0.75 6.05 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.325 0.185 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.605 1.53 0.725 1.75 ;
      RECT  1.85 1.425 1.98 1.75 ;
      RECT  2.415 1.415 2.535 1.75 ;
      RECT  2.945 1.35 3.065 1.75 ;
      RECT  3.735 1.435 3.855 1.75 ;
      RECT  4.255 1.435 4.375 1.75 ;
      RECT  5.845 1.62 6.015 1.75 ;
      RECT  6.555 1.42 6.675 1.75 ;
      RECT  7.075 1.385 7.195 1.75 ;
      RECT  7.595 1.21 7.715 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  0.86 0.05 1.03 0.19 ;
      RECT  2.125 0.05 2.245 0.225 ;
      RECT  2.665 0.05 2.785 0.225 ;
      RECT  3.185 0.05 3.305 0.225 ;
      RECT  3.725 0.05 3.845 0.225 ;
      RECT  4.255 0.05 4.375 0.37 ;
      RECT  6.035 0.05 6.155 0.375 ;
      RECT  7.075 0.05 7.195 0.42 ;
      RECT  7.595 0.05 7.715 0.59 ;
      RECT  6.555 0.05 6.66 0.625 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.405 0.21 2.505 0.315 ;
      RECT  2.405 0.315 3.905 0.405 ;
      RECT  3.815 0.405 3.905 0.795 ;
      RECT  2.74 0.405 2.83 1.055 ;
      RECT  3.815 0.795 4.33 0.905 ;
      RECT  1.695 1.055 2.83 1.155 ;
      RECT  2.66 1.155 2.83 1.185 ;
      RECT  0.31 0.28 1.28 0.38 ;
      RECT  0.955 0.38 1.045 1.33 ;
      RECT  0.31 1.33 1.045 1.365 ;
      RECT  0.31 1.365 1.27 1.44 ;
      RECT  0.955 1.44 1.27 1.475 ;
      RECT  1.37 0.315 2.315 0.405 ;
      RECT  2.215 0.405 2.315 0.745 ;
      RECT  4.515 0.4 5.22 0.46 ;
      RECT  3.995 0.46 5.22 0.505 ;
      RECT  3.995 0.505 4.635 0.57 ;
      RECT  3.995 0.57 4.115 0.655 ;
      RECT  4.515 0.57 4.635 0.985 ;
      RECT  4.515 0.985 5.145 1.035 ;
      RECT  3.945 1.035 5.145 1.16 ;
      RECT  0.075 0.375 0.195 0.47 ;
      RECT  0.075 0.47 0.765 0.59 ;
      RECT  1.53 0.495 1.63 0.605 ;
      RECT  1.14 0.605 1.63 0.695 ;
      RECT  1.14 0.695 1.25 1.15 ;
      RECT  1.14 1.15 1.32 1.25 ;
      RECT  3.13 0.495 3.63 0.615 ;
      RECT  3.13 0.615 3.23 0.885 ;
      RECT  3.13 0.885 3.49 0.985 ;
      RECT  3.4 0.985 3.49 1.24 ;
      RECT  3.4 1.24 3.625 1.36 ;
      RECT  1.75 0.51 1.85 0.85 ;
      RECT  1.405 0.85 1.85 0.965 ;
      RECT  6.49 0.785 7.06 0.895 ;
      RECT  6.49 0.895 6.58 1.24 ;
      RECT  4.73 0.21 5.705 0.31 ;
      RECT  5.615 0.31 5.705 1.24 ;
      RECT  5.415 1.24 6.58 1.33 ;
      RECT  5.415 1.33 5.505 1.44 ;
      RECT  4.73 1.44 5.505 1.56 ;
      RECT  5.795 0.965 5.895 1.045 ;
      RECT  5.795 1.045 6.4 1.15 ;
      RECT  6.285 0.21 6.4 1.045 ;
      RECT  5.415 0.51 5.525 1.06 ;
      RECT  2.94 0.495 3.04 1.085 ;
      RECT  2.94 1.085 3.31 1.175 ;
      RECT  3.205 1.175 3.31 1.44 ;
      RECT  1.435 1.245 2.365 1.335 ;
      RECT  2.115 1.335 2.365 1.34 ;
      RECT  1.435 1.335 1.53 1.45 ;
      RECT  2.115 1.34 2.235 1.605 ;
      RECT  1.36 1.45 1.53 1.565 ;
      RECT  0.815 1.565 1.53 1.57 ;
      RECT  0.815 1.57 1.455 1.66 ;
      RECT  5.595 1.42 6.33 1.53 ;
      RECT  5.595 1.53 5.705 1.615 ;
      LAYER M2 ;
      RECT  1.71 0.55 5.56 0.65 ;
      RECT  1.14 1.15 3.345 1.25 ;
      LAYER V1 ;
      RECT  1.75 0.55 1.85 0.65 ;
      RECT  3.13 0.55 3.23 0.65 ;
      RECT  5.42 0.55 5.52 0.65 ;
      RECT  1.18 1.15 1.28 1.25 ;
      RECT  3.205 1.15 3.305 1.25 ;
  END
END SEN_FDPRBQ_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBQ_D_1
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FDPRBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.52 0.69 ;
      RECT  4.35 0.69 4.45 1.095 ;
      RECT  4.35 1.095 4.52 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 3.65 0.71 ;
      RECT  3.35 0.71 3.65 0.89 ;
      RECT  2.135 0.67 2.295 0.965 ;
      LAYER M2 ;
      RECT  2.155 0.75 3.49 0.85 ;
      LAYER V1 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  2.195 0.75 2.295 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.042 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.84 1.45 0.97 1.75 ;
      RECT  1.795 1.63 1.965 1.75 ;
      RECT  2.29 1.63 2.46 1.75 ;
      RECT  3.455 1.295 3.585 1.75 ;
      RECT  4.17 1.21 4.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.3 0.05 2.47 0.185 ;
      RECT  3.34 0.05 3.51 0.19 ;
      RECT  0.82 0.05 0.99 0.2 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  4.145 0.05 4.275 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.22 0.16 2.165 0.25 ;
      RECT  2.075 0.25 2.165 0.295 ;
      RECT  1.22 0.25 1.335 0.3 ;
      RECT  2.075 0.295 3.105 0.385 ;
      RECT  3.005 0.16 3.105 0.295 ;
      RECT  0.34 0.3 1.335 0.39 ;
      RECT  0.34 0.39 0.445 0.785 ;
      RECT  0.34 0.785 0.66 0.895 ;
      RECT  0.34 0.895 0.43 1.21 ;
      RECT  0.065 1.21 0.43 1.305 ;
      RECT  0.065 1.305 0.185 1.43 ;
      RECT  3.195 0.3 4.02 0.4 ;
      RECT  3.9 0.4 4.02 0.6 ;
      RECT  3.9 0.6 4.08 0.69 ;
      RECT  3.99 0.69 4.08 0.785 ;
      RECT  3.99 0.785 4.26 0.895 ;
      RECT  3.99 0.895 4.08 1.32 ;
      RECT  3.68 1.32 4.08 1.44 ;
      RECT  1.48 0.34 1.985 0.445 ;
      RECT  1.895 0.445 1.985 0.475 ;
      RECT  1.895 0.475 2.495 0.565 ;
      RECT  2.385 0.565 2.495 0.825 ;
      RECT  1.895 0.565 1.985 0.875 ;
      RECT  1.41 0.875 1.985 0.965 ;
      RECT  1.41 0.965 1.5 1.235 ;
      RECT  1.33 1.235 1.5 1.355 ;
      RECT  2.585 0.475 2.755 0.595 ;
      RECT  2.585 0.595 2.675 1.055 ;
      RECT  1.8 1.055 2.705 1.145 ;
      RECT  2.6 1.145 2.705 1.3 ;
      RECT  2.845 0.48 3.085 0.6 ;
      RECT  2.98 0.6 3.085 1.115 ;
      RECT  2.98 1.115 3.9 1.205 ;
      RECT  3.79 0.84 3.9 1.115 ;
      RECT  2.98 1.205 3.1 1.46 ;
      RECT  2.765 0.695 2.885 0.865 ;
      RECT  2.795 0.865 2.885 1.45 ;
      RECT  0.545 0.485 1.25 0.605 ;
      RECT  1.15 0.605 1.25 0.695 ;
      RECT  1.15 0.695 1.78 0.785 ;
      RECT  1.67 0.585 1.78 0.695 ;
      RECT  1.15 0.785 1.3 0.925 ;
      RECT  1.15 0.925 1.24 1.24 ;
      RECT  0.55 1.24 1.24 1.36 ;
      RECT  1.15 1.36 1.24 1.45 ;
      RECT  1.15 1.45 2.885 1.54 ;
      RECT  2.795 1.54 2.885 1.55 ;
      RECT  2.795 1.55 3.25 1.64 ;
      RECT  1.59 1.235 2.25 1.355 ;
  END
END SEN_FDPRBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBQ_D_1P5
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBQ_D_1P5
  CLASS CORE ;
  FOREIGN SEN_FDPRBQ_D_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.935 ;
      RECT  0.07 0.935 0.25 1.105 ;
      RECT  0.15 1.105 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.08 0.2 4.255 0.32 ;
      RECT  4.15 0.32 4.255 0.51 ;
      RECT  4.15 0.51 4.45 0.69 ;
      RECT  4.35 0.69 4.45 1.11 ;
      RECT  4.15 1.11 4.45 1.29 ;
      RECT  4.15 1.29 4.25 1.385 ;
      RECT  4.065 1.385 4.25 1.505 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.085 0.14 3.135 0.23 ;
      RECT  3.045 0.23 3.135 0.31 ;
      RECT  2.085 0.23 2.175 0.395 ;
      RECT  3.045 0.31 3.25 0.4 ;
      RECT  1.78 0.395 2.175 0.485 ;
      RECT  3.15 0.4 3.25 0.61 ;
      RECT  1.78 0.485 1.89 0.635 ;
      RECT  3.15 0.61 3.855 0.7 ;
      RECT  3.745 0.7 3.855 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.051 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.385 0.19 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.785 1.43 0.905 1.75 ;
      RECT  2.12 1.64 2.29 1.75 ;
      RECT  3.305 1.225 3.425 1.75 ;
      RECT  3.835 1.405 3.955 1.75 ;
      RECT  4.385 1.38 4.505 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  3.225 0.05 3.345 0.22 ;
      RECT  1.875 0.05 1.995 0.305 ;
      RECT  3.82 0.05 3.99 0.325 ;
      RECT  0.06 0.05 0.18 0.42 ;
      RECT  0.765 0.05 0.885 0.42 ;
      RECT  4.385 0.05 4.505 0.42 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.17 0.24 1.66 0.36 ;
      RECT  1.55 0.36 1.66 0.74 ;
      RECT  1.345 0.74 2.2 0.83 ;
      RECT  2.1 0.615 2.2 0.74 ;
      RECT  1.345 0.83 1.435 1.17 ;
      RECT  1.195 1.17 1.435 1.275 ;
      RECT  2.47 0.32 2.955 0.41 ;
      RECT  2.865 0.41 2.955 0.79 ;
      RECT  2.865 0.79 3.605 0.865 ;
      RECT  2.87 0.865 3.605 0.895 ;
      RECT  2.87 0.895 2.96 1.2 ;
      RECT  2.84 1.2 2.96 1.37 ;
      RECT  2.265 0.32 2.38 0.49 ;
      RECT  2.29 0.49 2.38 0.92 ;
      RECT  1.58 0.92 2.565 1.01 ;
      RECT  2.46 1.01 2.565 1.19 ;
      RECT  3.35 0.415 4.045 0.515 ;
      RECT  3.955 0.515 4.045 0.78 ;
      RECT  3.955 0.78 4.24 0.89 ;
      RECT  3.955 0.89 4.045 1.01 ;
      RECT  3.115 1.01 4.045 1.13 ;
      RECT  3.565 1.13 3.685 1.635 ;
      RECT  1.355 0.46 1.46 0.55 ;
      RECT  1.15 0.55 1.46 0.64 ;
      RECT  1.15 0.64 1.255 0.99 ;
      RECT  0.505 0.21 0.645 0.38 ;
      RECT  0.53 0.38 0.645 0.99 ;
      RECT  0.53 0.99 1.255 1.08 ;
      RECT  0.53 1.08 0.645 1.16 ;
      RECT  2.66 0.5 2.775 0.91 ;
      RECT  2.66 0.91 2.78 1.08 ;
      RECT  2.66 1.08 2.75 1.28 ;
      RECT  1.75 1.28 2.75 1.365 ;
      RECT  0.315 0.465 0.44 0.645 ;
      RECT  0.34 0.645 0.44 1.25 ;
      RECT  0.34 1.25 1.095 1.34 ;
      RECT  1.005 1.34 1.095 1.365 ;
      RECT  0.34 1.34 0.45 1.54 ;
      RECT  1.005 1.365 2.75 1.37 ;
      RECT  1.005 1.37 1.84 1.465 ;
      RECT  1.525 1.1 2.185 1.19 ;
      RECT  1.525 1.19 1.635 1.275 ;
      RECT  1.935 1.46 3.075 1.55 ;
      RECT  1.935 1.55 2.03 1.555 ;
      RECT  1.545 1.555 2.03 1.66 ;
  END
END SEN_FDPRBQ_D_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBQ_D_2
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FDPRBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.325 0.51 4.65 0.69 ;
      RECT  4.55 0.69 4.65 1.11 ;
      RECT  4.35 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.5 0.51 3.6 0.71 ;
      RECT  3.3 0.71 3.6 0.89 ;
      RECT  2.085 0.67 2.245 0.965 ;
      LAYER M2 ;
      RECT  2.105 0.75 3.44 0.85 ;
      LAYER V1 ;
      RECT  3.3 0.75 3.4 0.85 ;
      RECT  2.145 0.75 2.245 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.79 1.45 0.92 1.75 ;
      RECT  1.745 1.63 1.915 1.75 ;
      RECT  2.24 1.63 2.41 1.75 ;
      RECT  3.405 1.295 3.535 1.75 ;
      RECT  4.12 1.21 4.23 1.75 ;
      RECT  4.62 1.41 4.75 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  2.25 0.05 2.42 0.185 ;
      RECT  3.29 0.05 3.46 0.19 ;
      RECT  0.77 0.05 0.94 0.2 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  4.1 0.05 4.23 0.39 ;
      RECT  4.62 0.05 4.75 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.21 0.16 2.115 0.25 ;
      RECT  2.025 0.25 2.115 0.295 ;
      RECT  1.21 0.25 1.32 0.3 ;
      RECT  2.025 0.295 3.055 0.385 ;
      RECT  2.955 0.16 3.055 0.295 ;
      RECT  0.34 0.19 0.445 0.3 ;
      RECT  0.34 0.3 1.32 0.39 ;
      RECT  0.34 0.39 0.445 0.785 ;
      RECT  0.34 0.785 0.64 0.895 ;
      RECT  0.34 0.895 0.43 1.21 ;
      RECT  0.065 1.21 0.43 1.305 ;
      RECT  0.065 1.305 0.185 1.43 ;
      RECT  3.145 0.3 3.97 0.4 ;
      RECT  3.85 0.4 3.97 0.6 ;
      RECT  3.85 0.6 4.03 0.69 ;
      RECT  3.94 0.69 4.03 0.785 ;
      RECT  3.94 0.785 4.46 0.895 ;
      RECT  3.94 0.895 4.03 1.32 ;
      RECT  3.63 1.32 4.03 1.44 ;
      RECT  1.435 0.34 1.935 0.445 ;
      RECT  1.845 0.445 1.935 0.475 ;
      RECT  1.845 0.475 2.445 0.565 ;
      RECT  2.335 0.565 2.445 0.825 ;
      RECT  1.845 0.565 1.935 0.875 ;
      RECT  1.36 0.875 1.935 0.965 ;
      RECT  1.36 0.965 1.45 1.21 ;
      RECT  1.32 1.21 1.45 1.4 ;
      RECT  2.535 0.475 2.705 0.595 ;
      RECT  2.535 0.595 2.625 1.055 ;
      RECT  1.75 1.055 2.655 1.145 ;
      RECT  2.55 1.145 2.655 1.3 ;
      RECT  2.795 0.48 3.035 0.6 ;
      RECT  2.93 0.6 3.035 1.115 ;
      RECT  2.93 1.115 3.85 1.205 ;
      RECT  3.74 0.835 3.85 1.115 ;
      RECT  2.93 1.205 3.05 1.46 ;
      RECT  2.715 0.695 2.835 0.865 ;
      RECT  2.745 0.865 2.835 1.45 ;
      RECT  1.565 1.45 2.835 1.54 ;
      RECT  2.745 1.54 2.835 1.55 ;
      RECT  1.565 1.54 1.655 1.57 ;
      RECT  2.745 1.55 3.2 1.64 ;
      RECT  0.535 0.5 1.24 0.62 ;
      RECT  0.535 0.62 0.63 0.695 ;
      RECT  1.14 0.62 1.24 0.695 ;
      RECT  1.14 0.695 1.73 0.785 ;
      RECT  1.62 0.585 1.73 0.695 ;
      RECT  1.14 0.785 1.265 0.955 ;
      RECT  1.14 0.955 1.23 1.24 ;
      RECT  0.525 1.01 0.645 1.24 ;
      RECT  0.525 1.24 1.23 1.36 ;
      RECT  1.14 1.36 1.23 1.57 ;
      RECT  1.14 1.57 1.655 1.66 ;
      RECT  1.54 1.235 2.2 1.355 ;
  END
END SEN_FDPRBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBQ_D_3
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBQ_D_3
  CLASS CORE ;
  FOREIGN SEN_FDPRBQ_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.925 ;
      RECT  0.075 0.925 0.25 1.095 ;
      RECT  0.15 1.095 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.08 0.2 4.255 0.32 ;
      RECT  4.15 0.32 4.255 0.51 ;
      RECT  4.15 0.51 4.745 0.69 ;
      RECT  4.55 0.69 4.65 1.11 ;
      RECT  4.15 1.11 4.745 1.29 ;
      RECT  4.15 1.29 4.25 1.385 ;
      RECT  4.05 1.385 4.25 1.505 ;
    END
    ANTENNADIFFAREA 0.358 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.085 0.14 3.135 0.23 ;
      RECT  3.045 0.23 3.135 0.31 ;
      RECT  2.085 0.23 2.175 0.395 ;
      RECT  3.045 0.31 3.25 0.4 ;
      RECT  1.78 0.395 2.175 0.485 ;
      RECT  3.15 0.4 3.25 0.61 ;
      RECT  1.78 0.485 1.89 0.65 ;
      RECT  3.15 0.61 3.855 0.7 ;
      RECT  3.745 0.7 3.855 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.38 0.19 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.785 1.43 0.905 1.75 ;
      RECT  2.12 1.64 2.29 1.75 ;
      RECT  3.305 1.225 3.425 1.75 ;
      RECT  3.835 1.41 3.955 1.75 ;
      RECT  4.365 1.385 4.485 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  3.225 0.05 3.345 0.22 ;
      RECT  1.875 0.05 1.995 0.305 ;
      RECT  3.82 0.05 3.99 0.325 ;
      RECT  0.765 0.05 0.885 0.41 ;
      RECT  0.06 0.05 0.18 0.415 ;
      RECT  4.365 0.05 4.485 0.415 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.175 0.24 1.66 0.36 ;
      RECT  1.55 0.36 1.66 0.74 ;
      RECT  1.345 0.74 2.2 0.83 ;
      RECT  2.1 0.625 2.2 0.74 ;
      RECT  1.345 0.83 1.435 1.17 ;
      RECT  1.2 1.17 1.435 1.275 ;
      RECT  2.49 0.32 2.955 0.41 ;
      RECT  2.865 0.41 2.955 0.79 ;
      RECT  2.865 0.79 3.635 0.865 ;
      RECT  2.87 0.865 3.635 0.895 ;
      RECT  2.87 0.895 2.96 1.2 ;
      RECT  2.84 1.2 2.96 1.37 ;
      RECT  2.265 0.32 2.38 0.49 ;
      RECT  2.29 0.49 2.38 0.92 ;
      RECT  1.58 0.92 2.565 1.01 ;
      RECT  2.46 1.01 2.565 1.19 ;
      RECT  3.35 0.415 4.045 0.52 ;
      RECT  3.955 0.52 4.045 0.785 ;
      RECT  3.955 0.785 4.44 0.895 ;
      RECT  3.955 0.895 4.045 1.01 ;
      RECT  3.115 1.01 4.045 1.13 ;
      RECT  3.565 1.13 3.685 1.635 ;
      RECT  1.355 0.46 1.46 0.55 ;
      RECT  1.15 0.55 1.46 0.64 ;
      RECT  1.15 0.64 1.255 0.99 ;
      RECT  0.485 0.21 0.645 0.38 ;
      RECT  0.53 0.38 0.645 0.99 ;
      RECT  0.53 0.99 1.255 1.08 ;
      RECT  0.53 1.08 0.645 1.16 ;
      RECT  2.66 0.5 2.775 0.91 ;
      RECT  2.66 0.91 2.78 1.08 ;
      RECT  2.66 1.08 2.75 1.28 ;
      RECT  1.75 1.28 2.75 1.365 ;
      RECT  0.315 0.475 0.44 0.645 ;
      RECT  0.34 0.645 0.44 1.25 ;
      RECT  0.34 1.25 1.095 1.34 ;
      RECT  1.005 1.34 1.095 1.365 ;
      RECT  0.34 1.34 0.45 1.54 ;
      RECT  1.005 1.365 2.75 1.37 ;
      RECT  1.005 1.37 1.84 1.465 ;
      RECT  1.53 1.1 2.19 1.19 ;
      RECT  1.53 1.19 1.635 1.275 ;
      RECT  1.935 1.46 3.075 1.55 ;
      RECT  1.935 1.55 2.03 1.555 ;
      RECT  1.545 1.555 2.03 1.66 ;
  END
END SEN_FDPRBQ_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBQ_D_4
#      Description : "D-Flip Flop, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FDPRBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.325 0.51 5.05 0.69 ;
      RECT  4.95 0.69 5.05 1.11 ;
      RECT  4.35 1.11 5.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.5 0.51 3.6 0.71 ;
      RECT  3.3 0.71 3.6 0.89 ;
      RECT  2.085 0.67 2.245 0.965 ;
      LAYER M2 ;
      RECT  2.105 0.75 3.44 0.85 ;
      LAYER V1 ;
      RECT  3.3 0.75 3.4 0.85 ;
      RECT  2.145 0.75 2.245 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  0.79 1.45 0.92 1.75 ;
      RECT  1.745 1.63 1.915 1.75 ;
      RECT  2.24 1.63 2.41 1.75 ;
      RECT  3.405 1.295 3.535 1.75 ;
      RECT  4.12 1.21 4.225 1.75 ;
      RECT  4.62 1.41 4.75 1.75 ;
      RECT  5.16 1.21 5.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  2.25 0.05 2.42 0.185 ;
      RECT  3.29 0.05 3.46 0.19 ;
      RECT  0.77 0.05 0.94 0.2 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  4.1 0.05 4.23 0.39 ;
      RECT  4.62 0.05 4.75 0.4 ;
      RECT  5.16 0.05 5.28 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.21 0.16 2.115 0.25 ;
      RECT  2.025 0.25 2.115 0.295 ;
      RECT  1.21 0.25 1.32 0.3 ;
      RECT  2.025 0.295 3.055 0.385 ;
      RECT  2.955 0.16 3.055 0.295 ;
      RECT  0.34 0.19 0.445 0.3 ;
      RECT  0.34 0.3 1.32 0.39 ;
      RECT  0.34 0.39 0.445 0.785 ;
      RECT  0.34 0.785 0.61 0.895 ;
      RECT  0.34 0.895 0.43 1.21 ;
      RECT  0.065 1.21 0.43 1.305 ;
      RECT  0.065 1.305 0.185 1.43 ;
      RECT  3.145 0.3 3.97 0.4 ;
      RECT  3.85 0.4 3.97 0.53 ;
      RECT  3.85 0.53 4.03 0.62 ;
      RECT  3.94 0.62 4.03 0.785 ;
      RECT  3.94 0.785 4.84 0.895 ;
      RECT  3.94 0.895 4.03 1.32 ;
      RECT  3.63 1.32 4.03 1.44 ;
      RECT  1.43 0.34 1.935 0.445 ;
      RECT  1.845 0.445 1.935 0.475 ;
      RECT  1.845 0.475 2.445 0.565 ;
      RECT  2.335 0.565 2.445 0.825 ;
      RECT  1.845 0.565 1.935 0.875 ;
      RECT  1.36 0.875 1.935 0.965 ;
      RECT  1.36 0.965 1.45 1.21 ;
      RECT  1.32 1.21 1.45 1.385 ;
      RECT  2.535 0.475 2.705 0.595 ;
      RECT  2.535 0.595 2.625 1.055 ;
      RECT  1.735 1.055 2.655 1.145 ;
      RECT  2.55 1.145 2.655 1.3 ;
      RECT  2.795 0.48 3.035 0.6 ;
      RECT  2.93 0.6 3.035 1.115 ;
      RECT  2.93 1.115 3.85 1.205 ;
      RECT  3.74 0.73 3.85 1.115 ;
      RECT  2.93 1.205 3.05 1.46 ;
      RECT  2.715 0.695 2.835 0.865 ;
      RECT  2.745 0.865 2.835 1.45 ;
      RECT  1.565 1.45 2.835 1.54 ;
      RECT  2.745 1.54 2.835 1.55 ;
      RECT  1.565 1.54 1.655 1.57 ;
      RECT  2.745 1.55 3.2 1.64 ;
      RECT  0.535 0.5 1.24 0.62 ;
      RECT  0.535 0.62 0.63 0.695 ;
      RECT  1.14 0.62 1.24 0.695 ;
      RECT  1.14 0.695 1.73 0.785 ;
      RECT  1.62 0.585 1.73 0.695 ;
      RECT  1.14 0.785 1.265 0.955 ;
      RECT  1.14 0.955 1.23 1.24 ;
      RECT  0.525 1.01 0.645 1.24 ;
      RECT  0.525 1.24 1.23 1.36 ;
      RECT  1.14 1.36 1.23 1.57 ;
      RECT  1.14 1.57 1.655 1.66 ;
      RECT  1.54 1.235 2.2 1.355 ;
  END
END SEN_FDPRBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBSBQ_1
#      Description : "D-Flip Flop pos-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBSBQ_1
  CLASS CORE ;
  FOREIGN SEN_FDPRBSBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.69 0.51 2.85 0.755 ;
      RECT  2.75 0.755 2.85 1.54 ;
      RECT  2.75 1.54 3.16 1.64 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0729 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0387 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.31 5.45 1.315 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.45 0.47 3.55 0.91 ;
      RECT  1.41 0.75 1.69 0.99 ;
      LAYER M2 ;
      RECT  1.51 0.75 3.59 0.85 ;
      LAYER V1 ;
      RECT  3.45 0.75 3.55 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.45 0.71 ;
      RECT  4.35 0.71 4.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0561 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  1.19 1.47 1.36 1.75 ;
      RECT  2.01 1.47 2.18 1.75 ;
      RECT  3.44 1.615 3.61 1.75 ;
      RECT  3.97 1.43 4.08 1.75 ;
      RECT  4.505 1.43 4.625 1.75 ;
      RECT  5.08 1.2 5.2 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  1.52 0.05 1.63 0.3 ;
      RECT  2.02 0.05 2.19 0.305 ;
      RECT  3.55 0.05 3.67 0.38 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  4.27 0.05 4.39 0.42 ;
      RECT  5.045 0.05 5.165 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.89 0.17 1.43 0.26 ;
      RECT  0.89 0.26 0.98 0.34 ;
      RECT  1.34 0.26 1.43 0.395 ;
      RECT  1.34 0.395 2.42 0.485 ;
      RECT  2.31 0.485 2.42 1.58 ;
      RECT  2.51 0.215 2.73 0.335 ;
      RECT  2.51 0.335 2.6 0.91 ;
      RECT  2.51 0.91 2.645 1.41 ;
      RECT  2.82 0.215 3.04 0.335 ;
      RECT  2.94 0.335 3.04 1.2 ;
      RECT  3.76 0.34 3.945 0.46 ;
      RECT  3.76 0.46 3.86 1.04 ;
      RECT  3.76 1.04 4.41 1.16 ;
      RECT  1.75 0.575 2.22 0.68 ;
      RECT  2.12 0.68 2.22 1.28 ;
      RECT  0.89 1.28 2.22 1.38 ;
      RECT  0.89 1.38 0.98 1.52 ;
      RECT  1.775 1.38 1.895 1.525 ;
      RECT  0.52 0.555 0.61 1.52 ;
      RECT  0.52 1.52 0.98 1.625 ;
      RECT  4.035 0.31 4.135 0.935 ;
      RECT  1.15 0.47 1.25 0.98 ;
      RECT  3.245 0.83 3.355 1.065 ;
      RECT  3.245 1.065 3.55 1.155 ;
      RECT  3.46 1.155 3.55 1.25 ;
      RECT  3.46 1.25 4.895 1.34 ;
      RECT  4.775 0.165 4.895 1.25 ;
      RECT  0.93 0.43 1.06 1.08 ;
      RECT  0.93 1.08 1.67 1.19 ;
      RECT  5.085 0.675 5.185 1.105 ;
      RECT  0.7 0.31 0.8 1.395 ;
      RECT  3.145 1.29 3.34 1.405 ;
      RECT  3.25 1.405 3.34 1.435 ;
      RECT  3.25 1.435 3.88 1.525 ;
      RECT  0.34 0.245 0.43 1.415 ;
      LAYER M2 ;
      RECT  0.66 0.35 4.175 0.45 ;
      RECT  1.11 0.55 3.9 0.65 ;
      RECT  0.915 0.95 2.65 1.05 ;
      RECT  2.9 0.95 5.225 1.05 ;
      LAYER V1 ;
      RECT  0.7 0.35 0.8 0.45 ;
      RECT  4.035 0.35 4.135 0.45 ;
      RECT  1.15 0.55 1.25 0.65 ;
      RECT  3.76 0.55 3.86 0.65 ;
      RECT  0.955 0.95 1.055 1.05 ;
      RECT  2.51 0.95 2.61 1.05 ;
      RECT  2.94 0.95 3.04 1.05 ;
      RECT  5.085 0.95 5.185 1.05 ;
  END
END SEN_FDPRBSBQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBSBQ_2
#      Description : "D-Flip Flop pos-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBSBQ_2
  CLASS CORE ;
  FOREIGN SEN_FDPRBSBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.935 0.185 4.45 0.275 ;
      RECT  3.935 0.275 4.025 0.735 ;
      RECT  4.35 0.275 4.45 1.34 ;
      RECT  3.935 0.735 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0939 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.67 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.3 6.85 1.3 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.51 5.05 0.71 ;
      RECT  4.945 0.71 5.05 0.89 ;
      RECT  4.95 0.89 5.05 1.09 ;
      RECT  2.55 0.71 2.65 0.785 ;
      RECT  2.01 0.785 2.65 0.895 ;
      LAYER M2 ;
      RECT  2.51 0.75 5.085 0.85 ;
      LAYER V1 ;
      RECT  4.945 0.75 5.045 0.85 ;
      RECT  2.55 0.75 2.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0822 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0645 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.18 0.185 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  1.225 1.5 1.345 1.75 ;
      RECT  2.08 1.5 2.2 1.75 ;
      RECT  2.805 1.61 2.975 1.75 ;
      RECT  4.675 1.63 4.845 1.75 ;
      RECT  5.235 1.44 5.355 1.75 ;
      RECT  5.765 1.44 5.885 1.75 ;
      RECT  6.445 1.09 6.565 1.75 ;
      RECT  7.005 1.21 7.125 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  2.015 0.05 2.135 0.225 ;
      RECT  2.535 0.05 2.655 0.225 ;
      RECT  3.175 0.05 3.345 0.305 ;
      RECT  4.985 0.05 5.105 0.39 ;
      RECT  5.765 0.05 5.885 0.39 ;
      RECT  0.065 0.05 0.185 0.58 ;
      RECT  7.005 0.05 7.125 0.61 ;
      RECT  6.485 0.05 6.605 0.655 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.715 0.14 1.84 0.24 ;
      RECT  1.75 0.24 1.84 0.315 ;
      RECT  1.75 0.315 3.045 0.395 ;
      RECT  1.75 0.395 3.605 0.405 ;
      RECT  3.5 0.23 3.605 0.395 ;
      RECT  2.955 0.405 3.605 0.485 ;
      RECT  3.515 0.485 3.605 1.02 ;
      RECT  3.3 1.02 3.605 1.14 ;
      RECT  6.025 0.24 6.38 0.36 ;
      RECT  6.025 0.36 6.145 1.26 ;
      RECT  4.58 0.685 4.68 1.26 ;
      RECT  4.58 1.26 6.145 1.35 ;
      RECT  6.025 1.35 6.145 1.595 ;
      RECT  0.61 0.35 0.79 0.45 ;
      RECT  0.7 0.45 0.79 1.41 ;
      RECT  4.115 0.365 4.25 0.535 ;
      RECT  4.15 0.535 4.25 1.52 ;
      RECT  3.56 1.43 3.65 1.52 ;
      RECT  3.56 1.52 4.25 1.61 ;
      RECT  1.25 0.51 2.43 0.625 ;
      RECT  1.25 0.625 1.34 0.715 ;
      RECT  2.745 0.575 3.425 0.675 ;
      RECT  2.745 0.675 2.835 1.07 ;
      RECT  2.745 1.07 3.105 1.16 ;
      RECT  1.06 0.51 1.16 0.83 ;
      RECT  1.06 0.83 1.415 0.93 ;
      RECT  6.25 0.785 6.66 0.895 ;
      RECT  6.25 0.895 6.35 1.51 ;
      RECT  5.435 0.31 5.545 0.9 ;
      RECT  5.245 0.39 5.345 1.02 ;
      RECT  5.245 1.02 5.66 1.14 ;
      RECT  3.75 0.315 3.845 1.24 ;
      RECT  3.75 1.24 3.975 1.25 ;
      RECT  0.88 0.33 1.655 0.42 ;
      RECT  0.88 0.42 0.97 1.085 ;
      RECT  0.88 1.085 2.655 1.205 ;
      RECT  2.565 1.205 2.655 1.25 ;
      RECT  2.565 1.25 3.975 1.34 ;
      RECT  0.34 0.285 0.43 1.315 ;
      RECT  0.955 1.32 2.455 1.41 ;
      RECT  2.355 1.41 2.455 1.43 ;
      RECT  0.955 1.41 1.045 1.53 ;
      RECT  2.355 1.43 3.46 1.52 ;
      RECT  0.52 0.61 0.61 1.53 ;
      RECT  0.52 1.53 1.045 1.63 ;
      RECT  4.39 1.44 5.14 1.54 ;
      LAYER M2 ;
      RECT  0.61 0.35 5.58 0.45 ;
      RECT  1.02 0.55 5.385 0.65 ;
      RECT  4.11 1.35 6.39 1.45 ;
      LAYER V1 ;
      RECT  0.65 0.35 0.75 0.45 ;
      RECT  5.44 0.35 5.54 0.45 ;
      RECT  1.06 0.55 1.16 0.65 ;
      RECT  5.245 0.55 5.345 0.65 ;
      RECT  4.15 1.35 4.25 1.45 ;
      RECT  6.25 1.35 6.35 1.45 ;
  END
END SEN_FDPRBSBQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPRBSBQ_4
#      Description : "D-Flip Flop pos-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPRBSBQ_4
  CLASS CORE ;
  FOREIGN SEN_FDPRBSBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.315 0.14 4.945 0.25 ;
      RECT  4.855 0.25 4.945 0.71 ;
      RECT  4.855 0.71 5.05 0.8 ;
      RECT  4.95 0.8 5.05 1.11 ;
      RECT  4.83 1.11 5.05 1.29 ;
      RECT  4.83 1.29 4.935 1.325 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1215 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.675 0.25 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.965 0.51 8.65 0.69 ;
      RECT  8.35 0.69 8.45 1.11 ;
      RECT  7.95 1.11 8.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.71 5.45 0.91 ;
      RECT  5.15 0.91 5.45 1.09 ;
      RECT  2.975 0.69 3.075 1.005 ;
      RECT  2.5 1.005 3.075 1.115 ;
      LAYER M2 ;
      RECT  2.935 0.75 5.49 0.85 ;
      LAYER V1 ;
      RECT  5.35 0.75 5.45 0.85 ;
      RECT  2.975 0.75 3.075 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1143 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.71 7.05 0.91 ;
      RECT  6.75 0.91 7.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0762 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.215 0.185 1.75 ;
      RECT  0.0 1.75 9.0 1.85 ;
      RECT  1.5 1.62 1.67 1.75 ;
      RECT  2.09 1.62 2.26 1.75 ;
      RECT  2.725 1.63 2.895 1.75 ;
      RECT  3.295 1.63 3.465 1.75 ;
      RECT  5.165 1.615 5.345 1.75 ;
      RECT  6.21 1.425 6.33 1.75 ;
      RECT  6.775 1.425 6.895 1.75 ;
      RECT  7.725 1.15 7.845 1.75 ;
      RECT  8.26 1.38 8.38 1.75 ;
      RECT  8.81 1.21 8.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      RECT  2.495 0.05 2.605 0.285 ;
      RECT  3.025 0.05 3.145 0.285 ;
      RECT  3.595 0.05 3.715 0.33 ;
      RECT  7.035 0.05 7.155 0.395 ;
      RECT  8.275 0.05 8.395 0.42 ;
      RECT  5.375 0.05 5.495 0.44 ;
      RECT  6.53 0.05 6.635 0.44 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  8.81 0.05 8.93 0.59 ;
      RECT  7.755 0.05 7.875 0.64 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.34 0.14 0.98 0.23 ;
      RECT  0.865 0.23 0.98 0.385 ;
      RECT  0.34 0.23 0.445 1.345 ;
      RECT  5.625 0.14 6.44 0.24 ;
      RECT  5.625 0.24 5.745 0.41 ;
      RECT  6.35 0.24 6.44 0.53 ;
      RECT  6.35 0.53 6.895 0.62 ;
      RECT  6.775 0.31 6.895 0.53 ;
      RECT  1.115 0.14 2.405 0.25 ;
      RECT  2.315 0.25 2.405 0.375 ;
      RECT  2.315 0.375 3.175 0.42 ;
      RECT  2.315 0.42 4.02 0.465 ;
      RECT  3.085 0.465 4.02 0.51 ;
      RECT  3.68 0.51 4.02 0.53 ;
      RECT  3.68 0.53 3.77 1.255 ;
      RECT  3.555 1.255 3.77 1.36 ;
      RECT  7.245 0.24 7.66 0.36 ;
      RECT  7.245 0.36 7.365 1.245 ;
      RECT  5.035 0.15 5.135 0.53 ;
      RECT  5.035 0.53 5.69 0.62 ;
      RECT  5.6 0.62 5.69 1.245 ;
      RECT  5.6 1.245 7.365 1.335 ;
      RECT  7.245 1.335 7.365 1.6 ;
      RECT  0.535 0.35 0.74 0.45 ;
      RECT  0.535 0.45 0.625 1.44 ;
      RECT  0.535 1.44 0.73 1.61 ;
      RECT  6.08 0.35 6.26 0.45 ;
      RECT  6.16 0.45 6.26 0.925 ;
      RECT  1.07 0.35 1.52 0.46 ;
      RECT  1.615 0.34 2.225 0.46 ;
      RECT  2.135 0.46 2.225 0.56 ;
      RECT  2.135 0.56 2.875 0.665 ;
      RECT  2.755 0.665 2.875 0.82 ;
      RECT  4.115 0.4 4.765 0.49 ;
      RECT  4.115 0.49 4.235 0.595 ;
      RECT  4.64 0.49 4.765 0.605 ;
      RECT  4.64 0.605 4.74 1.48 ;
      RECT  4.07 1.48 4.74 1.6 ;
      RECT  1.045 0.55 1.225 0.65 ;
      RECT  1.125 0.65 1.225 0.825 ;
      RECT  1.125 0.825 1.845 0.935 ;
      RECT  3.29 0.6 3.59 0.7 ;
      RECT  3.5 0.7 3.59 0.95 ;
      RECT  3.41 0.95 3.59 1.145 ;
      RECT  7.535 0.785 8.24 0.895 ;
      RECT  7.535 0.895 7.635 1.51 ;
      RECT  5.89 0.39 5.99 1.04 ;
      RECT  5.89 1.04 6.65 1.155 ;
      RECT  3.885 0.95 4.285 1.09 ;
      RECT  3.165 0.79 3.305 1.17 ;
      RECT  0.75 0.54 0.85 1.21 ;
      RECT  0.75 1.21 0.92 1.32 ;
      RECT  0.83 1.32 0.92 1.44 ;
      RECT  0.83 1.44 3.21 1.53 ;
      RECT  4.385 0.665 4.52 1.25 ;
      RECT  3.86 1.25 4.52 1.37 ;
      RECT  3.86 1.37 3.975 1.45 ;
      RECT  1.335 0.55 2.045 0.67 ;
      RECT  1.955 0.67 2.045 1.23 ;
      RECT  1.19 1.23 2.045 1.26 ;
      RECT  1.19 1.26 3.39 1.35 ;
      RECT  3.3 1.35 3.39 1.45 ;
      RECT  3.3 1.45 3.975 1.54 ;
      RECT  4.87 1.425 5.655 1.525 ;
      LAYER M2 ;
      RECT  0.535 0.35 6.26 0.45 ;
      RECT  1.045 0.55 6.03 0.65 ;
      RECT  0.71 0.95 4.18 1.05 ;
      RECT  4.6 1.35 7.675 1.45 ;
      LAYER V1 ;
      RECT  0.575 0.35 0.675 0.45 ;
      RECT  1.35 0.35 1.45 0.45 ;
      RECT  6.12 0.35 6.22 0.45 ;
      RECT  1.085 0.55 1.185 0.65 ;
      RECT  5.89 0.55 5.99 0.65 ;
      RECT  0.75 0.95 0.85 1.05 ;
      RECT  3.45 0.95 3.55 1.05 ;
      RECT  4.03 0.95 4.13 1.05 ;
      RECT  4.64 1.35 4.74 1.45 ;
      RECT  7.535 1.35 7.635 1.45 ;
  END
END SEN_FDPRBSBQ_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPSBQ_D_1
#      Description : "D-Flip Flop pos-edge triggered, lo-async-set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,preset=!SD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPSBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FDPSBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.1 0.68 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.31 4.51 0.49 ;
      RECT  4.35 0.49 4.45 1.11 ;
      RECT  4.35 1.11 4.51 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.69 0.915 ;
      RECT  1.84 0.705 2.18 0.905 ;
      LAYER M2 ;
      RECT  1.8 0.75 3.725 0.85 ;
      LAYER V1 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  3.585 0.75 3.685 0.85 ;
      RECT  1.84 0.75 1.94 0.85 ;
      RECT  2.04 0.75 2.14 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.425 0.45 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.775 1.425 0.905 1.75 ;
      RECT  1.745 1.415 1.875 1.75 ;
      RECT  2.35 1.415 2.52 1.75 ;
      RECT  3.385 1.425 3.515 1.75 ;
      RECT  4.14 1.21 4.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.745 0.05 0.915 0.19 ;
      RECT  1.9 0.05 2.07 0.19 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  3.645 0.05 3.775 0.39 ;
      RECT  4.14 0.05 4.26 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.26 0.16 3.16 0.25 ;
      RECT  2.26 0.25 2.35 0.28 ;
      RECT  2.66 0.25 2.75 0.745 ;
      RECT  3.07 0.25 3.16 0.96 ;
      RECT  1.16 0.15 1.76 0.26 ;
      RECT  1.67 0.26 1.76 0.28 ;
      RECT  1.16 0.26 1.25 0.3 ;
      RECT  1.67 0.28 2.35 0.37 ;
      RECT  0.585 0.3 1.25 0.39 ;
      RECT  0.585 0.39 0.705 0.63 ;
      RECT  1.16 0.39 1.25 1.015 ;
      RECT  0.56 1.015 1.25 1.135 ;
      RECT  1.365 0.355 1.485 0.46 ;
      RECT  1.365 0.46 2.37 0.55 ;
      RECT  2.275 0.55 2.37 0.715 ;
      RECT  1.365 0.55 1.47 1.255 ;
      RECT  2.275 0.715 2.38 0.905 ;
      RECT  1.21 1.255 1.47 1.375 ;
      RECT  3.29 0.41 3.4 0.52 ;
      RECT  3.29 0.52 4.03 0.61 ;
      RECT  3.91 0.225 4.03 0.52 ;
      RECT  3.91 0.61 4.03 0.785 ;
      RECT  3.91 0.785 4.25 0.895 ;
      RECT  3.96 0.895 4.05 1.255 ;
      RECT  3.88 1.255 4.05 1.45 ;
      RECT  2.46 0.39 2.56 0.585 ;
      RECT  2.47 0.585 2.56 1.03 ;
      RECT  1.59 0.73 1.7 1.03 ;
      RECT  1.59 1.03 2.75 1.145 ;
      RECT  2.86 0.365 2.965 1.065 ;
      RECT  2.86 1.065 3.87 1.155 ;
      RECT  3.76 0.98 3.87 1.065 ;
      RECT  2.86 1.155 2.965 1.31 ;
      RECT  1.56 1.235 2.77 1.325 ;
      RECT  1.56 1.325 1.65 1.52 ;
      RECT  2.66 1.325 2.77 1.65 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 0.45 0.59 ;
      RECT  0.36 0.59 0.45 0.755 ;
      RECT  0.36 0.755 0.53 0.925 ;
      RECT  0.36 0.925 0.45 1.225 ;
      RECT  0.065 1.225 1.11 1.315 ;
      RECT  0.065 1.315 0.185 1.455 ;
      RECT  1.02 1.315 1.11 1.52 ;
      RECT  1.02 1.52 1.65 1.64 ;
      RECT  3.13 1.245 3.77 1.335 ;
      RECT  3.13 1.335 3.25 1.62 ;
      RECT  3.65 1.335 3.77 1.62 ;
  END
END SEN_FDPSBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPSBQ_D_2
#      Description : "D-Flip Flop pos-edge triggered, lo-async-set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,preset=!SD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPSBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FDPSBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.1 0.68 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.31 4.65 0.49 ;
      RECT  4.55 0.49 4.65 1.11 ;
      RECT  4.35 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.67 0.915 ;
      RECT  1.84 0.705 2.18 0.905 ;
      LAYER M2 ;
      RECT  1.8 0.75 3.69 0.85 ;
      LAYER V1 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  1.84 0.75 1.94 0.85 ;
      RECT  2.04 0.75 2.14 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.425 0.45 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.775 1.425 0.905 1.75 ;
      RECT  1.745 1.415 1.875 1.75 ;
      RECT  2.35 1.415 2.52 1.75 ;
      RECT  3.385 1.425 3.515 1.75 ;
      RECT  4.14 1.21 4.26 1.75 ;
      RECT  4.74 1.21 4.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.745 0.05 0.915 0.19 ;
      RECT  1.9 0.05 2.07 0.19 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  3.645 0.05 3.775 0.39 ;
      RECT  4.14 0.05 4.26 0.59 ;
      RECT  4.74 0.05 4.86 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.26 0.16 3.16 0.25 ;
      RECT  2.26 0.25 2.35 0.28 ;
      RECT  2.66 0.25 2.75 0.745 ;
      RECT  3.07 0.25 3.16 0.96 ;
      RECT  1.16 0.15 1.76 0.26 ;
      RECT  1.67 0.26 1.76 0.28 ;
      RECT  1.16 0.26 1.25 0.3 ;
      RECT  1.67 0.28 2.35 0.37 ;
      RECT  0.585 0.3 1.25 0.39 ;
      RECT  0.585 0.39 0.705 0.63 ;
      RECT  1.16 0.39 1.25 1.015 ;
      RECT  0.56 1.015 1.25 1.135 ;
      RECT  1.365 0.355 1.485 0.46 ;
      RECT  1.365 0.46 2.37 0.55 ;
      RECT  2.275 0.55 2.37 0.715 ;
      RECT  1.365 0.55 1.47 1.255 ;
      RECT  2.275 0.715 2.38 0.905 ;
      RECT  1.21 1.255 1.47 1.375 ;
      RECT  3.29 0.41 3.4 0.52 ;
      RECT  3.29 0.52 4.05 0.61 ;
      RECT  3.91 0.225 4.05 0.52 ;
      RECT  3.96 0.61 4.05 0.785 ;
      RECT  3.96 0.785 4.46 0.895 ;
      RECT  3.96 0.895 4.05 1.255 ;
      RECT  3.88 1.255 4.05 1.45 ;
      RECT  2.46 0.39 2.56 0.585 ;
      RECT  2.47 0.585 2.56 1.03 ;
      RECT  1.59 0.715 1.7 1.03 ;
      RECT  1.59 1.03 2.75 1.145 ;
      RECT  2.86 0.365 2.965 1.065 ;
      RECT  2.86 1.065 3.87 1.155 ;
      RECT  3.76 0.88 3.87 1.065 ;
      RECT  2.86 1.155 2.965 1.31 ;
      RECT  1.56 1.235 2.77 1.325 ;
      RECT  1.56 1.325 1.65 1.52 ;
      RECT  2.66 1.325 2.77 1.65 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 0.45 0.59 ;
      RECT  0.36 0.59 0.45 0.755 ;
      RECT  0.36 0.755 0.53 0.925 ;
      RECT  0.36 0.925 0.45 1.225 ;
      RECT  0.065 1.225 1.11 1.315 ;
      RECT  0.065 1.315 0.185 1.455 ;
      RECT  1.02 1.315 1.11 1.52 ;
      RECT  1.02 1.52 1.65 1.64 ;
      RECT  3.13 1.245 3.77 1.335 ;
      RECT  3.13 1.335 3.25 1.62 ;
      RECT  3.65 1.335 3.77 1.62 ;
  END
END SEN_FDPSBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FDPSBQ_D_4
#      Description : "D-Flip Flop pos-edge triggered, lo-async-set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=D,preset=!SD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FDPSBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FDPSBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.1 0.68 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 5.05 0.69 ;
      RECT  4.95 0.69 5.05 1.11 ;
      RECT  4.35 1.11 5.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.345 0.71 3.67 0.915 ;
      RECT  1.84 0.705 2.18 0.905 ;
      LAYER M2 ;
      RECT  1.8 0.75 3.69 0.85 ;
      LAYER V1 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  1.84 0.75 1.94 0.85 ;
      RECT  2.04 0.75 2.14 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END SD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.425 0.45 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  0.775 1.41 0.905 1.75 ;
      RECT  1.745 1.415 1.875 1.75 ;
      RECT  2.35 1.415 2.52 1.75 ;
      RECT  3.385 1.425 3.515 1.75 ;
      RECT  4.14 1.21 4.26 1.75 ;
      RECT  4.655 1.41 4.785 1.75 ;
      RECT  5.18 1.21 5.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  0.745 0.05 0.915 0.19 ;
      RECT  1.9 0.05 2.07 0.19 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  3.645 0.05 3.775 0.39 ;
      RECT  4.655 0.05 4.785 0.39 ;
      RECT  4.14 0.05 4.26 0.59 ;
      RECT  5.18 0.05 5.3 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.26 0.16 3.16 0.25 ;
      RECT  2.26 0.25 2.35 0.28 ;
      RECT  2.66 0.25 2.75 0.745 ;
      RECT  3.07 0.25 3.16 0.96 ;
      RECT  1.16 0.15 1.76 0.26 ;
      RECT  1.67 0.26 1.76 0.28 ;
      RECT  1.16 0.26 1.25 0.3 ;
      RECT  1.67 0.28 2.35 0.37 ;
      RECT  0.585 0.3 1.25 0.39 ;
      RECT  0.585 0.39 0.705 0.63 ;
      RECT  1.16 0.39 1.25 1.015 ;
      RECT  0.56 1.015 1.25 1.135 ;
      RECT  1.365 0.355 1.485 0.46 ;
      RECT  1.365 0.46 2.37 0.55 ;
      RECT  2.275 0.55 2.37 0.715 ;
      RECT  1.365 0.55 1.47 1.255 ;
      RECT  2.275 0.715 2.38 0.905 ;
      RECT  1.21 1.255 1.47 1.375 ;
      RECT  3.29 0.41 3.4 0.52 ;
      RECT  3.29 0.52 4.05 0.61 ;
      RECT  3.91 0.2 4.05 0.52 ;
      RECT  3.96 0.61 4.05 0.785 ;
      RECT  3.96 0.785 4.86 0.895 ;
      RECT  3.96 0.895 4.05 1.255 ;
      RECT  3.88 1.255 4.05 1.45 ;
      RECT  2.46 0.39 2.56 0.585 ;
      RECT  2.47 0.585 2.56 1.03 ;
      RECT  1.59 0.73 1.7 1.03 ;
      RECT  1.59 1.03 2.75 1.145 ;
      RECT  2.86 0.365 2.965 1.065 ;
      RECT  2.86 1.065 3.87 1.155 ;
      RECT  3.76 0.735 3.87 1.065 ;
      RECT  2.86 1.155 2.965 1.31 ;
      RECT  1.56 1.235 2.77 1.325 ;
      RECT  1.56 1.325 1.65 1.52 ;
      RECT  2.66 1.325 2.77 1.65 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 0.45 0.59 ;
      RECT  0.36 0.59 0.45 0.755 ;
      RECT  0.36 0.755 0.53 0.925 ;
      RECT  0.36 0.925 0.45 1.225 ;
      RECT  0.065 1.225 1.11 1.315 ;
      RECT  0.065 1.315 0.185 1.455 ;
      RECT  1.02 1.315 1.11 1.52 ;
      RECT  1.02 1.52 1.65 1.64 ;
      RECT  3.13 1.245 3.77 1.335 ;
      RECT  3.13 1.335 3.25 1.62 ;
      RECT  3.65 1.335 3.77 1.62 ;
  END
END SEN_FDPSBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FILL1
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FILL1
  CLASS CORE SPACER ;
  FOREIGN SEN_FILL1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.2 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.2 0.05 ;
    END
  END VSS
END SEN_FILL1
#-----------------------------------------------------------------------
#      Cell        : SEN_FILL16
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FILL16
  CLASS CORE SPACER ;
  FOREIGN SEN_FILL16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
END SEN_FILL16
#-----------------------------------------------------------------------
#      Cell        : SEN_FILL2
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FILL2
  CLASS CORE SPACER ;
  FOREIGN SEN_FILL2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.4 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.4 0.05 ;
    END
  END VSS
END SEN_FILL2
#-----------------------------------------------------------------------
#      Cell        : SEN_FILL32
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FILL32
  CLASS CORE SPACER ;
  FOREIGN SEN_FILL32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
END SEN_FILL32
#-----------------------------------------------------------------------
#      Cell        : SEN_FILL4
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FILL4
  CLASS CORE SPACER ;
  FOREIGN SEN_FILL4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
    END
  END VSS
END SEN_FILL4
#-----------------------------------------------------------------------
#      Cell        : SEN_FILL64
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FILL64
  CLASS CORE SPACER ;
  FOREIGN SEN_FILL64 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
END SEN_FILL64
#-----------------------------------------------------------------------
#      Cell        : SEN_FILL8
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FILL8
  CLASS CORE SPACER ;
  FOREIGN SEN_FILL8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
END SEN_FILL8
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPNW1
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPNW1
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPNW1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
END SEN_CAPNW1
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPNW16
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPNW16
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPNW16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
END SEN_CAPNW16
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPNW2
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPNW2
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPNW2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
END SEN_CAPNW2
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPNW32
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPNW32
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPNW32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
END SEN_CAPNW32
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPNW4
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPNW4
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPNW4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
END SEN_CAPNW4
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPNW64
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPNW64
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPNW64 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
END SEN_CAPNW64
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPNW8
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPNW8
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPNW8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
END SEN_CAPNW8
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPCRNI10
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPCRNI10
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPCRNI10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
END SEN_CAPCRNI10
#-----------------------------------------------------------------------
#      Cell        : SEN_CAPLR10
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_CAPLR10
  CLASS CORE SPACER ;
  FOREIGN SEN_CAPLR10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.305 0.05 0.405 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.305 -0.05 0.405 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.255 0.665 1.865 0.755 ;
  END
END SEN_CAPLR10
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD1
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD1
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 0.2 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 0.2 0.05 ;
    END
  END VSS
END SEN_RAIL2TD1
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD128
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD128
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD128 0 0 ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 25.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 25.6 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 25.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 25.6 0.05 ;
    END
  END VSS
END SEN_RAIL2TD128
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD16
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD16
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 3.2 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 3.2 0.05 ;
    END
  END VSS
END SEN_RAIL2TD16
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD2
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD2
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 0.4 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 0.4 0.05 ;
    END
  END VSS
END SEN_RAIL2TD2
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD256
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD256
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD256 0 0 ;
  ORIGIN 0 0 ;
  SIZE 51.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 51.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 51.2 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 51.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 51.2 0.05 ;
    END
  END VSS
END SEN_RAIL2TD256
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD32
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD32
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 6.4 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 6.4 0.05 ;
    END
  END VSS
END SEN_RAIL2TD32
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD4
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD4
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 0.8 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 0.8 0.05 ;
    END
  END VSS
END SEN_RAIL2TD4
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD64
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD64
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD64 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 12.8 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 12.8 0.05 ;
    END
  END VSS
END SEN_RAIL2TD64
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TD8
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TD8
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TD8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.65 1.6 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.15 1.6 0.05 ;
    END
  END VSS
END SEN_RAIL2TD8
#-----------------------------------------------------------------------
#      Cell        : SEN_FILL_ECO1
#      Description : "Filler cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FILL_ECO1
  CLASS CORE SPACER ;
  FOREIGN SEN_FILL_ECO1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
END SEN_FILL_ECO1
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T1
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T1
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.2 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.2 0.05 ;
    END
  END VSS
END SEN_RAIL1T1
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T128
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T128
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T128 0 0 ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 25.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 25.6 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 25.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 25.6 0.05 ;
    END
  END VSS
END SEN_RAIL1T128
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T16
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T16
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
    END
  END VSS
END SEN_RAIL1T16
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T2
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T2
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.4 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.4 0.05 ;
    END
  END VSS
END SEN_RAIL1T2
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T256
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T256
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T256 0 0 ;
  ORIGIN 0 0 ;
  SIZE 51.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 51.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 51.2 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 51.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 51.2 0.05 ;
    END
  END VSS
END SEN_RAIL1T256
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T32
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T32
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
    END
  END VSS
END SEN_RAIL1T32
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T4
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T4
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
    END
  END VSS
END SEN_RAIL1T4
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T64
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T64
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T64 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
    END
  END VSS
END SEN_RAIL1T64
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL1T8
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL1T8
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL1T8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
    END
  END VSS
END SEN_RAIL1T8
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T1
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T1
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 0.2 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 0.2 0.2 ;
    END
  END VSS
END SEN_RAIL3T1
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T128
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T128
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T128 0 0 ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 25.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 25.6 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 25.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 25.6 0.2 ;
    END
  END VSS
END SEN_RAIL3T128
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T16
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T16
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 3.2 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 3.2 0.2 ;
    END
  END VSS
END SEN_RAIL3T16
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T2
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T2
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 0.4 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 0.4 0.2 ;
    END
  END VSS
END SEN_RAIL3T2
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T256
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T256
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T256 0 0 ;
  ORIGIN 0 0 ;
  SIZE 51.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 51.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 51.2 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 51.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 51.2 0.2 ;
    END
  END VSS
END SEN_RAIL3T256
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T32
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T32
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 6.4 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 6.4 0.2 ;
    END
  END VSS
END SEN_RAIL3T32
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T4
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T4
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 0.8 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 0.8 0.2 ;
    END
  END VSS
END SEN_RAIL3T4
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T64
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T64
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T64 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 12.8 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 12.8 0.2 ;
    END
  END VSS
END SEN_RAIL3T64
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL3T8
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL3T8
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL3T8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.6 1.6 2.0 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.2 1.6 0.2 ;
    END
  END VSS
END SEN_RAIL3T8
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU1
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU1
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.2 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.2 0.15 ;
    END
  END VSS
END SEN_RAIL2TU1
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU128
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU128
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU128 0 0 ;
  ORIGIN 0 0 ;
  SIZE 25.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 25.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 25.6 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 25.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 25.6 0.15 ;
    END
  END VSS
END SEN_RAIL2TU128
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU16
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU16
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.15 ;
    END
  END VSS
END SEN_RAIL2TU16
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU2
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU2
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.4 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.4 0.15 ;
    END
  END VSS
END SEN_RAIL2TU2
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU256
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU256
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU256 0 0 ;
  ORIGIN 0 0 ;
  SIZE 51.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 51.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 51.2 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 51.2 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 51.2 0.15 ;
    END
  END VSS
END SEN_RAIL2TU256
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU32
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU32
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.15 ;
    END
  END VSS
END SEN_RAIL2TU32
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU4
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU4
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.15 ;
    END
  END VSS
END SEN_RAIL2TU4
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU64
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU64
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU64 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.15 ;
    END
  END VSS
END SEN_RAIL2TU64
#-----------------------------------------------------------------------
#      Cell        : SEN_RAIL2TU8
#      Description : "Rail cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_RAIL2TU8
  CLASS CORE SPACER ;
  FOREIGN SEN_RAIL2TU8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.95 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.15 ;
    END
  END VSS
END SEN_RAIL2TU8
#-----------------------------------------------------------------------
#      Cell        : SEN_TAP_DS
#      Description : "Tap cell"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_TAP_DS
  CLASS CORE WELLTAP ;
  FOREIGN SEN_TAP_DS 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.15 1.25 0.25 1.75 ;
      RECT  0.0 1.75 0.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.4 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.4 0.05 ;
      RECT  0.15 0.05 0.25 0.55 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.4 0.05 ;
    END
  END VSS
END SEN_TAP_DS
#-----------------------------------------------------------------------
#      Cell        : SEN_DCAP16
#      Description : "Filler cell with De-coupling"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DCAP16
  CLASS CORE SPACER ;
  FOREIGN SEN_DCAP16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 0.41 2.825 0.59 ;
      RECT  0.055 0.59 0.175 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  2.965 0.05 3.085 1.075 ;
      RECT  0.315 1.075 3.085 1.255 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
END SEN_DCAP16
#-----------------------------------------------------------------------
#      Cell        : SEN_DCAP32
#      Description : "Filler cell with De-coupling"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DCAP32
  CLASS CORE SPACER ;
  FOREIGN SEN_DCAP32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 0.41 5.945 0.59 ;
      RECT  0.055 0.59 0.175 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  6.085 0.05 6.205 1.075 ;
      RECT  0.315 1.075 6.205 1.255 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
END SEN_DCAP32
#-----------------------------------------------------------------------
#      Cell        : SEN_DCAP4
#      Description : "Filler cell with De-coupling"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DCAP4
  CLASS CORE SPACER ;
  FOREIGN SEN_DCAP4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 0.41 0.535 0.59 ;
      RECT  0.055 0.59 0.175 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.625 0.05 0.745 1.01 ;
      RECT  0.265 1.01 0.745 1.19 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
END SEN_DCAP4
#-----------------------------------------------------------------------
#      Cell        : SEN_DCAP64
#      Description : "Filler cell with De-coupling"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DCAP64
  CLASS CORE SPACER ;
  FOREIGN SEN_DCAP64 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 0.41 12.445 0.59 ;
      RECT  0.055 0.59 0.175 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  12.585 0.05 12.705 1.075 ;
      RECT  0.315 1.075 12.705 1.255 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
END SEN_DCAP64
#-----------------------------------------------------------------------
#      Cell        : SEN_DCAP8
#      Description : "Filler cell with De-coupling"
#      Equation    : None
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_DCAP8
  CLASS CORE SPACER ;
  FOREIGN SEN_DCAP8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 0.41 1.265 0.59 ;
      RECT  0.055 0.59 0.175 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  1.405 0.05 1.525 1.075 ;
      RECT  0.315 1.075 1.525 1.255 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
END SEN_DCAP8
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDAO22PQ_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&((A1&A2)|(B1&B2)))|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDAO22PQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDAO22PQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.695 ;
      RECT  0.55 0.695 0.85 0.785 ;
      RECT  0.7 0.785 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.885 ;
      RECT  0.35 0.885 0.585 0.985 ;
      RECT  0.35 0.985 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B2
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.215 0.825 5.38 1.035 ;
      RECT  5.28 1.035 5.38 1.29 ;
      RECT  3.12 0.625 3.22 1.315 ;
      LAYER M2 ;
      RECT  3.08 1.15 5.42 1.25 ;
      LAYER V1 ;
      RECT  5.28 1.15 5.38 1.25 ;
      RECT  3.12 1.15 3.22 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1239 ;
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.31 6.45 1.29 ;
    END
    ANTENNADIFFAREA 0.178 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.55 0.91 2.25 1.09 ;
      RECT  2.15 0.71 2.25 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.4 0.445 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.595 1.39 1.715 1.75 ;
      RECT  2.6 1.425 2.73 1.75 ;
      RECT  4.035 1.425 4.155 1.75 ;
      RECT  5.28 1.385 5.45 1.75 ;
      RECT  6.08 1.405 6.2 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  5.315 0.05 5.435 0.26 ;
      RECT  1.565 0.05 1.685 0.385 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  2.515 0.05 2.635 0.41 ;
      RECT  4.035 0.05 4.155 0.41 ;
      RECT  1.085 0.05 1.195 0.415 ;
      RECT  6.08 0.05 6.2 0.605 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.025 0.14 3.895 0.23 ;
      RECT  3.775 0.23 3.895 0.405 ;
      RECT  3.025 0.23 3.145 0.415 ;
      RECT  4.555 0.15 5.125 0.24 ;
      RECT  5.035 0.24 5.125 0.35 ;
      RECT  4.555 0.24 4.675 1.41 ;
      RECT  5.035 0.35 5.625 0.44 ;
      RECT  5.525 0.14 5.625 0.35 ;
      RECT  0.535 0.21 0.95 0.335 ;
      RECT  0.85 0.335 0.95 0.495 ;
      RECT  0.85 0.495 1.04 0.585 ;
      RECT  0.94 0.585 1.04 1.24 ;
      RECT  0.81 1.24 1.04 1.36 ;
      RECT  2.005 0.235 2.285 0.355 ;
      RECT  2.185 0.355 2.285 0.58 ;
      RECT  1.775 0.245 1.875 0.445 ;
      RECT  1.775 0.445 2.01 0.535 ;
      RECT  1.91 0.535 2.01 0.79 ;
      RECT  3.495 0.35 3.68 0.45 ;
      RECT  3.55 0.45 3.68 0.695 ;
      RECT  3.265 0.32 3.405 0.49 ;
      RECT  3.31 0.49 3.405 0.825 ;
      RECT  3.31 0.825 4.22 0.915 ;
      RECT  4.12 0.715 4.22 0.825 ;
      RECT  3.31 0.915 3.4 1.415 ;
      RECT  3.285 1.415 3.4 1.465 ;
      RECT  3.285 1.465 3.72 1.585 ;
      RECT  2.795 0.165 2.915 0.505 ;
      RECT  2.385 0.505 3.03 0.605 ;
      RECT  2.94 0.605 3.03 1.025 ;
      RECT  2.75 1.025 3.03 1.15 ;
      RECT  4.295 0.37 4.44 0.505 ;
      RECT  3.8 0.505 4.44 0.605 ;
      RECT  4.35 0.605 4.44 1.04 ;
      RECT  4.245 1.04 4.44 1.145 ;
      RECT  1.34 0.17 1.455 0.52 ;
      RECT  1.34 0.52 1.555 0.62 ;
      RECT  1.34 0.62 1.43 1.18 ;
      RECT  1.34 1.18 2.33 1.28 ;
      RECT  1.34 1.28 1.45 1.605 ;
      RECT  5.02 0.545 5.215 0.665 ;
      RECT  5.02 0.665 5.125 1.35 ;
      RECT  5.02 1.35 5.19 1.47 ;
      RECT  5.02 1.47 5.11 1.56 ;
      RECT  3.57 1.005 3.8 1.115 ;
      RECT  3.71 1.115 3.8 1.235 ;
      RECT  3.71 1.235 4.37 1.335 ;
      RECT  4.28 1.335 4.37 1.56 ;
      RECT  4.28 1.56 5.11 1.66 ;
      RECT  5.535 0.55 5.73 0.665 ;
      RECT  5.585 0.665 5.73 0.96 ;
      RECT  5.585 0.96 5.945 1.06 ;
      RECT  5.585 1.06 5.705 1.49 ;
      RECT  5.82 0.38 5.94 0.7 ;
      RECT  5.82 0.7 6.15 0.79 ;
      RECT  6.05 0.79 6.15 1.22 ;
      RECT  5.82 1.22 6.15 1.31 ;
      RECT  5.82 1.31 5.94 1.625 ;
      RECT  0.07 1.215 0.705 1.305 ;
      RECT  0.07 1.305 0.185 1.44 ;
      RECT  0.585 1.305 0.705 1.515 ;
      RECT  0.585 1.515 1.225 1.605 ;
      RECT  1.11 1.42 1.225 1.515 ;
      RECT  2.42 1.245 3.03 1.335 ;
      RECT  2.94 1.335 3.03 1.44 ;
      RECT  2.42 1.335 2.51 1.48 ;
      RECT  2.94 1.44 3.19 1.56 ;
      RECT  2.005 1.48 2.51 1.595 ;
      RECT  4.82 0.39 4.93 1.415 ;
      LAYER M2 ;
      RECT  0.81 0.35 1.915 0.45 ;
      RECT  2.145 0.35 3.675 0.45 ;
      RECT  4.79 0.95 6.19 1.05 ;
      LAYER V1 ;
      RECT  0.85 0.35 0.95 0.45 ;
      RECT  1.775 0.35 1.875 0.45 ;
      RECT  2.185 0.35 2.285 0.45 ;
      RECT  3.535 0.35 3.635 0.45 ;
      RECT  4.83 0.95 4.93 1.05 ;
      RECT  6.05 0.95 6.15 1.05 ;
  END
END SEN_FSDAO22PQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDAO22PQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&((A1&A2)|(B1&B2)))|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDAO22PQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDAO22PQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.665 ;
      RECT  0.55 0.665 0.85 0.755 ;
      RECT  0.705 0.755 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.845 ;
      RECT  0.35 0.845 0.525 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B2
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.215 0.865 5.38 1.04 ;
      RECT  5.28 1.04 5.38 1.29 ;
      RECT  3.12 0.625 3.22 1.315 ;
      LAYER M2 ;
      RECT  3.08 1.15 5.42 1.25 ;
      LAYER V1 ;
      RECT  5.28 1.15 5.38 1.25 ;
      RECT  3.12 1.15 3.22 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1239 ;
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.31 6.45 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.55 0.91 2.25 1.09 ;
      RECT  2.15 0.62 2.25 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.4 0.445 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.595 1.39 1.715 1.75 ;
      RECT  2.6 1.425 2.72 1.75 ;
      RECT  4.035 1.425 4.155 1.75 ;
      RECT  5.28 1.385 5.45 1.75 ;
      RECT  6.08 1.4 6.2 1.75 ;
      RECT  6.6 1.21 6.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  5.315 0.05 5.435 0.26 ;
      RECT  1.075 0.05 1.195 0.385 ;
      RECT  1.565 0.05 1.685 0.385 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  4.035 0.05 4.155 0.41 ;
      RECT  2.515 0.05 2.635 0.415 ;
      RECT  6.6 0.05 6.72 0.59 ;
      RECT  6.08 0.05 6.2 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.025 0.14 3.895 0.23 ;
      RECT  3.025 0.23 3.145 0.415 ;
      RECT  3.78 0.23 3.895 0.42 ;
      RECT  4.555 0.195 5.125 0.285 ;
      RECT  5.035 0.285 5.125 0.35 ;
      RECT  4.555 0.285 4.675 1.435 ;
      RECT  5.035 0.35 5.625 0.44 ;
      RECT  5.525 0.14 5.625 0.35 ;
      RECT  0.54 0.215 0.95 0.335 ;
      RECT  0.85 0.335 0.95 0.48 ;
      RECT  0.85 0.48 1.04 0.57 ;
      RECT  0.94 0.57 1.04 1.24 ;
      RECT  0.8 1.24 1.04 1.36 ;
      RECT  2.01 0.23 2.28 0.355 ;
      RECT  2.18 0.355 2.28 0.53 ;
      RECT  1.775 0.245 1.875 0.445 ;
      RECT  1.775 0.445 2.01 0.535 ;
      RECT  1.91 0.535 2.01 0.775 ;
      RECT  3.495 0.35 3.68 0.45 ;
      RECT  3.55 0.45 3.68 0.695 ;
      RECT  3.285 0.32 3.405 0.49 ;
      RECT  3.31 0.49 3.405 0.785 ;
      RECT  3.31 0.785 4.255 0.875 ;
      RECT  3.31 0.875 3.4 1.415 ;
      RECT  3.275 1.415 3.4 1.465 ;
      RECT  3.275 1.465 3.72 1.585 ;
      RECT  2.795 0.17 2.915 0.505 ;
      RECT  2.37 0.505 3.03 0.605 ;
      RECT  2.94 0.605 3.03 1.025 ;
      RECT  2.37 0.605 2.46 1.045 ;
      RECT  2.745 1.025 3.03 1.15 ;
      RECT  4.295 0.33 4.44 0.505 ;
      RECT  3.97 0.505 4.44 0.59 ;
      RECT  3.795 0.59 4.44 0.605 ;
      RECT  3.795 0.605 4.075 0.695 ;
      RECT  4.35 0.605 4.44 1.015 ;
      RECT  4.245 1.015 4.44 1.135 ;
      RECT  1.34 0.165 1.455 0.52 ;
      RECT  1.34 0.52 1.585 0.62 ;
      RECT  1.34 0.62 1.43 1.18 ;
      RECT  1.34 1.18 2.33 1.28 ;
      RECT  1.34 1.28 1.45 1.605 ;
      RECT  5.02 0.545 5.22 0.665 ;
      RECT  5.02 0.665 5.125 1.35 ;
      RECT  5.02 1.35 5.19 1.47 ;
      RECT  5.02 1.47 5.11 1.56 ;
      RECT  3.57 0.975 3.8 1.07 ;
      RECT  3.7 1.07 3.8 1.235 ;
      RECT  3.7 1.235 4.37 1.335 ;
      RECT  4.28 1.335 4.37 1.56 ;
      RECT  4.28 1.56 5.11 1.66 ;
      RECT  5.535 0.54 5.73 0.665 ;
      RECT  5.585 0.665 5.73 0.96 ;
      RECT  5.585 0.96 5.94 1.06 ;
      RECT  5.585 1.06 5.705 1.505 ;
      RECT  5.82 0.39 5.94 0.7 ;
      RECT  5.82 0.7 6.15 0.79 ;
      RECT  6.05 0.79 6.15 1.22 ;
      RECT  5.82 1.22 6.15 1.31 ;
      RECT  5.82 1.31 5.94 1.63 ;
      RECT  0.065 1.215 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.445 ;
      RECT  0.585 1.305 0.705 1.515 ;
      RECT  0.585 1.515 1.225 1.605 ;
      RECT  1.105 1.425 1.225 1.515 ;
      RECT  2.42 1.245 3.03 1.335 ;
      RECT  2.94 1.335 3.03 1.44 ;
      RECT  2.42 1.335 2.51 1.48 ;
      RECT  2.94 1.44 3.175 1.56 ;
      RECT  2.005 1.48 2.51 1.595 ;
      RECT  4.82 0.385 4.93 1.435 ;
      LAYER M2 ;
      RECT  0.81 0.35 1.915 0.45 ;
      RECT  2.14 0.35 3.675 0.45 ;
      RECT  4.79 0.95 6.19 1.05 ;
      LAYER V1 ;
      RECT  0.85 0.35 0.95 0.45 ;
      RECT  1.775 0.35 1.875 0.45 ;
      RECT  2.18 0.35 2.28 0.45 ;
      RECT  3.535 0.35 3.635 0.45 ;
      RECT  4.83 0.95 4.93 1.05 ;
      RECT  6.05 0.95 6.15 1.05 ;
  END
END SEN_FSDAO22PQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDAO22PQ_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&((A1&A2)|(B1&B2)))|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDAO22PQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDAO22PQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.71 ;
      RECT  0.55 0.71 0.85 0.9 ;
      RECT  0.705 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.0 ;
      RECT  0.35 1.0 0.575 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END B2
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.215 0.9 5.38 1.11 ;
      RECT  5.28 1.11 5.38 1.29 ;
      RECT  3.12 0.625 3.22 1.315 ;
      LAYER M2 ;
      RECT  3.08 1.15 5.42 1.25 ;
      LAYER V1 ;
      RECT  5.28 1.15 5.38 1.25 ;
      RECT  3.12 1.15 3.22 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1239 ;
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.575 6.565 0.665 ;
      RECT  6.35 0.665 6.45 1.11 ;
      RECT  6.35 1.11 7.05 1.29 ;
      RECT  6.95 0.45 7.05 1.11 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.55 0.91 2.25 1.09 ;
      RECT  2.15 0.61 2.25 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.395 0.445 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  1.595 1.39 1.715 1.75 ;
      RECT  2.6 1.43 2.73 1.75 ;
      RECT  4.035 1.44 4.155 1.75 ;
      RECT  5.28 1.38 5.45 1.75 ;
      RECT  6.16 1.4 6.28 1.75 ;
      RECT  6.68 1.38 6.8 1.75 ;
      RECT  7.2 1.21 7.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  5.315 0.05 5.435 0.26 ;
      RECT  6.135 0.05 6.305 0.305 ;
      RECT  6.655 0.05 6.825 0.305 ;
      RECT  1.565 0.05 1.685 0.385 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  1.075 0.05 1.195 0.405 ;
      RECT  2.515 0.05 2.635 0.41 ;
      RECT  4.035 0.05 4.155 0.415 ;
      RECT  7.2 0.05 7.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.025 0.14 3.895 0.23 ;
      RECT  3.775 0.23 3.895 0.405 ;
      RECT  3.025 0.23 3.145 0.415 ;
      RECT  4.555 0.15 5.125 0.24 ;
      RECT  5.035 0.24 5.125 0.35 ;
      RECT  4.555 0.24 4.675 1.405 ;
      RECT  5.035 0.35 5.92 0.395 ;
      RECT  5.525 0.14 5.625 0.35 ;
      RECT  5.035 0.395 6.745 0.44 ;
      RECT  5.83 0.44 6.745 0.485 ;
      RECT  6.655 0.485 6.745 0.755 ;
      RECT  6.545 0.755 6.855 0.925 ;
      RECT  0.53 0.215 0.95 0.335 ;
      RECT  0.85 0.335 0.95 0.495 ;
      RECT  0.85 0.495 1.04 0.585 ;
      RECT  0.94 0.585 1.04 1.24 ;
      RECT  0.805 1.24 1.04 1.36 ;
      RECT  2.0 0.235 2.28 0.355 ;
      RECT  2.18 0.355 2.28 0.52 ;
      RECT  1.775 0.245 1.875 0.445 ;
      RECT  1.775 0.445 2.01 0.535 ;
      RECT  1.91 0.535 2.01 0.785 ;
      RECT  3.495 0.35 3.68 0.45 ;
      RECT  3.55 0.45 3.68 0.695 ;
      RECT  3.27 0.32 3.405 0.49 ;
      RECT  3.31 0.49 3.405 0.795 ;
      RECT  3.31 0.795 4.26 0.885 ;
      RECT  3.31 0.885 3.4 1.415 ;
      RECT  3.285 1.415 3.4 1.465 ;
      RECT  3.285 1.465 3.71 1.585 ;
      RECT  2.795 0.165 2.915 0.505 ;
      RECT  2.37 0.505 3.03 0.605 ;
      RECT  2.94 0.605 3.03 1.025 ;
      RECT  2.37 0.605 2.46 1.07 ;
      RECT  2.77 1.025 3.03 1.15 ;
      RECT  4.295 0.32 4.44 0.505 ;
      RECT  3.8 0.505 4.44 0.605 ;
      RECT  4.35 0.605 4.44 1.015 ;
      RECT  4.25 1.015 4.44 1.135 ;
      RECT  1.34 0.18 1.455 0.52 ;
      RECT  1.34 0.52 1.585 0.62 ;
      RECT  1.34 0.62 1.43 1.18 ;
      RECT  1.34 1.18 2.33 1.28 ;
      RECT  1.34 1.28 1.45 1.61 ;
      RECT  5.02 0.545 5.22 0.665 ;
      RECT  5.02 0.665 5.125 1.35 ;
      RECT  5.02 1.35 5.19 1.47 ;
      RECT  5.02 1.47 5.11 1.56 ;
      RECT  3.63 0.975 3.74 1.235 ;
      RECT  3.63 1.235 4.37 1.335 ;
      RECT  4.28 1.335 4.37 1.56 ;
      RECT  4.28 1.56 5.11 1.66 ;
      RECT  5.53 0.55 5.73 0.665 ;
      RECT  5.585 0.665 5.73 0.96 ;
      RECT  5.585 0.96 6.005 1.06 ;
      RECT  5.585 1.06 5.705 1.49 ;
      RECT  5.83 0.575 6.035 0.68 ;
      RECT  5.935 0.68 6.035 0.74 ;
      RECT  5.935 0.74 6.205 0.83 ;
      RECT  6.105 0.83 6.205 1.22 ;
      RECT  5.875 1.22 6.205 1.31 ;
      RECT  5.875 1.31 5.995 1.635 ;
      RECT  0.065 1.215 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.435 ;
      RECT  0.585 1.305 0.705 1.515 ;
      RECT  0.585 1.515 1.225 1.605 ;
      RECT  1.105 1.425 1.225 1.515 ;
      RECT  2.42 1.245 3.03 1.335 ;
      RECT  2.94 1.335 3.03 1.44 ;
      RECT  2.42 1.335 2.51 1.48 ;
      RECT  2.94 1.44 3.175 1.56 ;
      RECT  2.0 1.48 2.51 1.595 ;
      RECT  4.82 0.415 4.93 1.405 ;
      LAYER M2 ;
      RECT  0.81 0.35 1.915 0.45 ;
      RECT  2.14 0.35 3.675 0.45 ;
      RECT  4.79 0.95 6.245 1.05 ;
      LAYER V1 ;
      RECT  0.85 0.35 0.95 0.45 ;
      RECT  1.775 0.35 1.875 0.45 ;
      RECT  2.18 0.35 2.28 0.45 ;
      RECT  3.535 0.35 3.635 0.45 ;
      RECT  4.83 0.95 4.93 1.05 ;
      RECT  6.105 0.95 6.205 1.05 ;
  END
END SEN_FSDAO22PQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDAO22PQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&((A1&A2)|(B1&B2)))|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDAO22PQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDAO22PQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.71 ;
      RECT  0.55 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.98 ;
      RECT  0.35 0.98 0.575 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 ;
  END B2
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.39 0.92 5.485 1.11 ;
      RECT  5.39 1.11 5.65 1.2 ;
      RECT  5.55 1.2 5.65 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0756 ;
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.31 7.465 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 0.91 ;
      RECT  1.55 0.91 1.85 0.985 ;
      RECT  1.55 0.985 2.465 1.09 ;
      RECT  2.35 0.87 2.465 0.985 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 2.965 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.785 0.575 7.05 0.68 ;
      RECT  6.95 0.68 7.05 1.2 ;
      RECT  6.81 1.2 7.05 1.29 ;
      RECT  6.81 1.29 6.93 1.62 ;
    END
    ANTENNADIFFAREA 0.105 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.4 0.445 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  1.595 1.38 1.715 1.75 ;
      RECT  2.775 1.425 2.905 1.75 ;
      RECT  4.21 1.425 4.33 1.75 ;
      RECT  5.465 1.58 5.635 1.75 ;
      RECT  6.28 1.295 6.4 1.75 ;
      RECT  7.085 1.375 7.205 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  5.49 0.05 5.61 0.24 ;
      RECT  6.28 0.05 6.4 0.24 ;
      RECT  7.07 0.05 7.24 0.305 ;
      RECT  1.075 0.05 1.195 0.385 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  2.69 0.05 2.81 0.41 ;
      RECT  4.21 0.05 4.33 0.43 ;
      RECT  1.75 0.05 1.87 0.625 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.2 0.14 4.07 0.23 ;
      RECT  3.2 0.23 3.32 0.415 ;
      RECT  3.95 0.23 4.07 0.43 ;
      RECT  4.73 0.15 5.37 0.24 ;
      RECT  5.28 0.24 5.37 0.33 ;
      RECT  4.73 0.24 4.85 1.405 ;
      RECT  5.28 0.33 6.885 0.395 ;
      RECT  6.085 0.14 6.185 0.33 ;
      RECT  5.28 0.395 7.26 0.42 ;
      RECT  6.795 0.42 7.26 0.485 ;
      RECT  7.165 0.485 7.26 0.95 ;
      RECT  0.54 0.215 0.95 0.335 ;
      RECT  0.85 0.335 0.95 0.495 ;
      RECT  0.85 0.495 1.035 0.585 ;
      RECT  0.945 0.585 1.035 1.24 ;
      RECT  0.805 1.24 1.035 1.36 ;
      RECT  2.175 0.235 2.46 0.355 ;
      RECT  2.36 0.355 2.46 0.69 ;
      RECT  2.36 0.69 2.66 0.78 ;
      RECT  2.57 0.78 2.66 1.245 ;
      RECT  2.57 1.245 3.205 1.335 ;
      RECT  3.115 1.335 3.205 1.44 ;
      RECT  2.57 1.335 2.66 1.48 ;
      RECT  3.115 1.44 3.37 1.56 ;
      RECT  2.165 1.48 2.66 1.595 ;
      RECT  1.34 0.175 1.64 0.36 ;
      RECT  1.34 0.36 1.43 1.18 ;
      RECT  1.34 1.18 2.47 1.28 ;
      RECT  2.37 1.28 2.47 1.35 ;
      RECT  1.34 1.28 1.45 1.6 ;
      RECT  1.98 0.245 2.08 0.445 ;
      RECT  1.98 0.445 2.18 0.535 ;
      RECT  2.08 0.535 2.18 0.79 ;
      RECT  2.08 0.79 2.25 0.885 ;
      RECT  3.67 0.35 3.855 0.45 ;
      RECT  3.725 0.45 3.855 0.695 ;
      RECT  4.95 0.35 5.19 0.45 ;
      RECT  4.95 0.45 5.095 0.545 ;
      RECT  4.95 0.545 5.05 1.24 ;
      RECT  4.95 1.24 5.105 1.41 ;
      RECT  3.46 0.32 3.58 0.49 ;
      RECT  3.485 0.49 3.58 0.785 ;
      RECT  3.485 0.785 4.43 0.875 ;
      RECT  3.485 0.875 3.575 1.365 ;
      RECT  3.46 1.365 3.575 1.465 ;
      RECT  3.46 1.465 3.895 1.585 ;
      RECT  2.97 0.19 3.09 0.505 ;
      RECT  2.56 0.505 3.145 0.6 ;
      RECT  3.055 0.6 3.145 1.025 ;
      RECT  2.945 1.025 3.145 1.15 ;
      RECT  4.47 0.305 4.615 0.595 ;
      RECT  3.97 0.595 4.615 0.695 ;
      RECT  4.525 0.695 4.615 1.025 ;
      RECT  4.42 1.025 4.615 1.145 ;
      RECT  6.31 0.54 6.695 0.655 ;
      RECT  6.605 0.655 6.695 0.88 ;
      RECT  6.605 0.88 6.83 0.99 ;
      RECT  6.605 0.99 6.695 1.22 ;
      RECT  6.56 1.22 6.695 1.505 ;
      RECT  5.195 0.545 5.645 0.665 ;
      RECT  5.555 0.665 5.645 0.77 ;
      RECT  5.195 0.665 5.3 1.35 ;
      RECT  5.555 0.77 5.72 0.86 ;
      RECT  5.62 0.86 5.72 1.02 ;
      RECT  5.195 1.35 5.39 1.47 ;
      RECT  5.195 1.47 5.285 1.56 ;
      RECT  3.745 0.965 3.975 1.065 ;
      RECT  3.885 1.065 3.975 1.235 ;
      RECT  3.885 1.235 4.545 1.335 ;
      RECT  4.455 1.335 4.545 1.56 ;
      RECT  4.455 1.56 5.285 1.66 ;
      RECT  5.735 0.55 5.915 0.67 ;
      RECT  5.825 0.67 5.915 1.28 ;
      RECT  5.76 1.28 5.915 1.505 ;
      RECT  6.01 0.52 6.155 0.95 ;
      RECT  6.01 0.95 6.505 1.05 ;
      RECT  6.01 1.05 6.13 1.5 ;
      RECT  3.27 0.51 3.37 1.165 ;
      RECT  0.065 1.215 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.445 ;
      RECT  0.585 1.305 0.705 1.515 ;
      RECT  0.585 1.515 1.225 1.605 ;
      RECT  1.105 1.42 1.225 1.515 ;
      LAYER M2 ;
      RECT  0.805 0.35 2.12 0.45 ;
      RECT  2.32 0.35 3.85 0.45 ;
      RECT  5.01 0.35 6.2 0.45 ;
      RECT  6.1 0.45 6.2 0.55 ;
      RECT  6.1 0.55 6.49 0.65 ;
      RECT  3.23 0.55 5.915 0.65 ;
      LAYER V1 ;
      RECT  0.85 0.35 0.95 0.45 ;
      RECT  1.98 0.35 2.08 0.45 ;
      RECT  2.36 0.35 2.46 0.45 ;
      RECT  3.71 0.35 3.81 0.45 ;
      RECT  5.05 0.35 5.15 0.45 ;
      RECT  3.27 0.55 3.37 0.65 ;
      RECT  5.775 0.55 5.875 0.65 ;
      RECT  6.35 0.55 6.45 0.65 ;
  END
END SEN_FSDAO22PQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDAO22PQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&((A1&A2)|(B1&B2)))|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDAO22PQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDAO22PQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.805 ;
      RECT  0.35 0.805 0.575 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0576 ;
  END B2
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.705 7.05 1.29 ;
      RECT  5.835 0.855 6.15 0.945 ;
      RECT  6.05 0.945 6.15 1.09 ;
      LAYER M2 ;
      RECT  6.01 0.95 7.09 1.05 ;
      LAYER V1 ;
      RECT  6.95 0.95 7.05 1.05 ;
      RECT  6.05 0.95 6.15 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0975 ;
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.205 0.295 8.325 0.41 ;
      RECT  8.205 0.41 8.45 0.505 ;
      RECT  8.35 0.505 8.45 1.06 ;
      RECT  8.18 1.06 8.45 1.175 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.51 3.095 0.8 ;
      RECT  2.825 0.8 3.095 0.89 ;
      RECT  2.825 0.89 2.915 0.94 ;
      RECT  1.965 0.94 2.915 1.03 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0906 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 3.65 0.835 ;
      RECT  3.55 0.835 3.7 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.75 0.31 8.88 1.49 ;
    END
    ANTENNADIFFAREA 0.121 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.395 0.445 1.75 ;
      RECT  0.0 1.75 9.0 1.85 ;
      RECT  1.59 1.38 1.74 1.75 ;
      RECT  2.1 1.48 2.27 1.75 ;
      RECT  3.36 1.59 3.53 1.75 ;
      RECT  4.675 1.48 4.845 1.75 ;
      RECT  5.205 1.6 5.385 1.75 ;
      RECT  6.68 1.575 6.85 1.75 ;
      RECT  7.195 1.395 7.315 1.75 ;
      RECT  7.93 1.445 8.08 1.75 ;
      RECT  8.47 1.445 8.62 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      RECT  6.73 0.05 6.88 0.225 ;
      RECT  7.27 0.05 7.42 0.225 ;
      RECT  3.385 0.05 3.505 0.25 ;
      RECT  2.12 0.05 2.27 0.26 ;
      RECT  8.52 0.05 8.625 0.35 ;
      RECT  1.13 0.05 1.245 0.385 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  5.475 0.05 5.625 0.395 ;
      RECT  4.955 0.05 5.105 0.405 ;
      RECT  7.945 0.05 8.075 0.42 ;
      RECT  1.605 0.05 1.725 0.545 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.87 0.15 4.83 0.25 ;
      RECT  4.71 0.25 4.83 0.395 ;
      RECT  6.24 0.215 6.35 0.315 ;
      RECT  6.24 0.315 7.855 0.405 ;
      RECT  7.685 0.2 7.855 0.315 ;
      RECT  7.765 0.405 7.855 0.82 ;
      RECT  6.24 0.405 6.33 1.3 ;
      RECT  7.765 0.82 8.03 0.91 ;
      RECT  7.94 0.91 8.03 1.265 ;
      RECT  7.75 1.265 8.66 1.355 ;
      RECT  8.56 0.77 8.66 1.265 ;
      RECT  6.205 1.3 6.33 1.48 ;
      RECT  7.75 1.355 7.84 1.44 ;
      RECT  7.655 1.44 7.84 1.53 ;
      RECT  2.395 0.26 3.27 0.34 ;
      RECT  2.395 0.34 4.59 0.39 ;
      RECT  3.19 0.39 4.59 0.43 ;
      RECT  2.395 0.39 2.505 0.44 ;
      RECT  4.47 0.43 4.59 0.51 ;
      RECT  3.19 0.43 3.28 1.41 ;
      RECT  2.905 1.41 3.76 1.43 ;
      RECT  2.905 1.43 4.05 1.48 ;
      RECT  3.93 1.425 4.05 1.43 ;
      RECT  2.36 1.48 4.05 1.5 ;
      RECT  3.645 1.5 4.05 1.52 ;
      RECT  2.36 1.5 3.025 1.585 ;
      RECT  3.93 1.52 4.05 1.65 ;
      RECT  0.545 0.24 1.04 0.355 ;
      RECT  0.94 0.355 1.04 1.205 ;
      RECT  0.845 1.205 1.04 1.295 ;
      RECT  0.845 1.295 0.96 1.405 ;
      RECT  1.825 0.35 2.305 0.46 ;
      RECT  2.215 0.46 2.305 0.53 ;
      RECT  2.215 0.53 2.805 0.62 ;
      RECT  2.62 0.48 2.805 0.53 ;
      RECT  5.725 0.355 5.84 0.495 ;
      RECT  4.78 0.495 5.84 0.585 ;
      RECT  4.78 0.585 5.285 0.6 ;
      RECT  5.195 0.6 5.285 1.105 ;
      RECT  4.935 1.105 5.285 1.21 ;
      RECT  5.195 1.21 5.285 1.24 ;
      RECT  5.195 1.24 5.745 1.33 ;
      RECT  5.655 1.33 5.745 1.36 ;
      RECT  5.655 1.36 5.845 1.46 ;
      RECT  3.93 0.52 4.375 0.6 ;
      RECT  3.93 0.6 4.69 0.62 ;
      RECT  4.285 0.62 4.69 0.69 ;
      RECT  3.93 0.62 4.02 1.24 ;
      RECT  4.6 0.69 4.96 0.78 ;
      RECT  4.87 0.78 4.96 0.88 ;
      RECT  4.87 0.88 5.105 0.99 ;
      RECT  3.93 1.24 4.32 1.335 ;
      RECT  4.2 1.335 4.32 1.52 ;
      RECT  6.715 0.495 7.19 0.615 ;
      RECT  6.715 0.615 6.805 0.815 ;
      RECT  6.655 0.815 6.805 0.985 ;
      RECT  6.715 0.985 6.805 1.395 ;
      RECT  6.425 1.395 7.055 1.485 ;
      RECT  6.425 1.485 6.515 1.57 ;
      RECT  6.94 1.485 7.055 1.605 ;
      RECT  4.34 0.87 4.73 0.97 ;
      RECT  4.64 0.97 4.73 1.3 ;
      RECT  4.64 1.3 5.06 1.39 ;
      RECT  4.97 1.39 5.06 1.42 ;
      RECT  4.97 1.42 5.565 1.51 ;
      RECT  5.475 1.51 5.565 1.57 ;
      RECT  5.475 1.57 6.515 1.66 ;
      RECT  3.37 0.52 3.84 0.62 ;
      RECT  3.37 0.62 3.46 1.21 ;
      RECT  3.37 1.21 3.84 1.32 ;
      RECT  7.945 0.51 8.045 0.625 ;
      RECT  7.945 0.625 8.255 0.715 ;
      RECT  8.155 0.715 8.255 0.925 ;
      RECT  6.44 0.52 6.62 0.64 ;
      RECT  6.44 0.64 6.555 1.305 ;
      RECT  1.945 0.55 2.125 0.65 ;
      RECT  2.025 0.65 2.125 0.75 ;
      RECT  2.025 0.75 2.735 0.85 ;
      RECT  5.99 0.255 6.105 0.675 ;
      RECT  5.655 0.675 6.105 0.765 ;
      RECT  5.655 0.765 5.745 1.055 ;
      RECT  5.39 1.055 5.935 1.15 ;
      RECT  5.845 1.15 5.935 1.18 ;
      RECT  5.845 1.18 6.065 1.27 ;
      RECT  5.945 1.27 6.065 1.48 ;
      RECT  7.555 0.615 7.675 1.0 ;
      RECT  7.555 1.0 7.85 1.09 ;
      RECT  7.75 1.09 7.85 1.17 ;
      RECT  7.555 1.09 7.66 1.255 ;
      RECT  7.465 1.255 7.66 1.345 ;
      RECT  7.465 1.345 7.565 1.615 ;
      RECT  4.11 0.735 4.2 1.06 ;
      RECT  4.11 1.06 4.54 1.15 ;
      RECT  4.44 1.15 4.54 1.31 ;
      RECT  1.34 0.51 1.45 1.12 ;
      RECT  1.34 1.12 3.1 1.21 ;
      RECT  1.76 0.65 1.85 1.12 ;
      RECT  3.005 0.98 3.1 1.12 ;
      RECT  1.34 1.21 1.45 1.61 ;
      RECT  7.355 0.51 7.455 1.165 ;
      RECT  0.065 1.215 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.445 ;
      RECT  0.585 1.305 0.705 1.52 ;
      RECT  0.585 1.52 1.225 1.61 ;
      RECT  1.105 1.42 1.225 1.52 ;
      RECT  1.83 1.3 2.81 1.39 ;
      LAYER M2 ;
      RECT  0.9 0.55 2.125 0.65 ;
      RECT  5.955 0.55 8.085 0.65 ;
      RECT  4.4 1.15 6.58 1.25 ;
      LAYER V1 ;
      RECT  0.94 0.55 1.04 0.65 ;
      RECT  1.985 0.55 2.085 0.65 ;
      RECT  5.995 0.55 6.095 0.65 ;
      RECT  7.355 0.55 7.455 0.65 ;
      RECT  7.945 0.55 8.045 0.65 ;
      RECT  4.44 1.15 4.54 1.25 ;
      RECT  6.44 1.15 6.54 1.25 ;
  END
END SEN_FSDAO22PQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDAO22PQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&((A1&A2)|(B1&B2)))|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDAO22PQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDAO22PQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.785 ;
      RECT  0.35 0.785 0.575 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.705 8.05 1.29 ;
      RECT  6.59 0.625 6.69 0.95 ;
      RECT  6.59 0.95 7.005 1.05 ;
      RECT  6.875 0.84 7.005 0.95 ;
      LAYER M2 ;
      RECT  6.825 0.95 8.09 1.05 ;
      LAYER V1 ;
      RECT  7.95 0.95 8.05 1.05 ;
      RECT  6.865 0.95 6.965 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1263 ;
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.135 0.41 9.85 0.53 ;
      RECT  9.75 0.53 9.85 1.06 ;
      RECT  9.125 1.06 9.85 1.175 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 0.71 ;
      RECT  2.95 0.71 3.25 0.9 ;
      RECT  2.95 0.9 3.04 0.94 ;
      RECT  1.965 0.94 3.04 1.03 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1149 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.25 0.885 ;
      RECT  3.75 0.885 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.15 0.31 10.335 0.49 ;
      RECT  10.245 0.49 10.335 1.11 ;
      RECT  10.15 1.11 10.335 1.49 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.395 0.445 1.75 ;
      RECT  0.0 1.75 10.4 1.85 ;
      RECT  1.59 1.375 1.74 1.75 ;
      RECT  2.1 1.49 2.27 1.75 ;
      RECT  3.6 1.6 3.77 1.75 ;
      RECT  5.12 1.48 5.29 1.75 ;
      RECT  5.64 1.48 5.81 1.75 ;
      RECT  7.55 1.575 7.72 1.75 ;
      RECT  8.145 1.39 8.265 1.75 ;
      RECT  8.9 1.445 9.05 1.75 ;
      RECT  9.42 1.445 9.57 1.75 ;
      RECT  9.94 1.445 10.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.4 0.05 ;
      RECT  7.715 0.05 7.835 0.225 ;
      RECT  8.255 0.05 8.375 0.225 ;
      RECT  2.135 0.05 2.255 0.26 ;
      RECT  3.625 0.05 3.745 0.265 ;
      RECT  9.41 0.05 9.58 0.32 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  5.4 0.05 5.55 0.405 ;
      RECT  5.92 0.05 6.07 0.405 ;
      RECT  1.13 0.05 1.245 0.41 ;
      RECT  8.915 0.05 9.045 0.415 ;
      RECT  9.955 0.05 10.06 0.575 ;
      RECT  1.605 0.05 1.725 0.595 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  6.195 0.17 6.87 0.26 ;
      RECT  6.7 0.26 6.87 0.335 ;
      RECT  6.195 0.26 6.31 0.495 ;
      RECT  5.2 0.495 6.31 0.615 ;
      RECT  6.08 0.615 6.17 1.09 ;
      RECT  5.405 1.035 5.525 1.09 ;
      RECT  5.405 1.09 6.17 1.21 ;
      RECT  6.08 1.21 6.17 1.355 ;
      RECT  6.08 1.355 6.68 1.47 ;
      RECT  4.065 0.15 5.275 0.265 ;
      RECT  5.155 0.265 5.275 0.38 ;
      RECT  0.54 0.24 1.04 0.355 ;
      RECT  0.94 0.355 1.04 1.205 ;
      RECT  0.845 1.205 1.04 1.295 ;
      RECT  0.845 1.295 0.96 1.4 ;
      RECT  2.615 0.24 3.43 0.355 ;
      RECT  2.615 0.355 4.785 0.36 ;
      RECT  3.34 0.36 4.785 0.445 ;
      RECT  4.67 0.445 4.785 0.615 ;
      RECT  3.34 0.445 3.43 1.42 ;
      RECT  3.16 1.42 4.01 1.49 ;
      RECT  2.605 1.49 4.01 1.51 ;
      RECT  3.92 1.51 4.01 1.57 ;
      RECT  2.605 1.51 3.275 1.6 ;
      RECT  3.92 1.57 4.505 1.66 ;
      RECT  4.385 1.455 4.505 1.57 ;
      RECT  6.96 0.255 7.075 0.425 ;
      RECT  6.4 0.425 7.075 0.53 ;
      RECT  6.4 0.53 6.5 0.77 ;
      RECT  6.26 0.77 6.5 0.86 ;
      RECT  6.26 0.86 6.365 1.14 ;
      RECT  6.26 1.14 6.915 1.265 ;
      RECT  1.825 0.35 2.525 0.45 ;
      RECT  1.825 0.45 3.045 0.46 ;
      RECT  2.405 0.46 3.045 0.54 ;
      RECT  2.925 0.54 3.045 0.62 ;
      RECT  7.685 0.495 8.16 0.615 ;
      RECT  7.685 0.615 7.775 0.765 ;
      RECT  7.57 0.765 7.775 0.935 ;
      RECT  7.685 0.935 7.775 1.395 ;
      RECT  7.135 1.395 8.01 1.485 ;
      RECT  7.135 1.485 7.225 1.57 ;
      RECT  7.89 1.485 8.01 1.595 ;
      RECT  4.755 0.91 5.305 1.0 ;
      RECT  5.215 1.0 5.305 1.3 ;
      RECT  5.215 1.3 5.99 1.39 ;
      RECT  5.9 1.39 5.99 1.57 ;
      RECT  5.9 1.57 7.225 1.66 ;
      RECT  8.915 0.51 9.015 0.625 ;
      RECT  8.915 0.625 9.19 0.715 ;
      RECT  9.09 0.715 9.19 0.795 ;
      RECT  9.09 0.795 9.605 0.905 ;
      RECT  7.39 0.52 7.59 0.64 ;
      RECT  7.39 0.64 7.48 0.8 ;
      RECT  7.275 0.8 7.48 0.89 ;
      RECT  7.275 0.89 7.39 1.305 ;
      RECT  1.985 0.55 2.25 0.65 ;
      RECT  2.15 0.65 2.25 0.75 ;
      RECT  2.15 0.75 2.805 0.85 ;
      RECT  3.525 0.55 4.065 0.66 ;
      RECT  3.525 0.66 3.615 1.21 ;
      RECT  3.525 1.21 4.04 1.33 ;
      RECT  4.375 0.555 4.515 0.73 ;
      RECT  4.375 0.73 5.575 0.77 ;
      RECT  4.93 0.375 5.04 0.73 ;
      RECT  4.375 0.77 5.9 0.82 ;
      RECT  5.49 0.82 5.9 0.88 ;
      RECT  4.375 0.82 4.465 1.27 ;
      RECT  4.13 1.27 4.79 1.365 ;
      RECT  4.13 1.365 4.245 1.48 ;
      RECT  1.775 0.67 1.895 0.84 ;
      RECT  1.775 0.84 1.865 1.12 ;
      RECT  1.34 0.51 1.45 1.12 ;
      RECT  1.34 1.12 3.25 1.21 ;
      RECT  3.15 1.035 3.25 1.12 ;
      RECT  1.34 1.21 1.45 1.585 ;
      RECT  9.965 0.77 10.155 0.94 ;
      RECT  9.965 0.94 10.055 1.265 ;
      RECT  7.21 0.21 7.335 0.315 ;
      RECT  7.21 0.315 8.825 0.405 ;
      RECT  8.655 0.2 8.825 0.315 ;
      RECT  7.21 0.405 7.3 0.62 ;
      RECT  8.735 0.405 8.825 0.82 ;
      RECT  7.095 0.62 7.3 0.71 ;
      RECT  7.095 0.71 7.185 1.145 ;
      RECT  8.735 0.82 9.0 0.91 ;
      RECT  8.91 0.91 9.0 1.265 ;
      RECT  7.015 1.145 7.185 1.265 ;
      RECT  8.66 1.265 10.055 1.355 ;
      RECT  8.66 1.355 8.77 1.61 ;
      RECT  8.325 0.51 8.425 1.0 ;
      RECT  8.525 0.615 8.645 1.0 ;
      RECT  8.525 1.0 8.82 1.09 ;
      RECT  8.405 1.09 8.82 1.11 ;
      RECT  8.405 1.11 8.625 1.18 ;
      RECT  8.405 1.18 8.525 1.62 ;
      RECT  4.555 0.935 4.645 1.09 ;
      RECT  4.555 1.09 5.125 1.18 ;
      RECT  5.025 1.18 5.125 1.32 ;
      RECT  0.065 1.215 0.705 1.305 ;
      RECT  0.065 1.305 0.185 1.44 ;
      RECT  0.585 1.305 0.705 1.52 ;
      RECT  0.585 1.52 1.225 1.61 ;
      RECT  1.105 1.385 1.225 1.52 ;
      RECT  1.84 1.3 3.07 1.4 ;
      LAYER M2 ;
      RECT  0.9 0.55 2.165 0.65 ;
      RECT  6.36 0.55 9.055 0.65 ;
      RECT  4.985 1.15 7.415 1.25 ;
      LAYER V1 ;
      RECT  0.94 0.55 1.04 0.65 ;
      RECT  2.025 0.55 2.125 0.65 ;
      RECT  6.4 0.55 6.5 0.65 ;
      RECT  8.325 0.55 8.425 0.65 ;
      RECT  8.915 0.55 9.015 0.65 ;
      RECT  5.025 1.15 5.125 1.25 ;
      RECT  7.275 1.15 7.375 1.25 ;
  END
END SEN_FSDAO22PQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNQ_D_1
#      Description : "D-Flip Flop w/scan, neg-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDNQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.7 1.65 0.8 ;
      RECT  1.55 0.8 1.85 0.97 ;
      RECT  1.75 0.97 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.3 5.49 0.59 ;
      RECT  5.35 0.59 5.45 1.21 ;
      RECT  5.35 1.21 5.49 1.5 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.405 1.05 0.495 ;
      RECT  0.95 0.495 1.05 0.6 ;
      RECT  0.26 0.495 0.355 0.75 ;
      RECT  0.95 0.6 1.145 0.8 ;
      RECT  0.245 0.75 0.355 0.97 ;
      RECT  0.95 0.8 1.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.305 0.6 1.45 0.91 ;
      RECT  1.15 0.91 1.45 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.24 0.44 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  1.425 1.615 1.605 1.75 ;
      RECT  1.885 1.615 2.065 1.75 ;
      RECT  3.31 1.425 3.45 1.75 ;
      RECT  4.58 1.405 4.71 1.75 ;
      RECT  5.11 1.2 5.23 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  1.895 0.05 2.075 0.185 ;
      RECT  0.295 0.05 0.475 0.305 ;
      RECT  1.375 0.05 1.555 0.305 ;
      RECT  4.595 0.05 4.71 0.4 ;
      RECT  3.28 0.05 3.41 0.59 ;
      RECT  5.11 0.05 5.23 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.485 0.16 2.605 0.285 ;
      RECT  1.68 0.285 2.605 0.375 ;
      RECT  1.68 0.375 1.77 0.395 ;
      RECT  0.8 0.215 1.25 0.305 ;
      RECT  1.16 0.305 1.25 0.395 ;
      RECT  1.16 0.395 1.77 0.485 ;
      RECT  3.89 0.225 4.505 0.325 ;
      RECT  4.415 0.325 4.505 0.72 ;
      RECT  4.415 0.72 4.765 0.85 ;
      RECT  4.08 0.85 4.765 0.94 ;
      RECT  4.08 0.94 4.17 1.415 ;
      RECT  4.08 1.415 4.23 1.64 ;
      RECT  2.69 0.43 2.93 0.53 ;
      RECT  2.84 0.53 2.93 0.705 ;
      RECT  2.84 0.705 3.525 0.795 ;
      RECT  3.36 0.795 3.525 0.955 ;
      RECT  2.84 0.795 2.93 1.44 ;
      RECT  3.52 0.47 3.715 0.57 ;
      RECT  3.625 0.57 3.715 1.045 ;
      RECT  3.115 1.045 3.81 1.135 ;
      RECT  3.72 1.135 3.81 1.44 ;
      RECT  1.74 0.575 2.105 0.665 ;
      RECT  2.015 0.665 2.105 1.2 ;
      RECT  1.595 1.2 2.105 1.305 ;
      RECT  0.45 0.61 0.64 0.73 ;
      RECT  0.55 0.73 0.64 1.06 ;
      RECT  0.065 0.16 0.18 0.36 ;
      RECT  0.065 0.36 0.155 1.06 ;
      RECT  0.065 1.06 0.64 1.15 ;
      RECT  0.55 1.15 0.64 1.55 ;
      RECT  0.065 1.15 0.185 1.64 ;
      RECT  0.55 1.55 1.185 1.64 ;
      RECT  3.9 0.545 4.325 0.74 ;
      RECT  3.9 0.74 3.99 0.75 ;
      RECT  3.815 0.75 3.99 0.955 ;
      RECT  3.9 0.955 3.99 1.55 ;
      RECT  3.09 1.245 3.63 1.335 ;
      RECT  3.09 1.335 3.18 1.55 ;
      RECT  3.54 1.335 3.63 1.55 ;
      RECT  2.3 0.485 2.42 0.68 ;
      RECT  2.3 0.68 2.75 0.79 ;
      RECT  2.3 0.79 2.41 0.935 ;
      RECT  2.66 0.79 2.75 1.55 ;
      RECT  2.235 0.935 2.41 1.05 ;
      RECT  2.235 1.05 2.355 1.345 ;
      RECT  2.66 1.55 3.18 1.64 ;
      RECT  3.54 1.55 3.99 1.64 ;
      RECT  4.855 0.27 4.97 0.755 ;
      RECT  4.855 0.755 5.17 0.925 ;
      RECT  4.855 0.925 4.965 1.12 ;
      RECT  4.36 1.12 4.965 1.22 ;
      RECT  4.845 1.22 4.965 1.48 ;
      RECT  0.94 1.25 1.07 1.35 ;
      RECT  0.94 1.35 1.385 1.435 ;
      RECT  0.94 1.435 2.57 1.46 ;
      RECT  2.47 1.29 2.57 1.435 ;
      RECT  1.295 1.46 2.57 1.525 ;
  END
END SEN_FSDNQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNQ_D_2
#      Description : "D-Flip Flop w/scan, neg-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDNQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.8 ;
      RECT  1.55 0.8 1.85 0.97 ;
      RECT  1.75 0.97 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.5 5.46 1.3 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.405 1.05 0.495 ;
      RECT  0.95 0.495 1.05 0.6 ;
      RECT  0.26 0.495 0.355 0.75 ;
      RECT  0.95 0.6 1.145 0.8 ;
      RECT  0.245 0.75 0.355 0.97 ;
      RECT  0.95 0.8 1.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.305 0.6 1.45 0.91 ;
      RECT  1.15 0.91 1.45 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.24 0.44 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  1.425 1.615 1.605 1.75 ;
      RECT  1.885 1.615 2.065 1.75 ;
      RECT  3.34 1.435 3.45 1.75 ;
      RECT  4.58 1.41 4.71 1.75 ;
      RECT  5.095 1.2 5.215 1.75 ;
      RECT  5.615 1.21 5.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  1.895 0.05 2.075 0.185 ;
      RECT  0.295 0.05 0.475 0.305 ;
      RECT  1.375 0.05 1.555 0.305 ;
      RECT  4.595 0.05 4.71 0.4 ;
      RECT  3.28 0.05 3.41 0.575 ;
      RECT  5.615 0.05 5.735 0.59 ;
      RECT  5.095 0.05 5.215 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.485 0.16 2.605 0.285 ;
      RECT  1.68 0.285 2.605 0.375 ;
      RECT  1.68 0.375 1.77 0.395 ;
      RECT  0.8 0.215 1.25 0.305 ;
      RECT  1.16 0.305 1.25 0.395 ;
      RECT  1.16 0.395 1.77 0.485 ;
      RECT  3.93 0.225 4.505 0.325 ;
      RECT  4.415 0.325 4.505 0.71 ;
      RECT  4.415 0.71 4.765 0.85 ;
      RECT  4.08 0.85 4.765 0.94 ;
      RECT  4.08 0.94 4.185 1.64 ;
      RECT  2.69 0.43 2.93 0.53 ;
      RECT  2.84 0.53 2.93 0.705 ;
      RECT  2.84 0.705 3.525 0.795 ;
      RECT  3.36 0.795 3.525 0.955 ;
      RECT  2.84 0.795 2.95 1.46 ;
      RECT  3.52 0.45 3.715 0.55 ;
      RECT  3.625 0.55 3.715 1.045 ;
      RECT  3.12 1.045 3.81 1.135 ;
      RECT  3.72 1.135 3.81 1.44 ;
      RECT  1.74 0.575 2.105 0.665 ;
      RECT  2.015 0.665 2.105 1.2 ;
      RECT  1.595 1.2 2.105 1.305 ;
      RECT  3.9 0.51 4.325 0.735 ;
      RECT  3.9 0.735 3.99 0.75 ;
      RECT  3.815 0.75 3.99 0.955 ;
      RECT  3.9 0.955 3.99 1.55 ;
      RECT  3.08 1.245 3.63 1.335 ;
      RECT  3.08 1.335 3.19 1.55 ;
      RECT  3.54 1.335 3.63 1.55 ;
      RECT  2.3 0.485 2.42 0.68 ;
      RECT  2.3 0.68 2.75 0.79 ;
      RECT  2.3 0.79 2.41 0.935 ;
      RECT  2.66 0.79 2.75 1.55 ;
      RECT  2.235 0.935 2.41 1.05 ;
      RECT  2.235 1.05 2.355 1.345 ;
      RECT  2.66 1.55 3.19 1.64 ;
      RECT  3.54 1.55 3.99 1.64 ;
      RECT  0.455 0.605 0.64 0.78 ;
      RECT  0.55 0.78 0.64 1.06 ;
      RECT  0.065 0.16 0.18 0.36 ;
      RECT  0.065 0.36 0.155 1.06 ;
      RECT  0.065 1.06 0.64 1.15 ;
      RECT  0.55 1.15 0.64 1.55 ;
      RECT  0.065 1.15 0.185 1.64 ;
      RECT  0.55 1.55 1.185 1.64 ;
      RECT  4.855 0.34 4.965 0.79 ;
      RECT  4.855 0.79 5.24 0.89 ;
      RECT  4.855 0.89 4.965 1.12 ;
      RECT  4.36 1.12 4.965 1.22 ;
      RECT  4.845 1.22 4.965 1.38 ;
      RECT  0.94 1.25 1.045 1.35 ;
      RECT  0.94 1.35 1.385 1.435 ;
      RECT  0.94 1.435 2.57 1.46 ;
      RECT  2.47 1.29 2.57 1.435 ;
      RECT  1.295 1.46 2.57 1.525 ;
  END
END SEN_FSDNQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNQ_D_4
#      Description : "D-Flip Flop w/scan, neg-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDNQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 0.71 ;
      RECT  1.55 0.71 1.945 0.89 ;
      RECT  1.55 0.89 1.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.4 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.36 0.51 6.05 0.69 ;
      RECT  5.95 0.69 6.05 1.11 ;
      RECT  5.385 1.11 6.09 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.65 0.435 ;
      RECT  0.26 0.435 1.1 0.51 ;
      RECT  0.26 0.51 1.25 0.525 ;
      RECT  0.95 0.525 1.25 0.69 ;
      RECT  0.26 0.525 0.355 0.73 ;
      RECT  0.95 0.69 1.05 1.095 ;
      RECT  0.245 0.73 0.355 0.94 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.2 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.24 0.45 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  1.49 1.6 1.67 1.75 ;
      RECT  1.85 1.6 2.03 1.75 ;
      RECT  3.395 1.435 3.52 1.75 ;
      RECT  4.665 1.24 4.785 1.75 ;
      RECT  5.175 1.21 5.295 1.75 ;
      RECT  5.69 1.41 5.82 1.75 ;
      RECT  6.215 1.21 6.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  1.405 0.05 1.585 0.2 ;
      RECT  2.105 0.05 2.285 0.2 ;
      RECT  0.31 0.05 0.48 0.22 ;
      RECT  5.675 0.05 5.805 0.39 ;
      RECT  4.615 0.05 4.735 0.545 ;
      RECT  5.145 0.05 5.265 0.59 ;
      RECT  6.21 0.05 6.33 0.59 ;
      RECT  3.505 0.05 3.625 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.84 0.235 1.3 0.31 ;
      RECT  0.84 0.31 2.82 0.325 ;
      RECT  2.7 0.16 2.82 0.31 ;
      RECT  1.21 0.325 2.82 0.4 ;
      RECT  4.02 0.225 4.445 0.325 ;
      RECT  4.355 0.325 4.445 0.655 ;
      RECT  4.355 0.655 4.875 0.745 ;
      RECT  4.78 0.745 4.875 0.93 ;
      RECT  4.355 0.745 4.445 1.3 ;
      RECT  4.15 1.3 4.445 1.39 ;
      RECT  4.15 1.39 4.255 1.63 ;
      RECT  4.825 0.425 5.055 0.525 ;
      RECT  4.965 0.525 5.055 0.79 ;
      RECT  4.965 0.79 5.84 0.89 ;
      RECT  4.965 0.89 5.065 1.04 ;
      RECT  4.555 0.835 4.645 1.04 ;
      RECT  4.555 1.04 5.065 1.13 ;
      RECT  4.925 1.13 5.065 1.26 ;
      RECT  1.795 0.5 2.21 0.59 ;
      RECT  2.11 0.59 2.21 1.12 ;
      RECT  1.74 1.12 2.21 1.21 ;
      RECT  3.765 0.49 3.98 0.59 ;
      RECT  3.765 0.59 3.88 1.075 ;
      RECT  3.28 0.885 3.445 1.075 ;
      RECT  3.28 1.075 3.88 1.165 ;
      RECT  3.79 1.165 3.88 1.44 ;
      RECT  2.98 0.35 3.07 0.705 ;
      RECT  2.98 0.705 3.675 0.795 ;
      RECT  3.585 0.795 3.675 0.965 ;
      RECT  2.98 0.795 3.075 1.28 ;
      RECT  2.91 1.28 3.075 1.46 ;
      RECT  0.445 0.635 0.635 0.8 ;
      RECT  0.545 0.8 0.635 1.06 ;
      RECT  0.065 0.19 0.17 0.44 ;
      RECT  0.065 0.44 0.155 1.06 ;
      RECT  0.065 1.06 0.635 1.15 ;
      RECT  0.54 1.15 0.635 1.55 ;
      RECT  0.065 1.15 0.185 1.64 ;
      RECT  0.54 1.55 1.215 1.64 ;
      RECT  4.13 0.505 4.255 0.8 ;
      RECT  3.97 0.8 4.255 0.97 ;
      RECT  3.97 0.97 4.06 1.55 ;
      RECT  3.17 1.255 3.7 1.345 ;
      RECT  3.17 1.345 3.26 1.55 ;
      RECT  3.61 1.345 3.7 1.55 ;
      RECT  2.445 0.525 2.82 0.625 ;
      RECT  2.73 0.625 2.82 0.95 ;
      RECT  2.33 0.95 2.82 1.07 ;
      RECT  2.33 1.07 2.44 1.185 ;
      RECT  2.73 1.07 2.82 1.55 ;
      RECT  2.73 1.55 3.26 1.64 ;
      RECT  3.61 1.55 4.06 1.64 ;
      RECT  0.94 1.21 1.045 1.335 ;
      RECT  0.94 1.335 1.415 1.4 ;
      RECT  0.94 1.4 2.635 1.43 ;
      RECT  1.325 1.43 2.635 1.49 ;
      RECT  2.53 1.49 2.635 1.62 ;
  END
END SEN_FSDNQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDNQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.905 0.14 4.665 0.235 ;
      RECT  4.495 0.235 4.665 0.27 ;
      RECT  3.905 0.235 3.995 0.71 ;
      RECT  3.625 0.71 3.995 0.89 ;
      RECT  3.625 0.89 3.85 0.925 ;
      RECT  3.75 0.925 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0885 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.795 ;
      RECT  0.75 0.795 0.985 0.965 ;
      RECT  0.75 0.965 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.195 6.34 0.395 ;
      RECT  6.15 0.395 6.26 1.19 ;
      RECT  6.15 1.19 6.34 1.375 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.795 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0714 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.445 0.465 1.05 0.555 ;
      RECT  0.95 0.555 1.05 0.615 ;
      RECT  0.445 0.555 0.55 0.685 ;
      RECT  0.95 0.615 1.25 0.705 ;
      RECT  1.15 0.705 1.25 1.03 ;
      RECT  1.15 1.03 1.465 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.74 0.31 5.85 1.49 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.61 0.545 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  1.485 1.515 1.6 1.75 ;
      RECT  2.88 1.44 3.0 1.75 ;
      RECT  3.675 1.48 3.845 1.75 ;
      RECT  5.075 1.605 5.245 1.75 ;
      RECT  5.43 1.605 5.6 1.75 ;
      RECT  5.955 1.425 6.075 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  4.945 0.05 5.065 0.275 ;
      RECT  5.455 0.05 5.575 0.275 ;
      RECT  1.34 0.05 1.46 0.345 ;
      RECT  0.3 0.05 0.47 0.375 ;
      RECT  5.955 0.05 6.06 0.41 ;
      RECT  2.835 0.05 3.005 0.455 ;
      RECT  3.7 0.05 3.815 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.56 0.14 2.23 0.23 ;
      RECT  2.06 0.23 2.23 0.355 ;
      RECT  1.56 0.23 1.65 0.435 ;
      RECT  0.72 0.255 1.245 0.375 ;
      RECT  1.155 0.375 1.245 0.435 ;
      RECT  1.155 0.435 1.65 0.525 ;
      RECT  1.56 0.525 1.65 1.305 ;
      RECT  0.91 1.305 1.65 1.335 ;
      RECT  0.91 1.335 2.02 1.425 ;
      RECT  1.93 1.425 2.02 1.465 ;
      RECT  1.93 1.465 2.175 1.565 ;
      RECT  4.68 0.365 5.575 0.455 ;
      RECT  4.68 0.455 4.79 0.615 ;
      RECT  5.485 0.455 5.575 0.78 ;
      RECT  5.485 0.78 5.625 0.95 ;
      RECT  5.485 0.95 5.575 1.425 ;
      RECT  4.885 1.425 5.575 1.465 ;
      RECT  4.78 1.465 5.575 1.515 ;
      RECT  4.78 1.515 4.975 1.555 ;
      RECT  4.385 0.415 4.56 0.505 ;
      RECT  4.385 0.505 4.475 0.81 ;
      RECT  4.385 0.81 4.575 0.91 ;
      RECT  4.475 0.91 4.575 1.05 ;
      RECT  4.475 1.05 4.645 1.14 ;
      RECT  1.95 0.45 2.54 0.54 ;
      RECT  1.95 0.54 2.04 0.975 ;
      RECT  1.95 0.975 2.38 1.065 ;
      RECT  2.29 1.065 2.38 1.17 ;
      RECT  3.15 0.33 3.26 0.545 ;
      RECT  2.73 0.545 3.26 0.635 ;
      RECT  2.73 0.635 2.82 0.655 ;
      RECT  2.205 0.655 2.82 0.745 ;
      RECT  2.205 0.745 2.58 0.755 ;
      RECT  2.205 0.755 2.295 0.84 ;
      RECT  2.49 0.755 2.58 1.065 ;
      RECT  2.49 1.065 3.26 1.16 ;
      RECT  3.165 0.985 3.26 1.065 ;
      RECT  5.115 0.545 5.395 0.68 ;
      RECT  5.115 0.68 5.205 0.86 ;
      RECT  4.87 0.86 5.205 0.965 ;
      RECT  5.115 0.965 5.205 1.225 ;
      RECT  3.445 0.44 3.535 0.73 ;
      RECT  2.91 0.73 3.535 0.82 ;
      RECT  3.445 0.82 3.535 1.26 ;
      RECT  3.445 1.26 4.83 1.35 ;
      RECT  4.735 1.13 4.83 1.26 ;
      RECT  3.445 1.35 4.235 1.39 ;
      RECT  4.11 0.345 4.21 1.0 ;
      RECT  3.975 1.0 4.21 1.075 ;
      RECT  3.975 1.075 4.385 1.17 ;
      RECT  1.74 0.32 1.86 1.155 ;
      RECT  1.74 1.155 2.2 1.245 ;
      RECT  2.11 1.245 2.2 1.26 ;
      RECT  2.11 1.26 3.335 1.35 ;
      RECT  3.245 1.35 3.335 1.49 ;
      RECT  2.655 1.35 2.765 1.61 ;
      RECT  3.245 1.49 3.37 1.66 ;
      RECT  5.94 0.72 6.04 1.195 ;
      RECT  5.295 0.77 5.395 1.235 ;
      RECT  0.065 0.24 0.185 1.43 ;
      RECT  0.065 1.43 0.78 1.52 ;
      RECT  0.67 1.52 0.78 1.545 ;
      RECT  0.065 1.52 0.2 1.595 ;
      RECT  0.67 1.545 1.265 1.65 ;
      LAYER M2 ;
      RECT  4.435 0.95 6.08 1.05 ;
      LAYER V1 ;
      RECT  4.475 0.95 4.575 1.05 ;
      RECT  5.295 0.95 5.395 1.05 ;
      RECT  5.94 0.95 6.04 1.05 ;
  END
END SEN_FSDNQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDNQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.62 0.675 5.45 0.77 ;
      RECT  4.62 0.77 4.85 0.89 ;
      RECT  5.35 0.77 5.45 1.05 ;
      RECT  5.35 1.05 5.88 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1131 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.69 0.85 0.795 ;
      RECT  0.75 0.795 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0816 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.31 8.085 0.505 ;
      RECT  7.95 0.505 8.25 0.595 ;
      RECT  8.15 0.595 8.25 1.11 ;
      RECT  7.95 1.11 8.25 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.275 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.084 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.685 2.65 0.9 ;
      RECT  2.35 0.9 2.65 1.09 ;
      RECT  2.55 1.09 2.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.31 7.305 0.48 ;
      RECT  7.15 0.48 7.25 0.87 ;
      RECT  7.15 0.87 7.33 0.96 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.615 0.48 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  1.375 1.395 1.495 1.75 ;
      RECT  2.405 1.63 2.575 1.75 ;
      RECT  3.885 1.405 4.005 1.75 ;
      RECT  4.415 1.4 4.54 1.75 ;
      RECT  5.185 1.59 5.355 1.75 ;
      RECT  6.875 1.62 7.045 1.75 ;
      RECT  7.705 1.44 7.825 1.75 ;
      RECT  8.215 1.41 8.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  1.84 0.05 2.01 0.25 ;
      RECT  5.195 0.05 5.365 0.35 ;
      RECT  2.625 0.05 2.745 0.38 ;
      RECT  0.07 0.05 0.21 0.39 ;
      RECT  8.215 0.05 8.345 0.39 ;
      RECT  3.885 0.05 4.005 0.42 ;
      RECT  6.91 0.05 7.035 0.43 ;
      RECT  4.675 0.05 4.795 0.46 ;
      RECT  7.705 0.05 7.825 0.63 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.57 0.175 1.49 0.27 ;
      RECT  0.57 0.27 0.67 0.435 ;
      RECT  0.57 0.435 0.66 1.01 ;
      RECT  0.57 1.01 1.995 1.1 ;
      RECT  0.57 1.1 1.02 1.125 ;
      RECT  1.905 1.1 1.995 1.45 ;
      RECT  1.87 1.45 2.79 1.48 ;
      RECT  1.87 1.48 3.225 1.54 ;
      RECT  2.72 1.54 3.225 1.595 ;
      RECT  1.87 1.54 1.98 1.63 ;
      RECT  3.33 0.225 3.57 0.335 ;
      RECT  3.33 0.335 3.42 0.96 ;
      RECT  3.33 0.96 4.115 1.05 ;
      RECT  4.025 0.835 4.115 0.96 ;
      RECT  3.33 1.05 3.42 1.21 ;
      RECT  2.365 0.19 2.485 0.345 ;
      RECT  1.945 0.345 2.485 0.36 ;
      RECT  0.79 0.36 2.485 0.435 ;
      RECT  0.79 0.435 2.015 0.45 ;
      RECT  2.86 0.25 3.06 0.355 ;
      RECT  2.97 0.355 3.06 0.86 ;
      RECT  2.84 0.86 3.06 0.95 ;
      RECT  2.84 0.95 2.93 1.19 ;
      RECT  2.765 1.19 2.93 1.3 ;
      RECT  2.765 1.3 3.625 1.36 ;
      RECT  3.535 1.18 3.625 1.3 ;
      RECT  2.86 1.36 3.625 1.39 ;
      RECT  0.335 0.2 0.455 0.37 ;
      RECT  0.365 0.37 0.455 1.215 ;
      RECT  0.365 1.215 1.815 1.305 ;
      RECT  1.725 1.19 1.815 1.215 ;
      RECT  1.64 1.305 1.815 1.36 ;
      RECT  1.64 1.36 1.75 1.625 ;
      RECT  6.56 0.25 6.79 0.37 ;
      RECT  6.7 0.37 6.79 0.565 ;
      RECT  6.7 0.565 7.055 0.655 ;
      RECT  6.955 0.655 7.055 0.795 ;
      RECT  6.7 0.655 6.79 1.015 ;
      RECT  6.56 1.015 6.79 1.135 ;
      RECT  4.905 0.44 5.83 0.56 ;
      RECT  5.74 0.56 5.83 0.87 ;
      RECT  5.74 0.87 6.08 0.96 ;
      RECT  5.99 0.96 6.08 1.305 ;
      RECT  5.99 1.305 6.2 1.315 ;
      RECT  5.35 1.315 6.2 1.4 ;
      RECT  4.89 1.4 6.2 1.405 ;
      RECT  4.89 1.405 5.46 1.5 ;
      RECT  2.57 0.47 2.88 0.595 ;
      RECT  2.745 0.595 2.88 0.77 ;
      RECT  4.165 0.435 4.3 0.605 ;
      RECT  4.21 0.605 4.3 1.14 ;
      RECT  3.795 1.14 4.3 1.22 ;
      RECT  3.795 1.22 5.12 1.31 ;
      RECT  5.03 0.86 5.12 1.22 ;
      RECT  1.0 0.54 2.305 0.64 ;
      RECT  5.97 0.445 6.125 0.78 ;
      RECT  3.565 0.43 3.71 0.87 ;
      RECT  7.675 0.785 8.06 0.895 ;
      RECT  7.675 0.895 7.765 1.26 ;
      RECT  7.475 1.26 7.765 1.35 ;
      RECT  7.475 1.35 7.565 1.44 ;
      RECT  6.215 0.175 6.305 1.01 ;
      RECT  6.215 1.01 6.445 1.13 ;
      RECT  6.325 1.13 6.445 1.44 ;
      RECT  6.325 1.44 7.565 1.53 ;
      RECT  6.325 1.53 6.445 1.545 ;
      RECT  5.71 1.545 6.445 1.66 ;
      RECT  6.395 0.51 6.535 0.9 ;
      RECT  4.42 0.23 4.525 1.02 ;
      RECT  4.42 1.02 4.86 1.13 ;
      RECT  3.15 0.315 3.24 1.04 ;
      RECT  3.07 1.04 3.24 1.21 ;
      RECT  7.445 0.19 7.545 1.08 ;
      RECT  7.295 1.08 7.545 1.17 ;
      RECT  7.295 1.17 7.385 1.24 ;
      RECT  6.665 1.24 7.385 1.35 ;
      RECT  0.065 1.3 0.185 1.395 ;
      RECT  0.065 1.395 1.26 1.525 ;
      RECT  1.15 1.525 1.26 1.61 ;
      LAYER M2 ;
      RECT  2.71 0.55 6.575 0.65 ;
      LAYER V1 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  3.565 0.55 3.665 0.65 ;
      RECT  4.42 0.55 4.52 0.65 ;
      RECT  6.025 0.55 6.125 0.65 ;
      RECT  6.435 0.55 6.535 0.65 ;
  END
END SEN_FSDNQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDNQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.05 0.82 ;
      RECT  5.75 0.82 6.05 0.89 ;
      RECT  5.15 0.82 5.25 0.92 ;
      RECT  5.95 0.89 6.05 1.045 ;
      RECT  5.95 1.045 6.705 1.135 ;
      RECT  6.615 0.965 6.705 1.045 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1506 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.82 ;
      RECT  0.75 0.82 2.25 0.92 ;
      RECT  2.15 0.92 2.25 1.305 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.35 0.3 9.465 0.47 ;
      RECT  8.815 0.47 9.465 0.59 ;
      RECT  9.35 0.59 9.465 1.11 ;
      RECT  8.825 1.11 9.465 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.48 0.275 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0993 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 2.65 0.7 ;
      RECT  2.35 0.7 2.65 0.79 ;
      RECT  2.35 0.79 2.45 1.31 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.07 0.285 8.17 0.435 ;
      RECT  8.07 0.435 8.25 0.53 ;
      RECT  8.15 0.53 8.25 0.865 ;
      RECT  8.025 0.865 8.25 0.965 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.615 0.48 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  1.375 1.435 1.495 1.75 ;
      RECT  2.42 1.63 2.59 1.75 ;
      RECT  4.35 1.425 4.52 1.75 ;
      RECT  4.87 1.425 5.04 1.75 ;
      RECT  5.4 1.425 5.57 1.75 ;
      RECT  5.69 1.15 5.81 1.75 ;
      RECT  6.185 1.485 6.355 1.75 ;
      RECT  7.765 1.58 7.935 1.75 ;
      RECT  8.57 1.44 8.7 1.75 ;
      RECT  9.1 1.385 9.22 1.75 ;
      RECT  9.61 1.41 9.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  1.855 0.05 2.025 0.21 ;
      RECT  9.08 0.05 9.23 0.38 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  2.635 0.05 2.805 0.39 ;
      RECT  4.94 0.05 5.06 0.39 ;
      RECT  5.97 0.05 6.09 0.39 ;
      RECT  9.61 0.05 9.74 0.39 ;
      RECT  7.79 0.05 7.91 0.415 ;
      RECT  4.42 0.05 4.54 0.425 ;
      RECT  5.45 0.05 5.57 0.445 ;
      RECT  8.58 0.05 8.7 0.63 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.56 0.14 1.51 0.23 ;
      RECT  0.56 0.23 0.68 0.37 ;
      RECT  0.56 0.37 0.655 1.04 ;
      RECT  0.56 1.04 2.06 1.13 ;
      RECT  0.56 1.13 1.56 1.165 ;
      RECT  1.97 1.13 2.06 1.435 ;
      RECT  1.84 1.435 2.06 1.45 ;
      RECT  1.84 1.45 2.935 1.48 ;
      RECT  1.84 1.48 3.94 1.54 ;
      RECT  2.865 1.54 3.94 1.595 ;
      RECT  3.185 0.155 3.81 0.245 ;
      RECT  3.71 0.245 3.81 0.495 ;
      RECT  3.185 0.245 3.29 1.21 ;
      RECT  2.405 0.21 2.505 0.335 ;
      RECT  0.795 0.335 2.505 0.43 ;
      RECT  8.315 0.19 8.465 0.36 ;
      RECT  8.37 0.36 8.465 1.07 ;
      RECT  7.77 1.07 8.465 1.17 ;
      RECT  7.77 1.17 7.86 1.21 ;
      RECT  7.56 1.21 7.86 1.3 ;
      RECT  0.34 0.19 0.455 0.39 ;
      RECT  0.365 0.39 0.455 1.255 ;
      RECT  0.365 1.255 1.87 1.345 ;
      RECT  1.7 1.23 1.87 1.255 ;
      RECT  1.65 1.345 1.74 1.63 ;
      RECT  2.895 0.27 3.095 0.39 ;
      RECT  3.005 0.39 3.095 1.19 ;
      RECT  2.775 1.19 3.095 1.3 ;
      RECT  2.775 1.3 4.12 1.36 ;
      RECT  3.005 1.36 4.12 1.39 ;
      RECT  4.03 1.39 4.12 1.595 ;
      RECT  7.495 0.285 7.68 0.4 ;
      RECT  7.59 0.4 7.68 0.6 ;
      RECT  7.59 0.6 8.01 0.69 ;
      RECT  7.92 0.69 8.01 0.77 ;
      RECT  7.59 0.69 7.68 0.955 ;
      RECT  7.49 0.955 7.68 1.06 ;
      RECT  5.21 0.31 5.31 0.48 ;
      RECT  4.945 0.48 5.31 0.57 ;
      RECT  4.945 0.57 5.045 1.045 ;
      RECT  4.945 1.045 5.325 1.155 ;
      RECT  6.745 0.415 6.915 0.505 ;
      RECT  6.825 0.505 6.915 0.785 ;
      RECT  5.715 0.365 5.825 0.48 ;
      RECT  5.715 0.48 6.335 0.585 ;
      RECT  6.23 0.31 6.335 0.48 ;
      RECT  6.245 0.585 6.335 0.785 ;
      RECT  6.245 0.785 6.915 0.875 ;
      RECT  6.825 0.875 6.915 1.285 ;
      RECT  5.925 1.285 7.155 1.395 ;
      RECT  3.94 0.2 4.04 0.62 ;
      RECT  3.94 0.62 4.605 0.71 ;
      RECT  4.515 0.71 4.605 0.915 ;
      RECT  3.94 0.71 4.035 1.08 ;
      RECT  3.44 0.335 3.55 1.08 ;
      RECT  3.44 1.08 4.035 1.21 ;
      RECT  1.045 0.52 2.295 0.625 ;
      RECT  7.2 0.55 7.455 0.65 ;
      RECT  7.355 0.65 7.455 0.87 ;
      RECT  6.45 0.47 6.655 0.695 ;
      RECT  8.575 0.79 9.255 0.89 ;
      RECT  8.575 0.89 8.665 1.26 ;
      RECT  8.32 1.26 8.665 1.35 ;
      RECT  8.32 1.35 8.41 1.4 ;
      RECT  6.45 0.215 7.39 0.325 ;
      RECT  7.01 0.325 7.1 0.96 ;
      RECT  7.01 0.96 7.365 1.06 ;
      RECT  7.265 1.06 7.365 1.4 ;
      RECT  7.265 1.4 8.41 1.485 ;
      RECT  6.68 1.485 8.41 1.49 ;
      RECT  6.68 1.49 7.355 1.58 ;
      RECT  2.815 0.51 2.915 0.93 ;
      RECT  2.63 0.93 2.915 1.02 ;
      RECT  5.485 0.91 5.655 1.0 ;
      RECT  5.485 1.0 5.575 1.245 ;
      RECT  4.25 0.855 4.34 1.215 ;
      RECT  4.25 1.215 4.79 1.245 ;
      RECT  4.695 0.3 4.79 1.215 ;
      RECT  4.25 1.245 5.575 1.335 ;
      RECT  0.065 1.285 0.185 1.435 ;
      RECT  0.065 1.435 1.25 1.525 ;
      RECT  1.16 1.525 1.25 1.64 ;
      LAYER M2 ;
      RECT  2.775 0.55 7.38 0.65 ;
      LAYER V1 ;
      RECT  2.815 0.55 2.915 0.65 ;
      RECT  4.945 0.55 5.045 0.65 ;
      RECT  6.49 0.55 6.59 0.65 ;
      RECT  7.24 0.55 7.34 0.65 ;
  END
END SEN_FSDNQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNRBQ_1
#      Description : "D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNRBQ_1
  CLASS CORE ;
  FOREIGN SEN_FSDNRBQ_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.655 4.65 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0357 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.51 7.09 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.04 0.29 6.14 0.51 ;
      RECT  6.04 0.51 6.37 0.69 ;
      RECT  6.27 0.69 6.37 0.925 ;
      RECT  3.255 0.29 3.355 0.55 ;
      RECT  3.255 0.55 3.49 0.65 ;
      RECT  1.55 0.31 1.65 0.77 ;
      RECT  1.55 0.77 1.83 0.86 ;
      LAYER M2 ;
      RECT  1.51 0.35 6.18 0.45 ;
      LAYER V1 ;
      RECT  6.04 0.35 6.14 0.45 ;
      RECT  3.255 0.35 3.355 0.45 ;
      RECT  1.55 0.35 1.65 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0684 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.92 0.51 2.02 0.76 ;
      RECT  1.92 0.76 2.09 0.86 ;
      RECT  0.47 0.35 0.65 0.45 ;
      RECT  0.55 0.45 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.47 0.35 1.41 0.45 ;
      RECT  1.31 0.45 1.41 0.55 ;
      RECT  1.31 0.55 2.06 0.65 ;
      LAYER V1 ;
      RECT  1.92 0.55 2.02 0.65 ;
      RECT  0.51 0.35 0.61 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.65 1.13 1.87 1.33 ;
      RECT  0.15 0.51 0.25 1.29 ;
      LAYER M2 ;
      RECT  0.11 1.15 1.87 1.25 ;
      LAYER V1 ;
      RECT  1.73 1.15 1.83 1.25 ;
      RECT  0.15 1.15 0.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  0.595 1.57 0.715 1.75 ;
      RECT  1.83 1.61 2.0 1.75 ;
      RECT  3.19 1.615 3.36 1.75 ;
      RECT  3.485 1.615 3.655 1.75 ;
      RECT  4.275 1.615 4.445 1.75 ;
      RECT  4.795 1.615 4.965 1.75 ;
      RECT  6.07 1.56 6.24 1.75 ;
      RECT  6.715 1.375 6.835 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  4.24 0.05 4.36 0.385 ;
      RECT  4.79 0.05 4.91 0.385 ;
      RECT  6.23 0.05 6.33 0.385 ;
      RECT  3.47 0.05 3.59 0.41 ;
      RECT  1.79 0.05 1.91 0.415 ;
      RECT  6.715 0.05 6.835 0.65 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.065 0.14 1.435 0.23 ;
      RECT  0.065 0.23 0.185 0.39 ;
      RECT  1.315 0.23 1.435 0.475 ;
      RECT  2.625 0.255 3.165 0.345 ;
      RECT  3.075 0.345 3.165 0.74 ;
      RECT  2.625 0.345 2.73 1.16 ;
      RECT  3.075 0.74 3.69 0.83 ;
      RECT  3.585 0.83 3.69 0.98 ;
      RECT  3.255 0.83 3.345 1.165 ;
      RECT  6.42 0.24 6.59 0.36 ;
      RECT  6.5 0.36 6.59 1.015 ;
      RECT  6.04 0.87 6.13 1.015 ;
      RECT  6.04 1.015 6.59 1.105 ;
      RECT  3.99 0.28 4.105 0.485 ;
      RECT  4.015 0.485 4.105 1.435 ;
      RECT  2.805 1.435 5.375 1.525 ;
      RECT  5.285 1.525 5.375 1.555 ;
      RECT  2.805 1.525 2.915 1.66 ;
      RECT  5.285 1.555 5.515 1.645 ;
      RECT  3.74 0.28 3.84 0.55 ;
      RECT  3.74 0.55 3.925 0.65 ;
      RECT  3.835 0.65 3.925 1.255 ;
      RECT  3.045 0.93 3.155 1.255 ;
      RECT  3.045 1.255 3.925 1.345 ;
      RECT  5.27 0.45 5.95 0.55 ;
      RECT  5.86 0.55 5.95 1.195 ;
      RECT  5.58 1.195 6.845 1.285 ;
      RECT  6.755 0.755 6.845 1.195 ;
      RECT  5.58 1.285 5.67 1.48 ;
      RECT  2.13 0.48 2.27 0.675 ;
      RECT  2.18 0.675 2.27 0.95 ;
      RECT  1.255 0.72 1.345 0.95 ;
      RECT  1.255 0.95 2.27 1.04 ;
      RECT  2.13 1.04 2.27 1.17 ;
      RECT  5.245 0.715 5.345 0.795 ;
      RECT  5.245 0.795 5.77 0.885 ;
      RECT  5.67 0.685 5.77 0.795 ;
      RECT  5.35 0.885 5.45 1.255 ;
      RECT  4.49 0.18 4.61 0.475 ;
      RECT  4.195 0.475 4.61 0.565 ;
      RECT  4.195 0.565 4.285 1.255 ;
      RECT  4.195 1.255 5.45 1.345 ;
      RECT  4.875 0.475 4.975 0.955 ;
      RECT  5.065 0.41 5.155 0.975 ;
      RECT  5.065 0.975 5.21 1.145 ;
      RECT  0.75 0.415 0.85 1.2 ;
      RECT  0.75 1.2 1.48 1.29 ;
      RECT  1.39 1.29 1.48 1.43 ;
      RECT  1.39 1.43 2.46 1.52 ;
      RECT  2.37 0.25 2.46 1.43 ;
      RECT  1.39 1.52 1.48 1.57 ;
      RECT  0.82 1.57 1.48 1.66 ;
      RECT  2.84 0.465 2.94 1.25 ;
      RECT  2.55 1.25 2.94 1.34 ;
      RECT  2.55 1.34 2.65 1.66 ;
      RECT  5.8 1.375 6.54 1.465 ;
      RECT  0.325 1.39 1.26 1.48 ;
      RECT  0.325 1.48 0.445 1.585 ;
      LAYER M2 ;
      RECT  3.745 0.55 5.015 0.65 ;
      RECT  2.8 1.15 5.49 1.25 ;
      LAYER V1 ;
      RECT  3.785 0.55 3.885 0.65 ;
      RECT  4.875 0.55 4.975 0.65 ;
      RECT  2.84 1.15 2.94 1.25 ;
      RECT  5.35 1.15 5.45 1.25 ;
  END
END SEN_FSDNRBQ_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNRBQ_2
#      Description : "D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNRBQ_2
  CLASS CORE ;
  FOREIGN SEN_FSDNRBQ_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.05 0.89 ;
      RECT  4.75 0.89 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.705 0.85 0.91 ;
      RECT  0.75 0.91 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 0.31 8.65 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.55 0.29 7.65 0.51 ;
      RECT  7.55 0.51 7.85 0.69 ;
      RECT  3.905 0.31 4.005 0.575 ;
      RECT  3.905 0.575 4.17 0.685 ;
      RECT  2.95 0.31 3.05 0.71 ;
      RECT  2.55 0.71 3.05 0.89 ;
      LAYER M2 ;
      RECT  2.91 0.35 7.69 0.45 ;
      LAYER V1 ;
      RECT  7.55 0.35 7.65 0.45 ;
      RECT  3.905 0.35 4.005 0.45 ;
      RECT  2.95 0.35 3.05 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0876 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.27 0.51 2.37 1.03 ;
      RECT  0.405 0.51 0.51 0.91 ;
      RECT  0.405 0.91 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.365 0.55 2.41 0.65 ;
      LAYER V1 ;
      RECT  2.27 0.55 2.37 0.65 ;
      RECT  0.405 0.55 0.505 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0849 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.89 0.8 1.99 1.31 ;
      RECT  0.15 0.71 0.25 1.29 ;
      LAYER M2 ;
      RECT  0.11 1.15 2.03 1.25 ;
      LAYER V1 ;
      RECT  1.89 1.15 1.99 1.25 ;
      RECT  0.15 1.15 0.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0276 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 9.0 1.85 ;
      RECT  0.585 1.45 0.705 1.75 ;
      RECT  2.07 1.615 2.24 1.75 ;
      RECT  3.905 1.575 4.01 1.75 ;
      RECT  4.19 1.575 4.31 1.75 ;
      RECT  4.73 1.575 4.85 1.75 ;
      RECT  5.28 1.575 5.4 1.75 ;
      RECT  6.085 1.575 6.205 1.75 ;
      RECT  7.735 1.615 7.905 1.75 ;
      RECT  8.28 1.43 8.4 1.75 ;
      RECT  8.81 1.21 8.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      RECT  2.32 0.05 2.49 0.185 ;
      RECT  2.86 0.05 3.03 0.215 ;
      RECT  4.095 0.05 4.2 0.36 ;
      RECT  6.19 0.05 6.305 0.39 ;
      RECT  7.74 0.05 7.86 0.39 ;
      RECT  4.64 0.05 4.76 0.425 ;
      RECT  5.15 0.05 5.27 0.425 ;
      RECT  5.67 0.05 5.79 0.435 ;
      RECT  8.28 0.05 8.4 0.59 ;
      RECT  8.81 0.05 8.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.56 0.2 2.17 0.275 ;
      RECT  1.56 0.275 2.725 0.32 ;
      RECT  2.08 0.32 2.725 0.395 ;
      RECT  2.625 0.395 2.725 0.51 ;
      RECT  0.78 0.225 1.47 0.325 ;
      RECT  1.38 0.325 1.47 0.415 ;
      RECT  1.38 0.415 1.99 0.515 ;
      RECT  6.395 0.22 7.375 0.325 ;
      RECT  7.285 0.325 7.375 0.81 ;
      RECT  7.285 0.81 7.56 0.9 ;
      RECT  7.47 0.9 7.56 1.25 ;
      RECT  7.285 1.25 8.445 1.34 ;
      RECT  8.355 0.725 8.445 1.25 ;
      RECT  7.285 1.34 7.375 1.38 ;
      RECT  6.615 1.38 7.375 1.48 ;
      RECT  4.31 0.23 4.54 0.34 ;
      RECT  4.44 0.34 4.54 0.55 ;
      RECT  4.44 0.55 4.63 0.65 ;
      RECT  4.54 0.65 4.63 1.21 ;
      RECT  3.725 0.96 3.815 1.21 ;
      RECT  3.725 1.21 4.63 1.3 ;
      RECT  0.065 0.2 0.185 0.35 ;
      RECT  0.065 0.35 0.33 0.45 ;
      RECT  3.34 0.25 3.815 0.35 ;
      RECT  3.725 0.35 3.815 0.775 ;
      RECT  3.34 0.35 3.43 1.21 ;
      RECT  3.725 0.775 4.43 0.865 ;
      RECT  3.91 0.865 4.03 1.12 ;
      RECT  2.74 1.21 3.43 1.3 ;
      RECT  2.74 1.3 2.845 1.425 ;
      RECT  5.41 0.215 5.53 0.385 ;
      RECT  5.41 0.385 5.5 1.395 ;
      RECT  3.725 1.395 6.41 1.485 ;
      RECT  3.725 1.485 3.815 1.57 ;
      RECT  6.32 1.485 6.41 1.57 ;
      RECT  3.365 1.57 3.815 1.66 ;
      RECT  6.32 1.57 6.985 1.66 ;
      RECT  6.54 0.42 6.86 0.51 ;
      RECT  6.54 0.51 6.63 1.015 ;
      RECT  5.94 0.44 6.04 1.01 ;
      RECT  5.79 1.01 6.04 1.015 ;
      RECT  5.79 1.015 7.015 1.105 ;
      RECT  6.925 0.9 7.015 1.015 ;
      RECT  4.9 0.21 5.02 0.53 ;
      RECT  4.9 0.53 5.25 0.62 ;
      RECT  5.15 0.62 5.25 1.2 ;
      RECT  4.96 1.2 5.25 1.29 ;
      RECT  2.085 0.51 2.18 0.61 ;
      RECT  1.55 0.61 2.18 0.7 ;
      RECT  1.55 0.7 1.65 0.9 ;
      RECT  2.09 0.7 2.18 1.255 ;
      RECT  2.09 1.255 2.47 1.345 ;
      RECT  2.37 1.16 2.47 1.255 ;
      RECT  6.145 0.5 6.255 0.71 ;
      RECT  6.145 0.71 6.45 0.89 ;
      RECT  6.73 0.67 7.195 0.76 ;
      RECT  7.105 0.76 7.195 0.99 ;
      RECT  7.105 0.99 7.38 1.16 ;
      RECT  7.105 1.16 7.195 1.2 ;
      RECT  5.6 1.11 5.7 1.2 ;
      RECT  5.6 1.2 7.195 1.29 ;
      RECT  8.01 0.215 8.13 0.81 ;
      RECT  7.65 0.81 8.13 0.98 ;
      RECT  8.01 0.98 8.13 1.16 ;
      RECT  3.15 0.38 3.24 1.03 ;
      RECT  2.56 1.03 3.24 1.12 ;
      RECT  2.56 1.12 2.65 1.435 ;
      RECT  0.47 0.3 0.69 0.415 ;
      RECT  0.6 0.415 0.69 0.42 ;
      RECT  0.6 0.42 1.285 0.535 ;
      RECT  1.195 0.535 1.285 0.665 ;
      RECT  1.195 0.665 1.455 0.755 ;
      RECT  1.365 0.755 1.455 1.09 ;
      RECT  1.365 1.09 1.73 1.18 ;
      RECT  1.64 1.18 1.73 1.435 ;
      RECT  1.64 1.435 2.65 1.525 ;
      RECT  1.64 1.525 1.73 1.57 ;
      RECT  1.105 1.45 1.225 1.57 ;
      RECT  1.105 1.57 1.73 1.66 ;
      RECT  0.34 1.27 1.48 1.36 ;
      RECT  1.37 1.36 1.48 1.48 ;
      RECT  0.34 1.36 0.44 1.485 ;
      RECT  0.85 1.36 0.96 1.485 ;
      RECT  3.535 0.47 3.635 1.39 ;
      RECT  2.945 1.39 3.635 1.48 ;
      RECT  2.945 1.48 3.055 1.625 ;
      RECT  7.465 1.43 8.175 1.525 ;
      LAYER M2 ;
      RECT  0.11 0.35 2.765 0.45 ;
      RECT  4.44 0.55 6.29 0.65 ;
      RECT  3.495 1.15 5.745 1.25 ;
      LAYER V1 ;
      RECT  0.15 0.35 0.25 0.45 ;
      RECT  2.625 0.35 2.725 0.45 ;
      RECT  4.48 0.55 4.58 0.65 ;
      RECT  6.15 0.55 6.25 0.65 ;
      RECT  3.535 1.15 3.635 1.25 ;
      RECT  5.15 1.15 5.25 1.25 ;
      RECT  5.6 1.15 5.7 1.25 ;
  END
END SEN_FSDNRBQ_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNRBQ_4
#      Description : "D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNRBQ_4
  CLASS CORE ;
  FOREIGN SEN_FSDNRBQ_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.25 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0714 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.885 ;
      RECT  0.75 0.885 1.18 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.35 0.51 10.05 0.69 ;
      RECT  9.95 0.69 10.05 1.11 ;
      RECT  9.35 1.11 10.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.34 0.29 8.44 0.54 ;
      RECT  8.34 0.54 8.685 0.65 ;
      RECT  4.305 0.2 4.405 0.51 ;
      RECT  4.305 0.51 4.45 0.74 ;
      RECT  3.185 0.29 3.285 0.83 ;
      RECT  2.56 0.83 3.285 0.92 ;
      LAYER M2 ;
      RECT  3.145 0.35 8.48 0.45 ;
      LAYER V1 ;
      RECT  8.34 0.35 8.44 0.45 ;
      RECT  4.305 0.35 4.405 0.45 ;
      RECT  3.185 0.35 3.285 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.114 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.55 2.53 0.65 ;
      RECT  2.35 0.65 2.45 1.085 ;
      RECT  0.35 0.49 0.45 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.31 0.55 2.53 0.65 ;
      LAYER V1 ;
      RECT  2.39 0.55 2.49 0.65 ;
      RECT  0.35 0.55 0.45 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.95 2.07 1.345 ;
      RECT  0.15 0.6 0.25 1.29 ;
      LAYER M2 ;
      RECT  0.11 1.15 2.09 1.25 ;
      LAYER V1 ;
      RECT  1.95 1.15 2.05 1.25 ;
      RECT  0.15 1.15 0.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0393 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 10.4 1.85 ;
      RECT  0.56 1.495 0.73 1.75 ;
      RECT  2.075 1.615 2.245 1.75 ;
      RECT  4.115 1.615 4.285 1.75 ;
      RECT  4.86 1.615 5.03 1.75 ;
      RECT  5.425 1.615 5.595 1.75 ;
      RECT  6.26 1.615 6.43 1.75 ;
      RECT  6.8 1.615 6.97 1.75 ;
      RECT  8.485 1.615 8.655 1.75 ;
      RECT  9.16 1.44 9.28 1.75 ;
      RECT  9.68 1.38 9.8 1.75 ;
      RECT  10.21 1.21 10.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.4 0.05 ;
      RECT  2.335 0.05 2.505 0.26 ;
      RECT  4.495 0.05 4.585 0.385 ;
      RECT  5.0 0.05 5.12 0.385 ;
      RECT  6.03 0.05 6.15 0.4 ;
      RECT  6.55 0.05 6.67 0.4 ;
      RECT  7.07 0.05 7.19 0.4 ;
      RECT  9.68 0.05 9.8 0.42 ;
      RECT  8.53 0.05 8.645 0.43 ;
      RECT  5.51 0.05 5.63 0.435 ;
      RECT  10.21 0.05 10.33 0.59 ;
      RECT  9.14 0.05 9.26 0.65 ;
      RECT  2.975 0.05 3.095 0.685 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.065 0.17 1.775 0.26 ;
      RECT  1.655 0.26 1.775 0.35 ;
      RECT  0.065 0.26 0.185 0.44 ;
      RECT  1.655 0.35 2.86 0.45 ;
      RECT  3.555 0.235 4.215 0.335 ;
      RECT  4.125 0.335 4.215 1.07 ;
      RECT  3.555 0.335 3.645 1.21 ;
      RECT  4.125 1.07 4.645 1.16 ;
      RECT  4.555 0.77 4.645 1.07 ;
      RECT  2.755 1.21 3.645 1.3 ;
      RECT  2.755 1.3 2.86 1.43 ;
      RECT  0.83 0.35 1.54 0.44 ;
      RECT  1.45 0.44 1.54 0.56 ;
      RECT  1.45 0.56 2.06 0.65 ;
      RECT  5.77 0.315 5.9 0.485 ;
      RECT  5.8 0.485 5.9 0.965 ;
      RECT  5.54 0.965 5.9 1.055 ;
      RECT  5.54 1.055 5.63 1.435 ;
      RECT  3.925 1.435 7.15 1.525 ;
      RECT  3.925 1.525 4.015 1.57 ;
      RECT  7.06 1.525 7.15 1.57 ;
      RECT  3.45 1.57 4.015 1.66 ;
      RECT  7.06 1.57 7.815 1.66 ;
      RECT  5.265 0.315 5.375 0.525 ;
      RECT  5.265 0.525 5.45 0.615 ;
      RECT  5.35 0.615 5.45 0.775 ;
      RECT  5.35 0.775 5.71 0.875 ;
      RECT  5.35 0.875 5.45 1.255 ;
      RECT  5.13 1.255 5.45 1.345 ;
      RECT  6.265 0.49 7.76 0.585 ;
      RECT  6.94 0.585 7.03 1.015 ;
      RECT  5.99 1.015 7.765 1.105 ;
      RECT  3.735 0.48 4.005 0.59 ;
      RECT  3.735 0.59 3.835 1.39 ;
      RECT  3.155 1.39 3.835 1.48 ;
      RECT  3.155 1.48 3.245 1.66 ;
      RECT  6.05 0.51 6.15 0.71 ;
      RECT  6.05 0.71 6.73 0.89 ;
      RECT  2.16 0.58 2.25 0.77 ;
      RECT  1.615 0.77 2.25 0.86 ;
      RECT  1.615 0.86 1.785 0.925 ;
      RECT  2.16 0.86 2.25 1.255 ;
      RECT  2.16 1.255 2.485 1.345 ;
      RECT  2.395 1.175 2.485 1.255 ;
      RECT  7.24 0.69 7.945 0.8 ;
      RECT  7.855 0.8 7.945 1.075 ;
      RECT  7.855 1.075 8.21 1.165 ;
      RECT  8.11 0.965 8.21 1.075 ;
      RECT  7.855 1.165 7.945 1.21 ;
      RECT  5.72 1.15 5.9 1.21 ;
      RECT  5.72 1.21 7.945 1.3 ;
      RECT  9.09 0.785 9.84 0.895 ;
      RECT  9.09 0.895 9.18 1.255 ;
      RECT  7.295 0.25 8.125 0.35 ;
      RECT  8.035 0.35 8.125 0.75 ;
      RECT  8.035 0.75 8.39 0.85 ;
      RECT  8.3 0.85 8.39 1.255 ;
      RECT  8.035 1.255 9.18 1.345 ;
      RECT  8.035 1.345 8.125 1.39 ;
      RECT  7.3 1.39 8.125 1.48 ;
      RECT  3.375 0.19 3.465 1.03 ;
      RECT  2.575 1.03 3.465 1.12 ;
      RECT  2.575 1.12 2.665 1.435 ;
      RECT  0.57 0.53 1.36 0.62 ;
      RECT  1.27 0.62 1.36 1.135 ;
      RECT  1.27 1.135 1.735 1.225 ;
      RECT  1.645 1.225 1.735 1.435 ;
      RECT  1.645 1.435 2.665 1.495 ;
      RECT  1.05 1.495 2.665 1.525 ;
      RECT  1.05 1.525 1.735 1.59 ;
      RECT  8.48 0.75 8.58 1.07 ;
      RECT  8.48 1.07 8.955 1.16 ;
      RECT  8.855 0.19 8.955 1.07 ;
      RECT  3.925 0.74 4.015 1.255 ;
      RECT  3.925 1.255 4.85 1.345 ;
      RECT  4.75 0.28 4.85 1.255 ;
      RECT  0.34 1.315 1.515 1.405 ;
      RECT  0.34 1.405 0.445 1.54 ;
      RECT  8.215 1.435 9.01 1.525 ;
      LAYER M2 ;
      RECT  4.71 0.55 6.19 0.65 ;
      RECT  3.695 1.15 5.9 1.25 ;
      LAYER V1 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  6.05 0.55 6.15 0.65 ;
      RECT  3.735 1.15 3.835 1.25 ;
      RECT  5.35 1.15 5.45 1.25 ;
      RECT  5.76 1.15 5.86 1.25 ;
  END
END SEN_FSDNRBQ_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNRBQ_D_1
#      Description : "D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNRBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDNRBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.745 ;
      RECT  1.915 0.745 2.05 0.915 ;
      RECT  1.95 0.915 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.585 0.83 0.785 0.91 ;
      RECT  0.35 0.91 0.785 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 5.93 0.68 ;
      RECT  5.75 0.68 5.85 1.31 ;
      RECT  5.75 1.31 5.93 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.91 5.09 1.29 ;
      RECT  3.855 1.035 3.955 1.31 ;
      RECT  3.525 1.31 3.955 1.41 ;
      LAYER M2 ;
      RECT  3.815 1.15 5.095 1.25 ;
      LAYER V1 ;
      RECT  4.955 1.15 5.055 1.25 ;
      RECT  3.855 1.15 3.955 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.042 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.495 ;
      RECT  0.35 0.495 1.25 0.595 ;
      RECT  0.35 0.595 0.65 0.7 ;
      RECT  1.15 0.595 1.25 0.95 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.26 0.18 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  1.28 1.54 1.45 1.75 ;
      RECT  1.935 1.57 2.06 1.75 ;
      RECT  3.325 1.515 3.495 1.75 ;
      RECT  3.78 1.5 3.95 1.75 ;
      RECT  4.9 1.43 5.005 1.75 ;
      RECT  5.485 1.235 5.6 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  1.03 0.05 1.2 0.21 ;
      RECT  1.89 0.05 2.06 0.21 ;
      RECT  3.635 0.05 3.745 0.31 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  4.835 0.05 4.965 0.39 ;
      RECT  5.545 0.05 5.675 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.835 0.14 4.285 0.23 ;
      RECT  3.835 0.23 3.925 0.415 ;
      RECT  4.195 0.23 4.285 0.655 ;
      RECT  2.68 0.14 3.375 0.23 ;
      RECT  3.275 0.23 3.375 0.415 ;
      RECT  2.68 0.23 2.78 1.03 ;
      RECT  3.275 0.415 3.925 0.505 ;
      RECT  4.195 0.655 4.315 0.765 ;
      RECT  4.225 0.765 4.315 0.95 ;
      RECT  4.225 0.95 4.63 1.05 ;
      RECT  4.53 1.05 4.63 1.275 ;
      RECT  0.555 0.18 0.675 0.3 ;
      RECT  0.555 0.3 2.575 0.39 ;
      RECT  2.445 0.16 2.575 0.3 ;
      RECT  4.375 0.19 4.495 0.36 ;
      RECT  4.405 0.36 4.495 0.725 ;
      RECT  4.405 0.725 5.31 0.815 ;
      RECT  5.205 0.815 5.31 0.925 ;
      RECT  4.72 0.815 4.81 1.365 ;
      RECT  4.37 1.365 4.81 1.455 ;
      RECT  4.37 1.455 4.49 1.63 ;
      RECT  5.3 0.22 5.42 0.48 ;
      RECT  4.68 0.48 5.505 0.61 ;
      RECT  5.415 0.61 5.505 0.755 ;
      RECT  5.415 0.755 5.65 0.925 ;
      RECT  5.415 0.925 5.505 1.015 ;
      RECT  5.295 1.015 5.505 1.105 ;
      RECT  5.295 1.105 5.385 1.45 ;
      RECT  5.12 1.45 5.385 1.57 ;
      RECT  1.545 0.515 1.795 0.635 ;
      RECT  1.695 0.635 1.795 1.38 ;
      RECT  1.64 1.38 2.24 1.47 ;
      RECT  2.15 1.47 2.24 1.57 ;
      RECT  1.64 1.47 1.76 1.62 ;
      RECT  2.15 1.57 2.575 1.66 ;
      RECT  2.87 0.36 2.985 0.635 ;
      RECT  2.87 0.635 3.91 0.725 ;
      RECT  2.87 0.725 2.975 1.415 ;
      RECT  2.265 0.525 2.58 0.715 ;
      RECT  2.265 0.715 2.4 1.14 ;
      RECT  2.265 1.14 2.78 1.23 ;
      RECT  2.69 1.23 2.78 1.57 ;
      RECT  2.69 1.57 3.185 1.66 ;
      RECT  4.015 0.34 4.105 0.835 ;
      RECT  3.2 0.835 4.135 0.925 ;
      RECT  4.045 0.925 4.135 1.23 ;
      RECT  4.045 1.23 4.23 1.4 ;
      RECT  1.35 0.5 1.445 0.99 ;
      RECT  1.35 0.99 1.605 1.16 ;
      RECT  1.35 1.16 1.445 1.2 ;
      RECT  0.905 0.705 0.995 1.2 ;
      RECT  0.905 1.2 1.445 1.3 ;
      RECT  0.905 1.3 0.995 1.57 ;
      RECT  0.345 1.57 0.995 1.66 ;
      RECT  3.115 1.035 3.765 1.125 ;
      RECT  3.655 1.125 3.765 1.21 ;
      RECT  3.115 1.125 3.235 1.38 ;
      RECT  0.685 1.2 0.785 1.34 ;
      RECT  0.53 1.34 0.785 1.46 ;
      RECT  2.33 1.32 2.6 1.48 ;
      LAYER M2 ;
      RECT  3.605 0.95 4.415 1.05 ;
      RECT  3.605 1.05 3.705 1.15 ;
      RECT  1.655 1.15 3.705 1.25 ;
      RECT  0.605 1.35 2.555 1.45 ;
      LAYER V1 ;
      RECT  4.265 0.95 4.365 1.05 ;
      RECT  1.695 1.15 1.795 1.25 ;
      RECT  0.645 1.35 0.745 1.45 ;
      RECT  2.415 1.35 2.515 1.45 ;
  END
END SEN_FSDNRBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNRBQ_D_2
#      Description : "D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNRBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDNRBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.745 ;
      RECT  1.915 0.745 2.05 0.915 ;
      RECT  1.95 0.915 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.585 0.83 0.785 0.91 ;
      RECT  0.35 0.91 0.785 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 6.05 0.69 ;
      RECT  5.95 0.69 6.05 1.11 ;
      RECT  5.75 1.11 6.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.91 5.09 1.29 ;
      RECT  3.855 1.035 3.955 1.31 ;
      RECT  3.525 1.31 3.955 1.41 ;
      LAYER M2 ;
      RECT  3.815 1.15 5.095 1.25 ;
      LAYER V1 ;
      RECT  4.955 1.15 5.055 1.25 ;
      RECT  3.855 1.15 3.955 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.495 ;
      RECT  0.35 0.495 1.25 0.595 ;
      RECT  0.35 0.595 0.65 0.7 ;
      RECT  1.15 0.595 1.25 0.945 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.26 0.18 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  1.28 1.54 1.45 1.75 ;
      RECT  1.935 1.57 2.06 1.75 ;
      RECT  3.325 1.515 3.495 1.75 ;
      RECT  3.78 1.5 3.95 1.75 ;
      RECT  4.9 1.43 5.005 1.75 ;
      RECT  5.485 1.235 5.6 1.75 ;
      RECT  6.02 1.41 6.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  1.03 0.05 1.2 0.21 ;
      RECT  1.89 0.05 2.06 0.21 ;
      RECT  3.635 0.05 3.745 0.325 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  4.855 0.05 4.985 0.39 ;
      RECT  5.5 0.05 5.63 0.39 ;
      RECT  6.02 0.05 6.145 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.835 0.14 4.285 0.23 ;
      RECT  3.835 0.23 3.925 0.415 ;
      RECT  4.195 0.23 4.285 0.655 ;
      RECT  2.68 0.14 3.375 0.23 ;
      RECT  3.275 0.23 3.375 0.415 ;
      RECT  2.68 0.23 2.78 1.03 ;
      RECT  3.275 0.415 3.925 0.505 ;
      RECT  4.195 0.655 4.315 0.765 ;
      RECT  4.225 0.765 4.315 0.95 ;
      RECT  4.225 0.95 4.63 1.05 ;
      RECT  4.53 1.05 4.63 1.265 ;
      RECT  0.555 0.18 0.675 0.3 ;
      RECT  0.555 0.3 2.575 0.39 ;
      RECT  2.445 0.16 2.575 0.3 ;
      RECT  4.375 0.19 4.495 0.36 ;
      RECT  4.405 0.36 4.495 0.725 ;
      RECT  4.405 0.725 5.31 0.815 ;
      RECT  5.205 0.815 5.31 0.925 ;
      RECT  4.72 0.815 4.81 1.365 ;
      RECT  4.37 1.365 4.81 1.455 ;
      RECT  4.37 1.455 4.49 1.63 ;
      RECT  4.65 0.48 5.505 0.61 ;
      RECT  5.415 0.61 5.505 0.785 ;
      RECT  5.415 0.785 5.86 0.895 ;
      RECT  5.415 0.895 5.505 1.015 ;
      RECT  5.295 1.015 5.505 1.105 ;
      RECT  5.295 1.105 5.385 1.45 ;
      RECT  5.12 1.45 5.385 1.57 ;
      RECT  1.545 0.515 1.795 0.635 ;
      RECT  1.695 0.635 1.795 1.38 ;
      RECT  1.64 1.38 2.24 1.47 ;
      RECT  2.15 1.47 2.24 1.57 ;
      RECT  1.64 1.47 1.76 1.62 ;
      RECT  2.15 1.57 2.575 1.66 ;
      RECT  2.87 0.36 2.985 0.635 ;
      RECT  2.87 0.635 3.91 0.725 ;
      RECT  2.87 0.725 2.975 1.415 ;
      RECT  2.265 0.525 2.58 0.715 ;
      RECT  2.265 0.715 2.4 1.14 ;
      RECT  2.265 1.14 2.78 1.23 ;
      RECT  2.69 1.23 2.78 1.57 ;
      RECT  2.69 1.57 3.185 1.66 ;
      RECT  4.015 0.35 4.105 0.835 ;
      RECT  3.17 0.835 4.135 0.925 ;
      RECT  4.045 0.925 4.135 1.23 ;
      RECT  4.045 1.23 4.23 1.4 ;
      RECT  1.35 0.5 1.445 0.99 ;
      RECT  1.35 0.99 1.605 1.16 ;
      RECT  1.35 1.16 1.445 1.2 ;
      RECT  0.905 0.71 0.995 1.2 ;
      RECT  0.905 1.2 1.445 1.3 ;
      RECT  0.905 1.3 0.995 1.57 ;
      RECT  0.345 1.57 0.995 1.66 ;
      RECT  3.115 1.035 3.765 1.125 ;
      RECT  3.655 1.125 3.765 1.21 ;
      RECT  3.115 1.125 3.235 1.38 ;
      RECT  0.685 1.2 0.785 1.34 ;
      RECT  0.53 1.34 0.785 1.46 ;
      RECT  2.33 1.32 2.6 1.48 ;
      LAYER M2 ;
      RECT  3.605 0.95 4.415 1.05 ;
      RECT  3.605 1.05 3.705 1.15 ;
      RECT  1.655 1.15 3.705 1.25 ;
      RECT  0.605 1.35 2.555 1.45 ;
      LAYER V1 ;
      RECT  4.265 0.95 4.365 1.05 ;
      RECT  1.695 1.15 1.795 1.25 ;
      RECT  0.645 1.35 0.745 1.45 ;
      RECT  2.415 1.35 2.515 1.45 ;
  END
END SEN_FSDNRBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDNRBQ_D_4
#      Description : "D-Flip Flop w/scan, neg-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=!CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDNRBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDNRBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.605 0.83 0.815 0.91 ;
      RECT  0.35 0.91 0.815 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 6.47 0.69 ;
      RECT  6.35 0.69 6.47 1.06 ;
      RECT  5.805 1.06 6.47 1.16 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.015 1.07 5.26 1.29 ;
      RECT  3.88 1.035 3.995 1.31 ;
      RECT  3.57 1.31 3.995 1.41 ;
      LAYER M2 ;
      RECT  3.84 1.15 5.155 1.25 ;
      LAYER V1 ;
      RECT  5.015 1.15 5.115 1.25 ;
      RECT  3.88 1.15 3.98 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.495 ;
      RECT  0.35 0.495 1.28 0.595 ;
      RECT  0.35 0.595 0.65 0.7 ;
      RECT  1.15 0.595 1.28 0.945 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.26 0.19 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.32 1.54 1.49 1.75 ;
      RECT  1.955 1.61 2.125 1.75 ;
      RECT  3.345 1.515 3.515 1.75 ;
      RECT  3.82 1.5 3.99 1.75 ;
      RECT  4.96 1.43 5.07 1.75 ;
      RECT  5.545 1.21 5.66 1.75 ;
      RECT  6.09 1.255 6.21 1.75 ;
      RECT  6.615 1.21 6.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  1.07 0.05 1.24 0.21 ;
      RECT  1.93 0.05 2.1 0.21 ;
      RECT  3.695 0.05 3.805 0.33 ;
      RECT  0.07 0.05 0.2 0.39 ;
      RECT  4.905 0.05 5.035 0.39 ;
      RECT  5.565 0.05 5.695 0.39 ;
      RECT  6.085 0.05 6.215 0.4 ;
      RECT  6.615 0.05 6.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.895 0.16 4.355 0.25 ;
      RECT  3.895 0.25 3.985 0.435 ;
      RECT  4.265 0.25 4.355 0.95 ;
      RECT  2.72 0.16 3.415 0.25 ;
      RECT  3.315 0.25 3.415 0.435 ;
      RECT  2.72 0.25 2.82 0.995 ;
      RECT  3.315 0.435 3.985 0.525 ;
      RECT  4.265 0.95 4.445 0.97 ;
      RECT  4.265 0.97 4.69 1.06 ;
      RECT  4.59 1.06 4.69 1.265 ;
      RECT  0.54 0.225 0.72 0.3 ;
      RECT  0.54 0.3 2.615 0.39 ;
      RECT  2.485 0.16 2.615 0.3 ;
      RECT  4.445 0.19 4.585 0.36 ;
      RECT  4.475 0.36 4.585 0.71 ;
      RECT  4.475 0.71 5.37 0.8 ;
      RECT  5.265 0.8 5.37 0.925 ;
      RECT  4.78 0.8 4.87 1.365 ;
      RECT  4.43 1.365 4.87 1.455 ;
      RECT  4.43 1.455 4.55 1.63 ;
      RECT  4.71 0.5 5.55 0.605 ;
      RECT  5.46 0.605 5.55 0.795 ;
      RECT  5.46 0.795 6.255 0.895 ;
      RECT  5.46 0.895 5.55 1.015 ;
      RECT  5.355 1.015 5.55 1.105 ;
      RECT  5.355 1.105 5.445 1.45 ;
      RECT  5.18 1.45 5.445 1.57 ;
      RECT  1.585 0.515 1.835 0.635 ;
      RECT  1.735 0.635 1.835 1.38 ;
      RECT  1.68 1.38 1.835 1.41 ;
      RECT  1.68 1.41 2.305 1.5 ;
      RECT  2.215 1.5 2.305 1.57 ;
      RECT  1.68 1.5 1.8 1.62 ;
      RECT  2.215 1.57 2.615 1.66 ;
      RECT  2.91 0.36 3.025 0.635 ;
      RECT  2.91 0.635 3.985 0.725 ;
      RECT  2.91 0.725 3.015 1.415 ;
      RECT  2.305 0.525 2.62 0.715 ;
      RECT  2.305 0.715 2.44 1.085 ;
      RECT  2.305 1.085 2.82 1.175 ;
      RECT  2.73 1.175 2.82 1.57 ;
      RECT  2.73 1.57 3.225 1.66 ;
      RECT  4.075 0.36 4.175 0.835 ;
      RECT  3.21 0.835 4.175 0.925 ;
      RECT  4.085 0.925 4.175 1.23 ;
      RECT  4.085 1.23 4.27 1.4 ;
      RECT  1.39 0.5 1.485 0.99 ;
      RECT  1.39 0.99 1.645 1.16 ;
      RECT  1.39 1.16 1.485 1.2 ;
      RECT  0.925 0.705 1.015 1.2 ;
      RECT  0.925 1.2 1.485 1.3 ;
      RECT  0.925 1.3 1.015 1.57 ;
      RECT  0.36 1.57 1.015 1.66 ;
      RECT  3.155 1.035 3.79 1.125 ;
      RECT  3.685 1.125 3.79 1.21 ;
      RECT  3.155 1.125 3.275 1.38 ;
      RECT  0.705 1.2 0.805 1.33 ;
      RECT  0.55 1.33 0.805 1.46 ;
      RECT  2.395 1.265 2.64 1.48 ;
      LAYER M2 ;
      RECT  3.64 0.95 4.455 1.05 ;
      RECT  3.64 1.05 3.74 1.15 ;
      RECT  1.695 1.15 3.74 1.25 ;
      RECT  0.53 1.35 2.595 1.45 ;
      LAYER V1 ;
      RECT  4.305 0.95 4.405 1.05 ;
      RECT  1.735 1.15 1.835 1.25 ;
      RECT  0.665 1.35 0.765 1.45 ;
      RECT  2.455 1.35 2.555 1.45 ;
  END
END SEN_FSDNRBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPC1BQ_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&D&RS)|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPC1BQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDPC1BQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.7 2.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.44 0.85 0.705 ;
      RECT  0.75 0.705 1.07 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.415 5.72 0.585 ;
      RECT  5.55 0.585 5.65 1.215 ;
      RECT  5.55 1.215 5.73 1.385 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.71 ;
      RECT  1.205 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RS
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.26 0.65 0.45 ;
      RECT  0.505 0.45 0.65 0.62 ;
      RECT  0.55 0.62 0.65 1.01 ;
      RECT  0.55 1.01 2.05 1.1 ;
      RECT  1.95 1.1 2.05 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.37 1.44 0.49 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  2.285 1.6 2.455 1.75 ;
      RECT  3.83 1.475 4.0 1.75 ;
      RECT  4.865 1.38 4.99 1.75 ;
      RECT  5.35 1.44 5.47 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  2.475 0.05 2.595 0.21 ;
      RECT  5.35 0.05 5.47 0.365 ;
      RECT  0.325 0.05 0.445 0.38 ;
      RECT  4.86 0.05 4.98 0.4 ;
      RECT  1.735 0.05 1.855 0.42 ;
      RECT  3.82 0.05 3.94 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.35 0.165 4.71 0.255 ;
      RECT  4.35 0.255 4.47 0.39 ;
      RECT  4.62 0.255 4.71 0.655 ;
      RECT  4.62 0.655 5.12 0.745 ;
      RECT  5.03 0.745 5.12 0.94 ;
      RECT  4.62 0.745 4.71 1.475 ;
      RECT  4.37 1.475 4.71 1.57 ;
      RECT  3.08 0.19 3.2 0.3 ;
      RECT  1.945 0.3 3.2 0.42 ;
      RECT  1.945 0.42 2.035 0.51 ;
      RECT  0.77 0.205 1.645 0.315 ;
      RECT  1.555 0.315 1.645 0.51 ;
      RECT  1.555 0.51 2.035 0.6 ;
      RECT  5.125 0.27 5.24 0.455 ;
      RECT  5.125 0.455 5.395 0.56 ;
      RECT  5.305 0.56 5.395 1.04 ;
      RECT  4.8 0.835 4.89 1.04 ;
      RECT  4.8 1.04 5.395 1.13 ;
      RECT  5.13 1.13 5.25 1.41 ;
      RECT  4.09 0.295 4.26 0.465 ;
      RECT  4.17 0.465 4.26 1.105 ;
      RECT  3.69 0.855 3.78 1.105 ;
      RECT  3.69 1.105 4.26 1.205 ;
      RECT  3.335 0.41 3.475 0.58 ;
      RECT  3.38 0.58 3.475 0.675 ;
      RECT  3.38 0.675 4.065 0.765 ;
      RECT  3.975 0.765 4.065 0.985 ;
      RECT  3.38 0.765 3.47 1.29 ;
      RECT  3.375 1.29 3.47 1.46 ;
      RECT  2.76 0.51 2.88 0.585 ;
      RECT  2.76 0.585 3.06 0.685 ;
      RECT  2.97 0.685 3.06 1.125 ;
      RECT  2.76 1.125 3.06 1.215 ;
      RECT  2.76 1.215 2.88 1.32 ;
      RECT  2.185 0.51 2.62 0.61 ;
      RECT  2.53 0.61 2.62 0.785 ;
      RECT  2.53 0.785 2.86 0.895 ;
      RECT  2.53 0.895 2.62 1.24 ;
      RECT  2.235 1.24 2.62 1.33 ;
      RECT  4.36 0.54 4.53 0.71 ;
      RECT  4.36 0.71 4.45 1.295 ;
      RECT  3.635 1.295 4.45 1.385 ;
      RECT  3.635 1.385 3.725 1.55 ;
      RECT  3.16 0.685 3.285 0.855 ;
      RECT  3.195 0.855 3.285 1.55 ;
      RECT  3.195 1.55 3.725 1.66 ;
      RECT  0.075 0.17 0.18 1.26 ;
      RECT  0.075 1.26 0.695 1.35 ;
      RECT  0.605 1.35 0.695 1.57 ;
      RECT  0.075 1.35 0.225 1.625 ;
      RECT  0.605 1.57 1.9 1.66 ;
      RECT  1.005 1.19 1.69 1.28 ;
      RECT  1.57 1.28 1.69 1.39 ;
      RECT  1.57 1.39 2.165 1.42 ;
      RECT  1.57 1.42 3.105 1.48 ;
      RECT  2.065 1.48 3.105 1.51 ;
      RECT  2.995 1.51 3.105 1.63 ;
      RECT  0.785 1.23 0.875 1.37 ;
      RECT  0.785 1.37 1.435 1.48 ;
  END
END SEN_FSDPC1BQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPC1BQ_D_1P5
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&D&RS)|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPC1BQ_D_1P5
  CLASS CORE ;
  FOREIGN SEN_FSDPC1BQ_D_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.7 2.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.44 0.85 0.71 ;
      RECT  0.75 0.71 1.07 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.215 5.675 0.385 ;
      RECT  5.55 0.385 5.66 1.315 ;
      RECT  5.55 1.315 5.68 1.5 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.425 1.45 0.71 ;
      RECT  1.205 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RS
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.675 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.26 0.65 0.485 ;
      RECT  0.38 0.485 0.65 0.585 ;
      RECT  0.55 0.585 0.65 1.01 ;
      RECT  0.55 1.01 1.96 1.1 ;
      RECT  1.87 1.1 1.96 1.22 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.37 1.44 0.495 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  2.215 1.6 2.385 1.75 ;
      RECT  3.78 1.495 3.95 1.75 ;
      RECT  4.82 1.415 4.94 1.75 ;
      RECT  5.295 1.405 5.415 1.75 ;
      RECT  5.815 1.33 5.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  2.425 0.05 2.545 0.21 ;
      RECT  5.295 0.05 5.415 0.38 ;
      RECT  0.325 0.05 0.445 0.39 ;
      RECT  1.745 0.05 1.865 0.405 ;
      RECT  5.815 0.05 5.935 0.43 ;
      RECT  4.81 0.05 4.93 0.515 ;
      RECT  3.77 0.05 3.89 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.035 0.18 3.145 0.3 ;
      RECT  1.955 0.3 3.145 0.42 ;
      RECT  1.955 0.42 2.045 0.495 ;
      RECT  0.77 0.21 1.63 0.31 ;
      RECT  1.54 0.31 1.63 0.495 ;
      RECT  1.54 0.495 2.045 0.585 ;
      RECT  4.275 0.315 4.66 0.42 ;
      RECT  4.57 0.42 4.66 0.72 ;
      RECT  4.57 0.72 5.07 0.81 ;
      RECT  4.98 0.81 5.07 1.03 ;
      RECT  4.57 0.81 4.66 1.495 ;
      RECT  4.3 1.495 4.66 1.595 ;
      RECT  4.045 0.25 4.16 0.485 ;
      RECT  4.045 0.485 4.21 0.58 ;
      RECT  4.12 0.58 4.21 1.12 ;
      RECT  3.64 0.865 3.73 1.12 ;
      RECT  3.64 1.12 4.21 1.225 ;
      RECT  3.29 0.41 3.425 0.58 ;
      RECT  3.33 0.58 3.425 0.675 ;
      RECT  3.33 0.675 4.015 0.765 ;
      RECT  3.925 0.765 4.015 1.01 ;
      RECT  3.33 0.765 3.42 1.29 ;
      RECT  3.325 1.29 3.42 1.46 ;
      RECT  2.71 0.51 2.83 0.585 ;
      RECT  2.71 0.585 3.015 0.685 ;
      RECT  2.925 0.685 3.015 1.09 ;
      RECT  2.71 1.09 3.015 1.185 ;
      RECT  2.71 1.185 2.83 1.33 ;
      RECT  2.135 0.52 2.57 0.61 ;
      RECT  2.48 0.61 2.57 0.785 ;
      RECT  2.48 0.785 2.81 0.895 ;
      RECT  2.48 0.895 2.57 1.24 ;
      RECT  2.185 1.24 2.57 1.33 ;
      RECT  5.045 0.515 5.29 0.625 ;
      RECT  5.2 0.625 5.29 0.785 ;
      RECT  5.2 0.785 5.44 0.895 ;
      RECT  5.2 0.895 5.29 1.195 ;
      RECT  4.75 0.905 4.84 1.195 ;
      RECT  4.75 1.195 5.29 1.3 ;
      RECT  4.3 0.54 4.48 0.73 ;
      RECT  4.3 0.73 4.39 1.315 ;
      RECT  3.585 1.315 4.39 1.405 ;
      RECT  3.585 1.405 3.675 1.55 ;
      RECT  3.12 0.67 3.21 1.245 ;
      RECT  3.12 1.245 3.235 1.335 ;
      RECT  3.145 1.335 3.235 1.55 ;
      RECT  3.145 1.55 3.675 1.66 ;
      RECT  0.075 0.165 0.175 1.26 ;
      RECT  0.075 1.26 0.69 1.35 ;
      RECT  0.6 1.35 0.69 1.57 ;
      RECT  0.075 1.35 0.22 1.625 ;
      RECT  0.6 1.57 1.85 1.66 ;
      RECT  1.005 1.19 1.625 1.28 ;
      RECT  1.53 1.28 1.625 1.39 ;
      RECT  1.53 1.39 2.115 1.42 ;
      RECT  1.53 1.42 3.055 1.48 ;
      RECT  2.015 1.48 3.055 1.51 ;
      RECT  2.945 1.51 3.055 1.63 ;
      RECT  0.78 1.23 0.88 1.37 ;
      RECT  0.78 1.37 1.435 1.48 ;
  END
END SEN_FSDPC1BQ_D_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPC1BQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&D&RS)|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPC1BQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPC1BQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.7 2.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.44 0.85 0.71 ;
      RECT  0.75 0.71 1.07 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.31 5.685 0.485 ;
      RECT  5.55 0.485 5.65 1.315 ;
      RECT  5.55 1.315 5.68 1.5 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.425 1.45 0.71 ;
      RECT  1.205 0.71 1.45 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RS
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.26 0.65 0.45 ;
      RECT  0.505 0.45 0.65 0.62 ;
      RECT  0.55 0.62 0.65 1.01 ;
      RECT  0.55 1.01 1.96 1.1 ;
      RECT  1.87 1.1 1.96 1.185 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.37 1.44 0.495 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  2.21 1.6 2.38 1.75 ;
      RECT  3.78 1.495 3.95 1.75 ;
      RECT  4.82 1.415 4.94 1.75 ;
      RECT  5.3 1.41 5.42 1.75 ;
      RECT  5.81 1.41 5.94 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  2.425 0.05 2.545 0.21 ;
      RECT  0.325 0.05 0.445 0.38 ;
      RECT  5.3 0.05 5.42 0.385 ;
      RECT  5.815 0.05 5.945 0.39 ;
      RECT  1.745 0.05 1.865 0.4 ;
      RECT  4.795 0.05 4.965 0.435 ;
      RECT  3.77 0.05 3.89 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.03 0.18 3.14 0.3 ;
      RECT  1.955 0.3 3.14 0.42 ;
      RECT  1.955 0.42 2.045 0.49 ;
      RECT  0.77 0.21 1.63 0.31 ;
      RECT  1.54 0.31 1.63 0.49 ;
      RECT  1.54 0.49 2.045 0.58 ;
      RECT  4.275 0.32 4.66 0.42 ;
      RECT  4.57 0.42 4.66 1.025 ;
      RECT  4.57 1.025 5.08 1.115 ;
      RECT  4.99 0.78 5.08 1.025 ;
      RECT  4.57 1.115 4.66 1.495 ;
      RECT  4.3 1.495 4.66 1.595 ;
      RECT  4.04 0.25 4.16 0.485 ;
      RECT  4.04 0.485 4.21 0.58 ;
      RECT  4.12 0.58 4.21 1.135 ;
      RECT  3.64 0.855 3.73 1.135 ;
      RECT  3.64 1.135 4.21 1.225 ;
      RECT  3.295 0.41 3.425 0.58 ;
      RECT  3.325 0.58 3.425 0.675 ;
      RECT  3.325 0.675 4.015 0.765 ;
      RECT  3.925 0.765 4.015 1.02 ;
      RECT  3.325 0.765 3.42 1.46 ;
      RECT  2.71 0.51 2.83 0.585 ;
      RECT  2.71 0.585 3.01 0.685 ;
      RECT  2.92 0.685 3.01 1.075 ;
      RECT  2.71 1.075 3.01 1.185 ;
      RECT  2.71 1.185 2.83 1.33 ;
      RECT  2.135 0.52 2.57 0.61 ;
      RECT  2.48 0.61 2.57 0.785 ;
      RECT  2.48 0.785 2.81 0.895 ;
      RECT  2.48 0.895 2.57 1.24 ;
      RECT  2.185 1.24 2.57 1.33 ;
      RECT  4.75 0.53 5.29 0.625 ;
      RECT  5.2 0.625 5.29 0.785 ;
      RECT  4.75 0.625 4.84 0.935 ;
      RECT  5.2 0.785 5.44 0.895 ;
      RECT  5.2 0.895 5.29 1.21 ;
      RECT  5.03 1.21 5.29 1.31 ;
      RECT  4.3 0.54 4.48 0.73 ;
      RECT  4.3 0.73 4.39 1.315 ;
      RECT  3.585 1.315 4.39 1.405 ;
      RECT  3.585 1.405 3.675 1.55 ;
      RECT  3.11 0.7 3.235 0.87 ;
      RECT  3.145 0.87 3.235 1.55 ;
      RECT  3.145 1.55 3.675 1.66 ;
      RECT  0.075 0.16 0.175 1.26 ;
      RECT  0.075 1.26 0.695 1.35 ;
      RECT  0.605 1.35 0.695 1.57 ;
      RECT  0.075 1.35 0.22 1.63 ;
      RECT  0.605 1.57 1.85 1.66 ;
      RECT  1.005 1.19 1.625 1.28 ;
      RECT  1.53 1.28 1.625 1.39 ;
      RECT  1.53 1.39 2.115 1.42 ;
      RECT  1.53 1.42 3.045 1.48 ;
      RECT  2.015 1.48 3.045 1.51 ;
      RECT  2.94 1.51 3.045 1.63 ;
      RECT  0.785 1.23 0.875 1.37 ;
      RECT  0.785 1.37 1.435 1.48 ;
  END
END SEN_FSDPC1BQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPC1BQ_D_3
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&D&RS)|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPC1BQ_D_3
  CLASS CORE ;
  FOREIGN SEN_FSDPC1BQ_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.44 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.3 6.125 0.49 ;
      RECT  5.46 0.49 6.125 0.5 ;
      RECT  5.46 0.5 6.05 0.595 ;
      RECT  5.95 0.595 6.05 1.1 ;
      RECT  5.95 1.1 6.13 1.11 ;
      RECT  5.35 1.11 6.13 1.29 ;
    END
    ANTENNADIFFAREA 0.392 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.425 1.25 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RS
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.26 0.65 0.465 ;
      RECT  0.405 0.465 0.65 0.555 ;
      RECT  0.55 0.555 0.65 1.01 ;
      RECT  0.55 1.01 1.92 1.1 ;
      RECT  1.75 1.1 1.92 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.37 1.44 0.475 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  2.19 1.58 2.36 1.75 ;
      RECT  3.74 1.495 3.91 1.75 ;
      RECT  4.78 1.4 4.9 1.75 ;
      RECT  5.225 1.415 5.35 1.75 ;
      RECT  5.745 1.38 5.865 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  2.315 0.05 2.485 0.21 ;
      RECT  0.325 0.05 0.445 0.375 ;
      RECT  1.705 0.05 1.825 0.4 ;
      RECT  5.225 0.05 5.345 0.4 ;
      RECT  5.745 0.05 5.86 0.4 ;
      RECT  4.755 0.05 4.925 0.425 ;
      RECT  3.73 0.05 3.85 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.995 0.19 3.11 0.3 ;
      RECT  1.915 0.3 3.11 0.42 ;
      RECT  1.915 0.42 2.005 0.49 ;
      RECT  0.75 0.2 1.59 0.315 ;
      RECT  1.5 0.315 1.59 0.49 ;
      RECT  1.5 0.49 2.005 0.58 ;
      RECT  4.235 0.325 4.62 0.425 ;
      RECT  4.53 0.425 4.62 1.02 ;
      RECT  4.53 1.02 5.04 1.11 ;
      RECT  4.95 0.7 5.04 1.02 ;
      RECT  4.53 1.11 4.62 1.495 ;
      RECT  4.26 1.495 4.62 1.59 ;
      RECT  4.015 0.25 4.105 0.49 ;
      RECT  4.015 0.49 4.17 0.585 ;
      RECT  4.08 0.585 4.17 1.135 ;
      RECT  3.6 0.87 3.69 1.135 ;
      RECT  3.6 1.135 4.17 1.225 ;
      RECT  3.25 0.41 3.385 0.58 ;
      RECT  3.29 0.58 3.385 0.675 ;
      RECT  3.29 0.675 3.975 0.765 ;
      RECT  3.885 0.765 3.975 1.02 ;
      RECT  3.29 0.765 3.38 1.29 ;
      RECT  3.285 1.29 3.38 1.46 ;
      RECT  2.62 0.51 2.72 0.585 ;
      RECT  2.62 0.585 2.97 0.685 ;
      RECT  2.88 0.685 2.97 1.175 ;
      RECT  2.64 1.175 2.97 1.275 ;
      RECT  4.71 0.515 5.245 0.605 ;
      RECT  5.145 0.605 5.245 0.785 ;
      RECT  4.71 0.605 4.8 0.925 ;
      RECT  5.145 0.785 5.84 0.895 ;
      RECT  5.145 0.895 5.245 1.205 ;
      RECT  4.99 1.205 5.245 1.305 ;
      RECT  2.095 0.51 2.53 0.62 ;
      RECT  2.44 0.62 2.53 0.785 ;
      RECT  2.44 0.785 2.77 0.895 ;
      RECT  2.44 0.895 2.53 1.21 ;
      RECT  2.145 1.21 2.53 1.3 ;
      RECT  4.26 0.54 4.44 0.73 ;
      RECT  4.26 0.73 4.35 1.315 ;
      RECT  3.545 1.315 4.35 1.405 ;
      RECT  3.545 1.405 3.635 1.55 ;
      RECT  3.07 0.7 3.195 0.87 ;
      RECT  3.105 0.87 3.195 1.55 ;
      RECT  3.105 1.55 3.635 1.66 ;
      RECT  0.075 0.165 0.175 1.26 ;
      RECT  0.075 1.26 0.655 1.35 ;
      RECT  0.565 1.35 0.655 1.57 ;
      RECT  0.075 1.35 0.22 1.63 ;
      RECT  0.565 1.57 1.81 1.66 ;
      RECT  0.965 1.19 1.585 1.28 ;
      RECT  1.49 1.28 1.585 1.39 ;
      RECT  1.49 1.39 3.015 1.48 ;
      RECT  2.905 1.48 3.015 1.63 ;
      RECT  0.745 1.23 0.85 1.37 ;
      RECT  0.745 1.37 1.395 1.48 ;
  END
END SEN_FSDPC1BQ_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPC1BQ_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&D&RS)|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPC1BQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDPC1BQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.13 0.705 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.415 0.48 6.07 0.595 ;
      RECT  5.95 0.595 6.07 1.11 ;
      RECT  5.435 1.11 6.07 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RS
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.26 0.65 0.46 ;
      RECT  0.405 0.46 0.65 0.56 ;
      RECT  0.55 0.56 0.65 1.01 ;
      RECT  0.55 1.01 1.92 1.1 ;
      RECT  1.75 1.1 1.92 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.365 1.44 0.475 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  2.18 1.6 2.35 1.75 ;
      RECT  3.695 1.495 3.865 1.75 ;
      RECT  4.735 1.4 4.855 1.75 ;
      RECT  5.18 1.4 5.3 1.75 ;
      RECT  5.7 1.38 5.82 1.75 ;
      RECT  6.21 1.41 6.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  2.315 0.05 2.485 0.21 ;
      RECT  0.325 0.05 0.445 0.37 ;
      RECT  5.7 0.05 5.82 0.39 ;
      RECT  6.21 0.05 6.345 0.39 ;
      RECT  5.18 0.05 5.3 0.41 ;
      RECT  1.705 0.05 1.825 0.42 ;
      RECT  4.71 0.05 4.88 0.425 ;
      RECT  3.685 0.05 3.805 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.945 0.19 3.065 0.3 ;
      RECT  1.915 0.3 3.065 0.42 ;
      RECT  1.915 0.42 2.005 0.51 ;
      RECT  0.75 0.21 1.59 0.315 ;
      RECT  1.5 0.315 1.59 0.51 ;
      RECT  1.5 0.51 2.005 0.6 ;
      RECT  3.955 0.25 4.075 0.485 ;
      RECT  3.955 0.485 4.125 0.58 ;
      RECT  4.035 0.58 4.125 1.135 ;
      RECT  3.555 0.855 3.645 1.135 ;
      RECT  3.555 1.135 4.125 1.225 ;
      RECT  3.205 0.41 3.34 0.58 ;
      RECT  3.245 0.58 3.34 0.675 ;
      RECT  3.245 0.675 3.93 0.765 ;
      RECT  3.84 0.765 3.93 1.01 ;
      RECT  3.245 0.765 3.335 1.29 ;
      RECT  3.24 1.29 3.335 1.46 ;
      RECT  2.62 0.51 2.72 0.585 ;
      RECT  2.62 0.585 2.945 0.685 ;
      RECT  2.855 0.685 2.945 1.015 ;
      RECT  2.855 1.015 2.97 1.19 ;
      RECT  2.64 1.19 2.97 1.3 ;
      RECT  4.665 0.515 5.215 0.605 ;
      RECT  5.115 0.605 5.215 0.785 ;
      RECT  4.665 0.605 4.755 0.935 ;
      RECT  5.115 0.785 5.84 0.895 ;
      RECT  5.115 0.895 5.215 1.205 ;
      RECT  4.94 1.205 5.215 1.305 ;
      RECT  2.095 0.51 2.53 0.61 ;
      RECT  2.44 0.61 2.53 0.785 ;
      RECT  2.44 0.785 2.74 0.895 ;
      RECT  2.44 0.895 2.53 1.21 ;
      RECT  2.12 1.21 2.53 1.3 ;
      RECT  4.215 0.54 4.395 0.71 ;
      RECT  4.215 0.71 4.305 1.315 ;
      RECT  3.5 1.315 4.305 1.405 ;
      RECT  3.5 1.405 3.59 1.55 ;
      RECT  3.035 0.7 3.15 0.87 ;
      RECT  3.06 0.87 3.15 1.55 ;
      RECT  3.06 1.55 3.59 1.66 ;
      RECT  4.845 0.75 4.995 0.92 ;
      RECT  4.845 0.92 4.935 1.025 ;
      RECT  4.19 0.325 4.575 0.42 ;
      RECT  4.485 0.42 4.575 1.025 ;
      RECT  4.485 1.025 4.935 1.115 ;
      RECT  4.485 1.115 4.575 1.495 ;
      RECT  4.215 1.495 4.575 1.595 ;
      RECT  0.075 0.165 0.18 1.26 ;
      RECT  0.075 1.26 0.655 1.35 ;
      RECT  0.565 1.35 0.655 1.57 ;
      RECT  0.075 1.35 0.225 1.625 ;
      RECT  0.565 1.57 1.81 1.66 ;
      RECT  0.965 1.19 1.595 1.28 ;
      RECT  1.49 1.28 1.595 1.39 ;
      RECT  1.49 1.39 2.96 1.48 ;
      RECT  2.855 1.48 2.96 1.63 ;
      RECT  0.745 1.23 0.85 1.37 ;
      RECT  0.745 1.37 1.395 1.48 ;
  END
END SEN_FSDPC1BQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPC1BQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&D&RS)|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPC1BQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDPC1BQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.175 0.71 5.275 1.19 ;
      RECT  4.63 0.46 4.73 0.89 ;
      RECT  3.385 0.69 3.485 0.88 ;
      RECT  3.385 0.88 4.155 0.98 ;
      LAYER M2 ;
      RECT  3.345 0.75 5.32 0.85 ;
      LAYER V1 ;
      RECT  5.175 0.75 5.275 0.85 ;
      RECT  4.63 0.75 4.73 0.85 ;
      RECT  3.385 0.75 3.485 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0717 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.86 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.31 6.25 1.16 ;
    END
    ANTENNADIFFAREA 0.166 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RS
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.655 1.85 0.915 ;
      RECT  1.75 0.915 1.93 1.01 ;
      RECT  0.55 0.31 0.65 0.5 ;
      RECT  0.405 0.5 0.65 0.615 ;
      RECT  0.55 0.615 0.65 1.01 ;
      RECT  0.55 1.01 1.93 1.1 ;
      RECT  1.75 1.1 1.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.165 6.47 0.475 ;
      RECT  6.35 0.475 6.745 0.69 ;
      RECT  6.625 0.69 6.745 1.38 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.355 1.44 0.46 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.935 1.57 2.055 1.75 ;
      RECT  3.395 1.465 3.515 1.75 ;
      RECT  4.2 1.43 4.32 1.75 ;
      RECT  5.64 1.48 5.81 1.75 ;
      RECT  6.365 1.43 6.485 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  1.74 0.05 1.86 0.24 ;
      RECT  5.26 0.05 5.43 0.245 ;
      RECT  3.375 0.05 3.495 0.345 ;
      RECT  5.9 0.05 6.005 0.36 ;
      RECT  6.625 0.05 6.745 0.385 ;
      RECT  0.325 0.05 0.445 0.4 ;
      RECT  4.2 0.05 4.32 0.43 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.065 0.195 2.625 0.285 ;
      RECT  2.065 0.285 2.16 0.33 ;
      RECT  2.505 0.285 2.625 0.43 ;
      RECT  0.74 0.205 1.47 0.32 ;
      RECT  1.38 0.32 1.47 0.33 ;
      RECT  1.38 0.33 2.16 0.42 ;
      RECT  2.07 0.42 2.16 1.39 ;
      RECT  0.935 1.2 1.585 1.3 ;
      RECT  1.47 1.3 1.585 1.39 ;
      RECT  1.47 1.39 2.465 1.465 ;
      RECT  1.47 1.465 2.67 1.48 ;
      RECT  2.375 1.48 2.67 1.57 ;
      RECT  5.0 0.2 5.09 0.335 ;
      RECT  5.0 0.335 5.81 0.425 ;
      RECT  5.72 0.425 5.81 0.45 ;
      RECT  5.72 0.45 6.015 0.54 ;
      RECT  5.925 0.54 6.015 1.25 ;
      RECT  5.925 1.25 6.49 1.34 ;
      RECT  6.4 0.78 6.49 1.25 ;
      RECT  5.925 1.34 6.025 1.51 ;
      RECT  4.45 0.18 4.58 0.35 ;
      RECT  4.45 0.35 4.54 0.99 ;
      RECT  4.45 0.99 4.825 1.16 ;
      RECT  4.72 0.18 4.91 0.35 ;
      RECT  4.82 0.35 4.91 0.52 ;
      RECT  4.82 0.52 5.085 0.61 ;
      RECT  4.975 0.61 5.085 1.3 ;
      RECT  4.975 1.3 5.815 1.39 ;
      RECT  5.725 0.725 5.815 1.3 ;
      RECT  3.675 0.19 3.775 0.435 ;
      RECT  3.205 0.435 3.775 0.525 ;
      RECT  3.205 0.525 3.295 0.77 ;
      RECT  2.995 0.77 3.295 0.94 ;
      RECT  3.205 0.94 3.295 1.105 ;
      RECT  3.205 1.105 3.815 1.195 ;
      RECT  5.24 0.515 5.63 0.615 ;
      RECT  5.525 0.615 5.63 1.165 ;
      RECT  3.89 0.535 4.355 0.655 ;
      RECT  3.89 0.655 3.98 0.69 ;
      RECT  4.265 0.655 4.355 1.245 ;
      RECT  3.575 0.69 3.98 0.79 ;
      RECT  3.925 1.165 4.025 1.245 ;
      RECT  3.925 1.245 4.355 1.25 ;
      RECT  3.925 1.25 4.695 1.34 ;
      RECT  4.605 1.34 4.695 1.66 ;
      RECT  2.78 0.42 2.87 0.685 ;
      RECT  2.43 0.685 2.87 0.855 ;
      RECT  2.735 0.855 2.87 1.06 ;
      RECT  2.735 1.06 2.925 1.18 ;
      RECT  2.25 0.385 2.34 1.14 ;
      RECT  2.25 1.14 2.645 1.23 ;
      RECT  2.555 1.23 2.645 1.285 ;
      RECT  2.555 1.285 3.8 1.375 ;
      RECT  3.71 1.375 3.8 1.495 ;
      RECT  3.185 1.375 3.285 1.59 ;
      RECT  3.71 1.495 3.985 1.66 ;
      RECT  0.07 0.18 0.18 1.26 ;
      RECT  0.07 1.26 0.64 1.35 ;
      RECT  0.55 1.35 0.64 1.57 ;
      RECT  0.07 1.35 0.21 1.61 ;
      RECT  0.55 1.57 1.745 1.66 ;
      RECT  0.73 1.22 0.82 1.39 ;
      RECT  0.73 1.39 1.38 1.48 ;
      RECT  4.785 1.29 4.885 1.48 ;
      RECT  4.785 1.48 5.42 1.595 ;
      LAYER M2 ;
      RECT  4.745 1.35 6.1 1.45 ;
      LAYER V1 ;
      RECT  4.785 1.35 4.885 1.45 ;
      RECT  5.925 1.35 6.025 1.45 ;
  END
END SEN_FSDPC1BQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPC1BQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&D&RS)|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPC1BQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDPC1BQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.535 0.51 6.65 1.115 ;
      RECT  5.98 0.55 6.08 0.785 ;
      RECT  5.8 0.785 6.08 0.89 ;
      RECT  4.705 0.59 4.84 0.915 ;
      LAYER M2 ;
      RECT  4.7 0.75 6.675 0.85 ;
      LAYER V1 ;
      RECT  6.535 0.75 6.635 0.85 ;
      RECT  5.98 0.75 6.08 0.85 ;
      RECT  4.74 0.75 4.84 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.4 ;
      RECT  0.35 0.4 0.65 0.49 ;
      RECT  0.55 0.49 0.65 0.945 ;
      RECT  0.55 0.945 0.98 1.045 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0846 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.495 0.195 7.65 0.365 ;
      RECT  7.55 0.365 7.65 0.99 ;
      RECT  7.51 0.99 7.65 1.165 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.285 0.745 1.59 0.975 ;
      LAYER M2 ;
      RECT  1.31 0.75 1.88 0.85 ;
      LAYER V1 ;
      RECT  1.42 0.75 1.52 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0846 ;
  END RS
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.665 0.555 2.765 1.13 ;
      RECT  0.35 0.58 0.45 1.045 ;
      LAYER M2 ;
      RECT  0.31 0.75 0.65 0.85 ;
      RECT  0.55 0.85 0.65 0.95 ;
      RECT  0.55 0.95 2.805 1.05 ;
      LAYER V1 ;
      RECT  2.665 0.95 2.765 1.05 ;
      RECT  0.35 0.75 0.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.087 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.135 ;
      RECT  0.15 1.135 2.345 1.225 ;
      RECT  2.255 1.055 2.345 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.29 8.145 0.51 ;
      RECT  8.055 0.51 8.145 1.11 ;
      RECT  7.95 1.11 8.145 1.37 ;
      RECT  7.95 1.37 8.05 1.49 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.56 1.495 0.73 1.75 ;
      RECT  2.34 1.495 2.51 1.75 ;
      RECT  2.73 1.495 2.9 1.75 ;
      RECT  4.265 1.365 4.435 1.75 ;
      RECT  5.045 1.39 5.215 1.75 ;
      RECT  5.575 1.61 5.745 1.75 ;
      RECT  6.88 1.44 7.0 1.75 ;
      RECT  7.235 1.44 7.355 1.75 ;
      RECT  7.745 1.435 7.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  6.695 0.05 6.865 0.2 ;
      RECT  7.155 0.05 7.325 0.2 ;
      RECT  1.895 0.05 2.015 0.23 ;
      RECT  2.74 0.05 2.87 0.23 ;
      RECT  4.525 0.05 4.695 0.32 ;
      RECT  5.56 0.05 5.68 0.375 ;
      RECT  0.11 0.05 0.25 0.39 ;
      RECT  4.06 0.05 4.18 0.405 ;
      RECT  5.07 0.05 5.19 0.435 ;
      RECT  7.755 0.05 7.86 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.565 0.14 1.705 0.23 ;
      RECT  0.565 0.23 0.735 0.31 ;
      RECT  1.615 0.23 1.705 0.32 ;
      RECT  1.615 0.32 3.49 0.41 ;
      RECT  2.875 0.41 3.49 0.425 ;
      RECT  2.875 0.425 2.965 1.315 ;
      RECT  1.98 1.315 3.08 1.405 ;
      RECT  2.99 1.405 3.08 1.44 ;
      RECT  1.98 1.405 2.08 1.495 ;
      RECT  2.99 1.44 3.675 1.53 ;
      RECT  3.505 1.425 3.675 1.44 ;
      RECT  0.84 1.495 2.08 1.6 ;
      RECT  5.795 0.225 5.94 0.395 ;
      RECT  5.795 0.395 5.885 0.465 ;
      RECT  5.275 0.465 5.885 0.555 ;
      RECT  5.275 0.555 5.595 0.585 ;
      RECT  5.505 0.585 5.595 1.0 ;
      RECT  5.285 1.0 6.235 1.12 ;
      RECT  6.08 0.225 6.26 0.395 ;
      RECT  6.17 0.395 6.26 0.47 ;
      RECT  6.17 0.47 6.44 0.56 ;
      RECT  6.34 0.56 6.44 1.22 ;
      RECT  5.78 1.22 6.44 1.25 ;
      RECT  5.78 1.25 6.455 1.34 ;
      RECT  6.365 1.34 6.455 1.42 ;
      RECT  0.855 0.32 1.525 0.41 ;
      RECT  0.855 0.41 0.965 0.84 ;
      RECT  4.81 0.28 4.93 0.41 ;
      RECT  4.525 0.41 4.93 0.5 ;
      RECT  4.525 0.5 4.615 0.72 ;
      RECT  4.46 0.72 4.615 1.005 ;
      RECT  4.46 1.005 4.835 1.095 ;
      RECT  4.745 1.095 4.835 1.21 ;
      RECT  4.745 1.21 5.495 1.3 ;
      RECT  5.405 1.3 5.495 1.43 ;
      RECT  5.405 1.43 6.075 1.52 ;
      RECT  5.975 1.52 6.075 1.545 ;
      RECT  5.975 1.545 6.265 1.655 ;
      RECT  4.32 0.3 4.435 0.495 ;
      RECT  3.8 0.495 4.435 0.585 ;
      RECT  3.8 0.585 3.89 0.895 ;
      RECT  3.67 0.895 3.89 0.985 ;
      RECT  3.8 0.985 3.89 1.065 ;
      RECT  3.8 1.065 4.075 1.155 ;
      RECT  3.985 1.155 4.075 1.185 ;
      RECT  3.985 1.185 4.655 1.275 ;
      RECT  4.55 1.275 4.655 1.48 ;
      RECT  3.59 0.425 3.71 0.555 ;
      RECT  3.245 0.555 3.71 0.645 ;
      RECT  3.245 0.645 3.355 1.245 ;
      RECT  3.245 1.245 3.895 1.335 ;
      RECT  3.245 1.335 3.415 1.35 ;
      RECT  3.805 1.335 3.895 1.415 ;
      RECT  1.065 0.5 2.35 0.59 ;
      RECT  6.94 0.515 7.14 0.615 ;
      RECT  6.94 0.615 7.04 0.76 ;
      RECT  6.74 0.76 7.04 0.945 ;
      RECT  6.94 0.945 7.04 1.16 ;
      RECT  2.47 0.505 2.575 0.845 ;
      RECT  1.86 0.845 2.575 0.945 ;
      RECT  2.47 0.945 2.575 1.16 ;
      RECT  4.93 0.75 5.4 0.86 ;
      RECT  4.93 0.86 5.03 1.095 ;
      RECT  7.875 0.74 7.965 0.86 ;
      RECT  7.755 0.86 7.965 0.95 ;
      RECT  7.755 0.95 7.845 1.255 ;
      RECT  6.37 0.17 6.49 0.29 ;
      RECT  6.37 0.29 7.36 0.38 ;
      RECT  7.27 0.38 7.36 0.455 ;
      RECT  7.27 0.455 7.42 0.545 ;
      RECT  7.33 0.545 7.42 1.255 ;
      RECT  6.62 1.255 7.845 1.345 ;
      RECT  6.62 1.345 6.74 1.61 ;
      RECT  3.98 0.675 4.07 0.885 ;
      RECT  3.98 0.885 4.265 0.975 ;
      RECT  4.165 0.975 4.265 1.095 ;
      RECT  7.14 0.71 7.24 1.16 ;
      RECT  3.055 0.52 3.155 1.17 ;
      RECT  0.325 1.315 1.82 1.405 ;
      RECT  0.325 1.405 0.445 1.545 ;
      LAYER M2 ;
      RECT  3.015 0.95 5.07 1.05 ;
      RECT  6.3 0.95 7.28 1.05 ;
      LAYER V1 ;
      RECT  3.055 0.95 3.155 1.05 ;
      RECT  4.165 0.95 4.265 1.05 ;
      RECT  4.93 0.95 5.03 1.05 ;
      RECT  6.34 0.95 6.44 1.05 ;
      RECT  7.14 0.95 7.24 1.05 ;
  END
END SEN_FSDPC1BQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPC1BQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-sync-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&D&RS)|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPC1BQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDPC1BQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.42 0.69 7.52 0.905 ;
      RECT  7.42 0.905 7.705 0.995 ;
      RECT  7.605 0.995 7.705 1.165 ;
      RECT  6.0 0.58 6.875 0.67 ;
      RECT  6.0 0.67 6.095 0.71 ;
      RECT  6.77 0.67 6.875 0.89 ;
      RECT  5.62 0.71 6.095 0.89 ;
      LAYER M2 ;
      RECT  6.73 0.75 7.56 0.85 ;
      LAYER V1 ;
      RECT  7.42 0.75 7.52 0.85 ;
      RECT  6.77 0.75 6.87 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.117 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1092 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 0.475 9.25 0.595 ;
      RECT  9.15 0.595 9.25 1.025 ;
      RECT  8.52 1.025 9.25 1.145 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.83 ;
      RECT  1.15 0.83 1.81 0.94 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1092 ;
  END RS
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.88 0.51 2.98 1.11 ;
      RECT  0.35 0.51 0.45 0.95 ;
      RECT  0.35 0.95 0.53 1.05 ;
      LAYER M2 ;
      RECT  0.35 0.95 3.02 1.05 ;
      LAYER V1 ;
      RECT  2.88 0.95 2.98 1.05 ;
      RECT  0.39 0.95 0.49 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1035 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.14 ;
      RECT  0.15 1.14 2.465 1.205 ;
      RECT  0.6 1.115 2.465 1.14 ;
      RECT  0.15 1.205 0.665 1.23 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.55 0.31 9.745 0.49 ;
      RECT  9.655 0.49 9.745 1.11 ;
      RECT  9.55 1.11 9.745 1.49 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.37 0.185 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  0.61 1.52 0.73 1.75 ;
      RECT  2.33 1.475 2.5 1.75 ;
      RECT  2.93 1.475 3.1 1.75 ;
      RECT  3.47 1.48 3.64 1.75 ;
      RECT  4.89 1.365 5.01 1.75 ;
      RECT  5.83 1.39 5.95 1.75 ;
      RECT  6.335 1.585 6.505 1.75 ;
      RECT  7.965 1.44 8.085 1.75 ;
      RECT  8.315 1.44 8.435 1.75 ;
      RECT  8.835 1.44 8.955 1.75 ;
      RECT  9.345 1.44 9.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  2.14 0.05 2.31 0.19 ;
      RECT  2.94 0.05 3.11 0.19 ;
      RECT  3.48 0.05 3.65 0.19 ;
      RECT  7.68 0.05 7.85 0.21 ;
      RECT  6.325 0.05 6.495 0.31 ;
      RECT  8.835 0.05 8.955 0.385 ;
      RECT  0.095 0.05 0.235 0.39 ;
      RECT  5.31 0.05 5.43 0.39 ;
      RECT  8.315 0.05 8.435 0.4 ;
      RECT  5.83 0.05 5.95 0.405 ;
      RECT  9.355 0.05 9.46 0.405 ;
      RECT  4.8 0.05 4.92 0.43 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.56 0.14 2.03 0.23 ;
      RECT  1.94 0.23 2.03 0.28 ;
      RECT  0.56 0.23 0.73 0.385 ;
      RECT  1.94 0.28 4.2 0.37 ;
      RECT  3.07 0.37 4.2 0.42 ;
      RECT  3.07 0.42 3.16 1.295 ;
      RECT  1.97 1.295 4.24 1.385 ;
      RECT  1.97 1.385 2.07 1.495 ;
      RECT  0.83 1.495 2.07 1.59 ;
      RECT  6.82 0.21 7.33 0.31 ;
      RECT  7.23 0.31 7.33 1.085 ;
      RECT  7.23 1.085 7.485 1.175 ;
      RECT  7.385 1.175 7.485 1.44 ;
      RECT  7.385 1.44 7.6 1.455 ;
      RECT  6.865 1.455 7.6 1.56 ;
      RECT  0.82 0.32 1.81 0.41 ;
      RECT  6.065 0.4 7.14 0.49 ;
      RECT  7.05 0.49 7.14 1.265 ;
      RECT  6.645 1.265 7.295 1.365 ;
      RECT  6.645 1.365 6.75 1.395 ;
      RECT  6.065 1.395 6.75 1.495 ;
      RECT  4.315 0.4 4.42 0.52 ;
      RECT  3.72 0.52 4.42 0.62 ;
      RECT  3.72 0.62 3.81 0.785 ;
      RECT  3.46 0.785 3.81 0.895 ;
      RECT  3.72 0.895 3.81 1.115 ;
      RECT  3.72 1.115 4.47 1.205 ;
      RECT  5.06 0.37 5.18 0.52 ;
      RECT  4.56 0.52 5.18 0.61 ;
      RECT  4.56 0.61 4.65 0.715 ;
      RECT  4.34 0.715 4.65 0.81 ;
      RECT  4.56 0.81 4.65 1.185 ;
      RECT  4.56 1.185 5.265 1.275 ;
      RECT  5.175 1.275 5.265 1.435 ;
      RECT  2.06 0.465 2.58 0.555 ;
      RECT  2.06 0.555 2.15 0.56 ;
      RECT  1.35 0.56 2.15 0.65 ;
      RECT  7.88 0.48 7.985 0.665 ;
      RECT  7.61 0.665 7.985 0.765 ;
      RECT  7.87 0.765 7.985 0.92 ;
      RECT  7.87 0.92 8.08 1.01 ;
      RECT  7.975 1.01 8.08 1.17 ;
      RECT  2.7 0.52 2.79 0.78 ;
      RECT  2.575 0.78 2.79 0.85 ;
      RECT  2.13 0.85 2.79 0.89 ;
      RECT  2.13 0.89 2.665 0.96 ;
      RECT  2.575 0.96 2.665 1.185 ;
      RECT  8.35 0.51 8.45 0.785 ;
      RECT  8.35 0.785 9.045 0.895 ;
      RECT  9.465 0.74 9.565 0.88 ;
      RECT  9.35 0.88 9.565 0.97 ;
      RECT  9.35 0.97 9.44 1.26 ;
      RECT  7.42 0.17 7.525 0.3 ;
      RECT  7.42 0.3 8.165 0.39 ;
      RECT  8.075 0.39 8.165 0.74 ;
      RECT  8.075 0.74 8.26 0.83 ;
      RECT  8.17 0.83 8.26 1.26 ;
      RECT  7.71 1.26 9.44 1.35 ;
      RECT  7.71 1.35 7.82 1.59 ;
      RECT  6.185 0.78 6.57 0.9 ;
      RECT  6.185 0.9 6.365 1.055 ;
      RECT  4.74 0.715 4.84 1.005 ;
      RECT  4.74 1.005 5.18 1.095 ;
      RECT  6.465 1.01 6.96 1.12 ;
      RECT  6.465 1.12 6.555 1.185 ;
      RECT  5.425 0.48 5.74 0.6 ;
      RECT  5.425 0.6 5.515 0.815 ;
      RECT  4.97 0.815 5.515 0.915 ;
      RECT  5.425 0.915 5.515 1.185 ;
      RECT  5.425 1.185 6.555 1.275 ;
      RECT  3.25 0.52 3.35 1.175 ;
      RECT  0.7 1.315 1.81 1.34 ;
      RECT  0.3 1.34 1.81 1.405 ;
      RECT  0.3 1.405 0.765 1.43 ;
      LAYER M2 ;
      RECT  7.19 0.55 8.49 0.65 ;
      RECT  3.21 0.95 6.365 1.05 ;
      LAYER V1 ;
      RECT  7.23 0.55 7.33 0.65 ;
      RECT  8.35 0.55 8.45 0.65 ;
      RECT  3.25 0.95 3.35 1.05 ;
      RECT  4.74 0.95 4.84 1.05 ;
      RECT  6.225 0.95 6.325 1.05 ;
  END
END SEN_FSDPC1BQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPHQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, sync hold, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(iq&EN&!SE)|(!EN&(!SE&D))|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPHQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPHQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.05 1.21 ;
      RECT  4.95 1.21 5.38 1.3 ;
      RECT  5.29 1.3 5.38 1.52 ;
      RECT  5.29 1.52 5.83 1.625 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1176 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.07 0.75 1.17 1.27 ;
      LAYER M2 ;
      RECT  0.655 0.95 1.21 1.05 ;
      LAYER V1 ;
      RECT  1.07 0.95 1.17 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.26 0.75 1.465 0.77 ;
      RECT  1.26 0.77 2.17 0.86 ;
      RECT  0.3 0.51 0.45 0.71 ;
      RECT  0.3 0.71 0.61 0.89 ;
      LAYER M2 ;
      RECT  0.47 0.75 1.44 0.85 ;
      LAYER V1 ;
      RECT  1.3 0.75 1.4 0.85 ;
      RECT  0.51 0.75 0.61 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0927 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.31 6.86 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.165 0.19 3.265 0.71 ;
      RECT  0.7 0.495 0.8 0.985 ;
      LAYER M2 ;
      RECT  0.66 0.55 3.305 0.65 ;
      LAYER V1 ;
      RECT  3.165 0.55 3.265 0.65 ;
      RECT  0.7 0.55 0.8 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.335 0.98 0.505 1.49 ;
      LAYER M2 ;
      RECT  0.365 1.35 1.02 1.45 ;
      LAYER V1 ;
      RECT  0.405 1.35 0.505 1.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.585 0.485 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  3.015 1.59 3.185 1.75 ;
      RECT  3.64 1.59 3.81 1.75 ;
      RECT  4.93 1.39 5.1 1.75 ;
      RECT  5.99 1.49 6.115 1.75 ;
      RECT  6.495 1.385 6.615 1.75 ;
      RECT  7.015 1.21 7.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  0.35 0.05 0.465 0.24 ;
      RECT  5.995 0.05 6.115 0.38 ;
      RECT  6.495 0.05 6.615 0.38 ;
      RECT  3.66 0.05 3.785 0.4 ;
      RECT  7.015 0.05 7.135 0.59 ;
      RECT  2.7 0.05 2.82 0.61 ;
      RECT  4.945 0.05 5.065 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.555 0.15 2.45 0.25 ;
      RECT  0.555 0.25 0.645 0.33 ;
      RECT  0.065 0.33 0.645 0.42 ;
      RECT  0.065 0.42 0.185 1.56 ;
      RECT  4.57 0.14 4.805 0.31 ;
      RECT  4.685 0.31 4.805 1.57 ;
      RECT  3.95 1.57 4.805 1.66 ;
      RECT  5.66 0.22 5.885 0.34 ;
      RECT  5.66 0.34 5.76 1.03 ;
      RECT  5.66 1.03 5.845 1.22 ;
      RECT  5.155 0.225 5.35 0.345 ;
      RECT  5.25 0.345 5.35 0.99 ;
      RECT  5.155 0.99 5.35 1.12 ;
      RECT  1.605 0.34 2.56 0.46 ;
      RECT  2.45 0.46 2.56 0.59 ;
      RECT  3.95 0.29 4.05 0.52 ;
      RECT  3.36 0.52 4.05 0.62 ;
      RECT  3.36 0.62 3.45 1.095 ;
      RECT  3.36 1.095 3.515 1.265 ;
      RECT  5.865 0.47 6.62 0.575 ;
      RECT  6.52 0.575 6.62 0.855 ;
      RECT  5.865 0.575 5.955 0.86 ;
      RECT  6.28 0.855 6.62 0.96 ;
      RECT  6.28 0.96 6.385 1.245 ;
      RECT  4.18 0.28 4.29 0.755 ;
      RECT  3.555 0.755 4.29 0.855 ;
      RECT  3.555 0.855 3.665 0.985 ;
      RECT  4.175 0.855 4.29 1.26 ;
      RECT  2.6 0.71 2.71 0.85 ;
      RECT  2.6 0.85 3.27 0.94 ;
      RECT  2.975 0.47 3.075 0.85 ;
      RECT  3.17 0.94 3.27 1.29 ;
      RECT  1.535 0.95 2.165 1.05 ;
      RECT  5.47 0.19 5.57 1.31 ;
      RECT  5.47 1.31 6.19 1.4 ;
      RECT  6.1 0.665 6.19 1.31 ;
      RECT  4.435 0.4 4.555 1.355 ;
      RECT  3.6 1.355 4.555 1.41 ;
      RECT  0.89 0.495 0.98 0.555 ;
      RECT  0.89 0.555 2.36 0.645 ;
      RECT  2.27 0.645 2.36 1.135 ;
      RECT  0.89 0.645 0.98 1.185 ;
      RECT  2.27 1.135 3.035 1.225 ;
      RECT  2.945 1.225 3.035 1.41 ;
      RECT  2.945 1.41 4.555 1.445 ;
      RECT  2.945 1.445 3.705 1.5 ;
      RECT  1.39 1.315 2.85 1.405 ;
      RECT  1.39 1.405 1.51 1.61 ;
      RECT  1.6 1.495 2.34 1.6 ;
      RECT  0.7 1.08 0.8 1.635 ;
      LAYER M2 ;
      RECT  3.91 0.35 5.39 0.45 ;
      RECT  1.71 0.95 5.8 1.05 ;
      RECT  0.66 1.15 3.31 1.25 ;
      LAYER V1 ;
      RECT  3.95 0.35 4.05 0.45 ;
      RECT  5.25 0.35 5.35 0.45 ;
      RECT  1.75 0.95 1.85 1.05 ;
      RECT  5.66 0.95 5.76 1.05 ;
      RECT  0.7 1.15 0.8 1.25 ;
      RECT  3.17 1.15 3.27 1.25 ;
  END
END SEN_FSDPHQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPHQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, sync hold, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(iq&EN&!SE)|(!EN&(!SE&D))|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPHQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDPHQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.25 0.71 7.35 0.795 ;
      RECT  7.25 0.795 7.45 0.885 ;
      RECT  7.25 0.885 7.35 1.085 ;
      RECT  6.75 0.69 6.895 1.2 ;
      LAYER M2 ;
      RECT  6.71 0.75 7.39 0.85 ;
      LAYER V1 ;
      RECT  7.25 0.75 7.35 0.85 ;
      RECT  6.75 0.75 6.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1059 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.825 0.71 4.105 0.895 ;
      LAYER M2 ;
      RECT  2.84 0.75 4.025 0.85 ;
      LAYER V1 ;
      RECT  3.885 0.75 3.985 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END EN
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.75 0.31 9.87 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.025 0.945 1.125 1.11 ;
      RECT  1.025 1.11 1.65 1.29 ;
      RECT  1.52 0.87 1.65 1.11 ;
      RECT  1.55 1.29 1.65 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1002 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.325 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.275 0.27 9.38 0.42 ;
      RECT  9.275 0.42 9.45 0.495 ;
      RECT  9.33 0.495 9.45 1.355 ;
    END
    ANTENNADIFFAREA 0.105 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.405 0.455 1.75 ;
      RECT  0.0 1.75 10.2 1.85 ;
      RECT  1.35 1.415 1.46 1.75 ;
      RECT  2.355 1.605 2.525 1.75 ;
      RECT  2.89 1.44 3.01 1.75 ;
      RECT  4.755 1.425 4.875 1.75 ;
      RECT  5.865 1.48 6.035 1.75 ;
      RECT  6.635 1.48 6.805 1.75 ;
      RECT  7.775 1.525 7.945 1.75 ;
      RECT  8.27 1.58 8.44 1.75 ;
      RECT  9.04 1.415 9.16 1.75 ;
      RECT  9.48 1.45 9.65 1.75 ;
      RECT  10.015 1.41 10.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      RECT  4.35 0.05 4.52 0.185 ;
      RECT  8.175 0.05 8.345 0.185 ;
      RECT  7.66 0.05 7.78 0.26 ;
      RECT  1.825 0.05 1.995 0.305 ;
      RECT  2.355 0.05 2.525 0.305 ;
      RECT  5.485 0.05 5.655 0.305 ;
      RECT  6.28 0.05 6.45 0.305 ;
      RECT  8.99 0.05 9.145 0.36 ;
      RECT  9.52 0.05 9.625 0.36 ;
      RECT  10.015 0.05 10.145 0.39 ;
      RECT  1.31 0.05 1.43 0.42 ;
      RECT  0.31 0.05 0.48 0.44 ;
      RECT  3.26 0.05 3.385 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.655 0.14 1.11 0.255 ;
      RECT  0.655 0.255 0.755 1.525 ;
      RECT  0.655 1.525 0.885 1.635 ;
      RECT  3.765 0.2 4.25 0.275 ;
      RECT  3.765 0.275 4.855 0.32 ;
      RECT  4.155 0.32 4.855 0.365 ;
      RECT  4.605 0.365 4.855 0.395 ;
      RECT  4.605 0.395 4.695 1.245 ;
      RECT  4.48 1.245 5.11 1.295 ;
      RECT  3.395 1.295 5.11 1.335 ;
      RECT  3.395 1.335 4.565 1.39 ;
      RECT  4.985 1.335 5.11 1.465 ;
      RECT  4.21 1.39 4.38 1.405 ;
      RECT  6.57 0.23 6.79 0.35 ;
      RECT  6.57 0.35 6.66 0.395 ;
      RECT  5.24 0.22 5.36 0.395 ;
      RECT  5.24 0.395 6.66 0.485 ;
      RECT  6.57 0.485 6.66 1.3 ;
      RECT  5.615 1.3 7.07 1.39 ;
      RECT  5.615 1.39 5.735 1.61 ;
      RECT  6.15 1.39 6.265 1.62 ;
      RECT  8.675 0.23 8.9 0.35 ;
      RECT  8.81 0.35 8.9 1.395 ;
      RECT  7.605 1.345 8.125 1.395 ;
      RECT  7.605 1.395 8.9 1.435 ;
      RECT  8.035 1.435 8.9 1.485 ;
      RECT  8.755 1.485 8.9 1.62 ;
      RECT  4.945 0.235 5.15 0.355 ;
      RECT  5.055 0.355 5.15 0.6 ;
      RECT  5.055 0.6 5.915 0.69 ;
      RECT  5.82 0.69 5.915 0.78 ;
      RECT  5.055 0.69 5.145 1.065 ;
      RECT  5.82 0.78 6.25 0.89 ;
      RECT  5.055 1.065 5.29 1.155 ;
      RECT  5.2 1.155 5.29 1.465 ;
      RECT  5.2 1.465 5.46 1.585 ;
      RECT  7.235 0.305 7.51 0.425 ;
      RECT  7.42 0.425 7.51 0.55 ;
      RECT  7.42 0.55 7.64 0.65 ;
      RECT  7.54 0.65 7.64 0.98 ;
      RECT  7.44 0.98 7.64 1.07 ;
      RECT  0.845 0.35 1.025 0.45 ;
      RECT  0.845 0.45 0.935 1.41 ;
      RECT  2.91 0.35 3.155 0.45 ;
      RECT  3.04 0.45 3.155 0.67 ;
      RECT  7.62 0.35 7.82 0.45 ;
      RECT  7.73 0.45 7.82 1.16 ;
      RECT  7.425 1.16 7.82 1.25 ;
      RECT  7.425 1.25 7.515 1.44 ;
      RECT  7.145 1.44 7.515 1.555 ;
      RECT  6.9 0.2 7.05 0.49 ;
      RECT  8.47 0.2 8.585 0.49 ;
      RECT  8.47 0.49 8.72 0.58 ;
      RECT  8.62 0.58 8.72 1.29 ;
      RECT  0.065 0.295 0.19 0.53 ;
      RECT  0.065 0.53 0.555 0.62 ;
      RECT  0.465 0.62 0.555 1.21 ;
      RECT  0.065 1.21 0.555 1.3 ;
      RECT  0.065 1.3 0.185 1.435 ;
      RECT  3.645 0.455 4.515 0.545 ;
      RECT  3.645 0.545 3.735 0.85 ;
      RECT  4.425 0.545 4.515 0.95 ;
      RECT  2.665 0.425 2.77 0.85 ;
      RECT  2.665 0.85 3.735 0.94 ;
      RECT  2.665 0.94 2.78 1.17 ;
      RECT  9.02 0.45 9.12 0.55 ;
      RECT  9.02 0.55 9.2 0.645 ;
      RECT  9.02 0.645 9.24 0.745 ;
      RECT  1.405 0.51 1.505 0.62 ;
      RECT  1.21 0.62 1.505 0.78 ;
      RECT  1.21 0.78 1.3 0.91 ;
      RECT  6.005 0.575 6.45 0.665 ;
      RECT  6.36 0.665 6.45 1.01 ;
      RECT  5.79 1.01 6.45 1.11 ;
      RECT  6.36 1.11 6.45 1.18 ;
      RECT  5.235 0.81 5.48 0.92 ;
      RECT  5.38 0.92 5.48 1.315 ;
      RECT  8.25 0.31 8.35 0.95 ;
      RECT  8.17 0.95 8.35 1.05 ;
      RECT  4.195 0.71 4.29 1.035 ;
      RECT  3.215 1.035 4.29 1.135 ;
      RECT  3.215 1.135 3.305 1.26 ;
      RECT  1.595 0.42 2.575 0.51 ;
      RECT  1.595 0.51 1.685 0.64 ;
      RECT  2.485 0.51 2.575 1.26 ;
      RECT  2.485 1.26 3.305 1.35 ;
      RECT  2.485 1.35 2.575 1.415 ;
      RECT  1.83 1.415 2.575 1.515 ;
      RECT  4.835 0.535 4.935 1.11 ;
      RECT  7.04 0.585 7.14 1.11 ;
      RECT  9.55 0.51 9.655 1.11 ;
      RECT  7.93 0.25 8.035 1.165 ;
      RECT  7.93 1.165 8.53 1.255 ;
      RECT  8.44 0.67 8.53 1.165 ;
      RECT  5.57 0.8 5.695 1.19 ;
      RECT  2.105 0.6 2.22 1.255 ;
      RECT  8.99 0.855 9.09 1.32 ;
      RECT  3.13 1.445 3.3 1.48 ;
      RECT  3.13 1.48 3.81 1.595 ;
      RECT  3.69 1.595 3.81 1.66 ;
      RECT  3.95 1.48 4.12 1.52 ;
      RECT  3.95 1.52 4.64 1.635 ;
      RECT  4.47 1.48 4.64 1.52 ;
      LAYER M2 ;
      RECT  0.845 0.35 3.09 0.45 ;
      RECT  6.91 0.35 8.39 0.45 ;
      RECT  1.365 0.55 9.21 0.65 ;
      RECT  0.615 0.95 2.255 1.05 ;
      RECT  4.795 0.95 8.07 1.05 ;
      RECT  8.17 0.95 9.69 1.05 ;
      RECT  5.34 1.15 8.76 1.25 ;
      LAYER V1 ;
      RECT  0.885 0.35 0.985 0.45 ;
      RECT  2.95 0.35 3.05 0.45 ;
      RECT  6.95 0.35 7.05 0.45 ;
      RECT  7.66 0.35 7.76 0.45 ;
      RECT  8.25 0.35 8.35 0.45 ;
      RECT  1.405 0.55 1.505 0.65 ;
      RECT  7.46 0.55 7.56 0.65 ;
      RECT  9.06 0.55 9.16 0.65 ;
      RECT  0.655 0.95 0.755 1.05 ;
      RECT  2.115 0.95 2.215 1.05 ;
      RECT  4.835 0.95 4.935 1.05 ;
      RECT  5.57 0.95 5.67 1.05 ;
      RECT  7.04 0.95 7.14 1.05 ;
      RECT  7.93 0.95 8.03 1.05 ;
      RECT  8.21 0.95 8.31 1.05 ;
      RECT  8.99 0.95 9.09 1.05 ;
      RECT  9.55 0.95 9.65 1.05 ;
      RECT  5.38 1.15 5.48 1.25 ;
      RECT  8.62 1.15 8.72 1.25 ;
  END
END SEN_FSDPHQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPMQ_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, 2-to-1 muxed data inputs, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D1&S&!SE)|(!S&(!SE&D0))|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPMQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDPMQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 4.85 1.25 ;
      RECT  4.75 1.25 5.105 1.34 ;
      RECT  5.01 1.34 5.105 1.55 ;
      RECT  5.01 1.55 5.5 1.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 ;
  END CK
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.075 0.71 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.105 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.51 6.545 0.685 ;
      RECT  6.35 0.685 6.45 1.015 ;
      RECT  6.35 1.015 6.545 1.185 ;
    END
    ANTENNADIFFAREA 0.139 ;
  END Q
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.64 ;
      RECT  0.27 0.64 0.45 0.82 ;
      RECT  1.11 0.35 1.45 0.45 ;
      RECT  1.34 0.45 1.45 0.71 ;
      RECT  1.34 0.71 1.86 0.89 ;
      LAYER M2 ;
      RECT  0.445 0.35 1.29 0.45 ;
      RECT  0.445 0.45 0.555 0.55 ;
      RECT  0.31 0.55 0.555 0.65 ;
      LAYER V1 ;
      RECT  0.35 0.55 0.45 0.65 ;
      RECT  1.15 0.35 1.25 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 ;
  END S
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.695 0.485 0.795 1.015 ;
      RECT  2.8 0.15 2.975 0.25 ;
      RECT  2.865 0.25 2.975 0.35 ;
      RECT  2.865 0.35 3.055 0.45 ;
      LAYER M2 ;
      RECT  1.41 0.35 3.055 0.45 ;
      RECT  1.41 0.45 1.51 0.55 ;
      RECT  0.655 0.55 1.51 0.65 ;
      LAYER V1 ;
      RECT  0.695 0.55 0.795 0.65 ;
      RECT  2.915 0.35 3.015 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.91 0.575 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  5.67 1.105 5.87 1.225 ;
      RECT  5.77 1.225 5.87 1.315 ;
      RECT  5.77 1.315 6.285 1.425 ;
      RECT  6.165 1.425 6.285 1.75 ;
      RECT  4.66 1.43 4.91 1.545 ;
      RECT  4.82 1.545 4.91 1.75 ;
      RECT  0.335 1.4 0.455 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  2.85 1.525 2.99 1.75 ;
      RECT  3.475 1.54 3.615 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.345 0.05 0.45 0.225 ;
      RECT  6.165 0.05 6.285 0.39 ;
      RECT  3.485 0.05 3.605 0.43 ;
      RECT  5.72 0.05 5.84 0.485 ;
      RECT  2.58 0.05 2.7 0.61 ;
      RECT  4.745 0.05 4.855 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.54 0.14 1.435 0.24 ;
      RECT  0.54 0.24 0.63 0.315 ;
      RECT  0.075 0.315 0.63 0.405 ;
      RECT  0.075 0.405 0.195 0.515 ;
      RECT  0.075 0.515 0.18 1.37 ;
      RECT  0.075 1.37 0.195 1.61 ;
      RECT  4.37 0.145 4.595 0.315 ;
      RECT  4.475 0.315 4.595 0.565 ;
      RECT  4.42 0.565 4.595 0.67 ;
      RECT  4.42 0.67 4.54 1.165 ;
      RECT  4.45 1.165 4.54 1.525 ;
      RECT  3.78 1.525 4.54 1.56 ;
      RECT  3.78 1.56 4.57 1.625 ;
      RECT  4.395 1.625 4.57 1.66 ;
      RECT  1.61 0.215 2.49 0.33 ;
      RECT  4.945 0.19 5.08 0.36 ;
      RECT  4.98 0.36 5.08 0.99 ;
      RECT  4.94 0.99 5.08 1.16 ;
      RECT  3.215 0.45 3.335 0.565 ;
      RECT  3.215 0.565 3.835 0.665 ;
      RECT  3.735 0.29 3.835 0.565 ;
      RECT  3.215 0.665 3.32 1.225 ;
      RECT  2.825 0.545 3.02 0.665 ;
      RECT  2.825 0.665 2.915 0.855 ;
      RECT  2.44 0.725 2.53 0.855 ;
      RECT  2.44 0.855 3.095 0.955 ;
      RECT  2.99 0.955 3.095 1.15 ;
      RECT  2.835 1.15 3.095 1.25 ;
      RECT  5.98 0.455 6.1 0.755 ;
      RECT  5.98 0.755 6.26 0.855 ;
      RECT  5.655 0.71 5.755 0.855 ;
      RECT  5.655 0.855 6.26 0.925 ;
      RECT  5.655 0.925 6.1 0.95 ;
      RECT  5.98 0.95 6.1 1.19 ;
      RECT  3.41 0.775 3.5 1.105 ;
      RECT  3.41 1.105 4.075 1.195 ;
      RECT  3.955 0.25 4.075 1.105 ;
      RECT  5.455 0.275 5.565 1.24 ;
      RECT  4.225 0.4 4.33 1.26 ;
      RECT  4.225 1.26 4.345 1.345 ;
      RECT  2.07 0.465 2.32 0.585 ;
      RECT  2.23 0.585 2.32 1.185 ;
      RECT  2.23 1.185 2.745 1.26 ;
      RECT  0.885 0.495 0.985 1.26 ;
      RECT  0.885 1.26 2.745 1.275 ;
      RECT  2.655 1.275 2.745 1.345 ;
      RECT  0.885 1.275 2.32 1.38 ;
      RECT  2.655 1.345 4.345 1.435 ;
      RECT  5.195 0.255 5.315 1.33 ;
      RECT  5.195 1.33 5.68 1.42 ;
      RECT  5.59 1.42 5.68 1.555 ;
      RECT  5.59 1.555 6.055 1.655 ;
      RECT  2.425 1.39 2.545 1.47 ;
      RECT  1.37 1.47 2.545 1.59 ;
      RECT  0.695 1.105 0.795 1.535 ;
      LAYER M2 ;
      RECT  3.695 0.35 5.12 0.45 ;
      RECT  0.655 1.15 3.015 1.25 ;
      LAYER V1 ;
      RECT  3.735 0.35 3.835 0.45 ;
      RECT  4.98 0.35 5.08 0.45 ;
      RECT  0.695 1.15 0.795 1.25 ;
      RECT  2.875 1.15 2.975 1.25 ;
  END
END SEN_FSDPMQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPMQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, 2-to-1 muxed data inputs, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D1&S&!SE)|(!S&(!SE&D0))|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPMQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPMQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 4.85 1.25 ;
      RECT  4.75 1.25 5.12 1.34 ;
      RECT  5.025 1.34 5.12 1.55 ;
      RECT  5.025 1.55 5.515 1.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 ;
  END CK
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.075 0.71 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.105 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.505 0.51 6.65 0.69 ;
      RECT  6.55 0.69 6.65 1.11 ;
      RECT  6.505 1.11 6.65 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.64 ;
      RECT  0.27 0.64 0.45 0.82 ;
      RECT  1.11 0.35 1.43 0.45 ;
      RECT  1.34 0.45 1.43 0.71 ;
      RECT  1.34 0.71 1.86 0.89 ;
      LAYER M2 ;
      RECT  0.445 0.35 1.29 0.45 ;
      RECT  0.445 0.45 0.555 0.55 ;
      RECT  0.31 0.55 0.555 0.65 ;
      LAYER V1 ;
      RECT  0.35 0.55 0.45 0.65 ;
      RECT  1.15 0.35 1.25 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 ;
  END S
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.695 0.485 0.795 0.92 ;
      RECT  2.815 0.15 2.99 0.25 ;
      RECT  2.88 0.25 2.99 0.35 ;
      RECT  2.88 0.35 3.07 0.45 ;
      LAYER M2 ;
      RECT  1.41 0.35 3.07 0.45 ;
      RECT  1.41 0.45 1.51 0.55 ;
      RECT  0.655 0.55 1.51 0.65 ;
      LAYER V1 ;
      RECT  0.695 0.55 0.795 0.65 ;
      RECT  2.93 0.35 3.03 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.91 0.45 1.11 ;
      RECT  0.35 1.11 0.565 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  5.685 1.105 5.905 1.225 ;
      RECT  5.8 1.225 5.905 1.315 ;
      RECT  5.8 1.315 6.365 1.425 ;
      RECT  6.245 1.425 6.365 1.75 ;
      RECT  4.69 1.43 4.925 1.545 ;
      RECT  4.835 1.545 4.925 1.75 ;
      RECT  0.335 1.38 0.455 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  2.865 1.525 3.005 1.75 ;
      RECT  3.49 1.525 3.63 1.75 ;
      RECT  6.79 1.21 6.91 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  0.345 0.05 0.45 0.225 ;
      RECT  5.735 0.05 5.855 0.42 ;
      RECT  3.5 0.05 3.62 0.43 ;
      RECT  6.79 0.05 6.91 0.59 ;
      RECT  2.595 0.05 2.715 0.61 ;
      RECT  4.76 0.05 4.87 0.61 ;
      RECT  6.245 0.05 6.365 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.54 0.14 1.435 0.24 ;
      RECT  0.54 0.24 0.63 0.315 ;
      RECT  0.075 0.315 0.63 0.405 ;
      RECT  0.075 0.405 0.195 0.515 ;
      RECT  0.075 0.515 0.18 1.37 ;
      RECT  0.075 1.37 0.195 1.61 ;
      RECT  4.385 0.145 4.61 0.315 ;
      RECT  4.49 0.315 4.61 0.565 ;
      RECT  4.435 0.565 4.61 0.67 ;
      RECT  4.435 0.67 4.555 1.165 ;
      RECT  4.465 1.165 4.555 1.525 ;
      RECT  3.79 1.525 4.555 1.56 ;
      RECT  3.79 1.56 4.585 1.625 ;
      RECT  4.41 1.625 4.585 1.66 ;
      RECT  1.61 0.215 2.48 0.33 ;
      RECT  4.965 0.19 5.095 0.36 ;
      RECT  4.995 0.36 5.095 0.99 ;
      RECT  4.945 0.99 5.095 1.16 ;
      RECT  3.23 0.45 3.35 0.565 ;
      RECT  3.23 0.565 3.85 0.665 ;
      RECT  3.75 0.29 3.85 0.565 ;
      RECT  3.23 0.665 3.335 1.2 ;
      RECT  2.84 0.545 3.035 0.665 ;
      RECT  2.84 0.665 2.93 0.855 ;
      RECT  2.45 0.725 2.55 0.855 ;
      RECT  2.45 0.855 3.11 0.955 ;
      RECT  3.005 0.955 3.11 1.15 ;
      RECT  2.85 1.15 3.11 1.25 ;
      RECT  5.995 0.42 6.115 0.79 ;
      RECT  5.995 0.79 6.45 0.855 ;
      RECT  5.67 0.7 5.77 0.855 ;
      RECT  5.67 0.855 6.45 0.89 ;
      RECT  5.67 0.89 6.115 0.95 ;
      RECT  5.995 0.95 6.115 1.19 ;
      RECT  3.425 0.775 3.515 1.105 ;
      RECT  3.425 1.105 4.09 1.195 ;
      RECT  3.97 0.245 4.09 1.105 ;
      RECT  4.24 0.4 4.345 1.26 ;
      RECT  4.24 1.26 4.36 1.345 ;
      RECT  2.07 0.465 2.32 0.585 ;
      RECT  2.23 0.585 2.32 1.185 ;
      RECT  2.23 1.185 2.76 1.26 ;
      RECT  0.885 0.52 0.985 1.26 ;
      RECT  0.885 1.26 2.76 1.275 ;
      RECT  2.67 1.275 2.76 1.345 ;
      RECT  0.885 1.275 2.32 1.38 ;
      RECT  2.67 1.345 4.36 1.435 ;
      RECT  5.47 0.2 5.58 1.265 ;
      RECT  5.21 0.2 5.33 1.355 ;
      RECT  5.21 1.355 5.695 1.445 ;
      RECT  5.605 1.445 5.695 1.55 ;
      RECT  5.605 1.55 6.095 1.655 ;
      RECT  2.44 1.39 2.56 1.47 ;
      RECT  1.37 1.47 2.56 1.59 ;
      RECT  0.695 1.105 0.795 1.535 ;
      LAYER M2 ;
      RECT  3.71 0.35 5.135 0.45 ;
      RECT  0.655 1.15 3.03 1.25 ;
      LAYER V1 ;
      RECT  3.75 0.35 3.85 0.45 ;
      RECT  4.995 0.35 5.095 0.45 ;
      RECT  0.695 1.15 0.795 1.25 ;
      RECT  2.89 1.15 2.99 1.25 ;
  END
END SEN_FSDPMQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPMQ_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, 2-to-1 muxed data inputs, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D1&S&!SE)|(!S&(!SE&D0))|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPMQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDPMQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 4.85 1.25 ;
      RECT  4.75 1.25 5.12 1.34 ;
      RECT  5.025 1.34 5.12 1.55 ;
      RECT  5.025 1.55 5.515 1.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12 ;
  END CK
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.075 0.71 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.105 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.51 7.095 0.69 ;
      RECT  6.95 0.69 7.05 1.11 ;
      RECT  6.44 1.11 7.095 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.64 ;
      RECT  0.27 0.64 0.45 0.82 ;
      RECT  1.11 0.35 1.435 0.45 ;
      RECT  1.34 0.45 1.435 0.71 ;
      RECT  1.34 0.71 1.86 0.89 ;
      LAYER M2 ;
      RECT  0.445 0.35 1.29 0.45 ;
      RECT  0.445 0.45 0.555 0.55 ;
      RECT  0.31 0.55 0.555 0.65 ;
      LAYER V1 ;
      RECT  0.35 0.55 0.45 0.65 ;
      RECT  1.15 0.35 1.25 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0888 ;
  END S
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.695 0.485 0.795 0.92 ;
      RECT  2.815 0.15 2.99 0.25 ;
      RECT  2.88 0.25 2.99 0.35 ;
      RECT  2.88 0.35 3.07 0.45 ;
      LAYER M2 ;
      RECT  1.41 0.35 3.07 0.45 ;
      RECT  1.41 0.45 1.51 0.55 ;
      RECT  0.655 0.55 1.51 0.65 ;
      LAYER V1 ;
      RECT  0.695 0.55 0.795 0.65 ;
      RECT  2.93 0.35 3.03 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.91 0.57 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  5.685 1.105 5.885 1.225 ;
      RECT  5.785 1.225 5.885 1.315 ;
      RECT  5.785 1.315 6.3 1.425 ;
      RECT  6.18 1.425 6.3 1.75 ;
      RECT  4.675 1.43 4.925 1.545 ;
      RECT  4.835 1.545 4.925 1.75 ;
      RECT  0.335 1.4 0.455 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  2.865 1.525 3.005 1.75 ;
      RECT  3.49 1.525 3.63 1.75 ;
      RECT  6.7 1.39 6.82 1.75 ;
      RECT  7.21 1.41 7.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  0.345 0.05 0.45 0.225 ;
      RECT  7.21 0.05 7.34 0.39 ;
      RECT  6.18 0.05 6.3 0.41 ;
      RECT  6.7 0.05 6.82 0.41 ;
      RECT  5.735 0.05 5.855 0.425 ;
      RECT  3.5 0.05 3.62 0.43 ;
      RECT  2.595 0.05 2.715 0.585 ;
      RECT  4.76 0.05 4.87 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.54 0.14 1.435 0.24 ;
      RECT  0.54 0.24 0.63 0.315 ;
      RECT  0.075 0.315 0.63 0.405 ;
      RECT  0.075 0.405 0.195 0.515 ;
      RECT  0.075 0.515 0.18 1.37 ;
      RECT  0.075 1.37 0.195 1.61 ;
      RECT  4.385 0.145 4.62 0.315 ;
      RECT  4.5 0.315 4.62 0.565 ;
      RECT  4.435 0.565 4.62 0.67 ;
      RECT  4.435 0.67 4.555 1.165 ;
      RECT  4.465 1.165 4.555 1.525 ;
      RECT  3.79 1.525 4.555 1.56 ;
      RECT  3.79 1.56 4.585 1.625 ;
      RECT  4.41 1.625 4.585 1.66 ;
      RECT  1.61 0.215 2.48 0.33 ;
      RECT  4.96 0.19 5.095 0.36 ;
      RECT  4.995 0.36 5.095 0.99 ;
      RECT  4.945 0.99 5.095 1.16 ;
      RECT  3.23 0.45 3.35 0.57 ;
      RECT  3.23 0.57 3.85 0.67 ;
      RECT  3.75 0.29 3.85 0.57 ;
      RECT  3.23 0.67 3.335 1.225 ;
      RECT  2.84 0.545 3.035 0.665 ;
      RECT  2.84 0.665 2.93 0.855 ;
      RECT  2.455 0.725 2.545 0.855 ;
      RECT  2.455 0.855 3.11 0.955 ;
      RECT  3.005 0.955 3.11 1.15 ;
      RECT  2.84 1.15 3.11 1.25 ;
      RECT  5.995 0.495 6.115 0.79 ;
      RECT  5.995 0.79 6.84 0.86 ;
      RECT  5.67 0.725 5.77 0.86 ;
      RECT  5.67 0.86 6.84 0.89 ;
      RECT  5.67 0.89 6.115 0.955 ;
      RECT  5.995 0.955 6.115 1.19 ;
      RECT  3.425 0.775 3.515 1.105 ;
      RECT  3.425 1.105 4.09 1.195 ;
      RECT  3.97 0.245 4.09 1.105 ;
      RECT  5.47 0.2 5.58 1.24 ;
      RECT  4.24 0.405 4.345 1.26 ;
      RECT  4.24 1.26 4.36 1.345 ;
      RECT  2.07 0.465 2.32 0.585 ;
      RECT  2.23 0.585 2.32 1.185 ;
      RECT  2.23 1.185 2.75 1.26 ;
      RECT  0.885 0.495 0.985 1.26 ;
      RECT  0.885 1.26 2.75 1.275 ;
      RECT  2.66 1.275 2.75 1.345 ;
      RECT  0.885 1.275 2.32 1.38 ;
      RECT  2.66 1.345 4.36 1.435 ;
      RECT  5.21 0.2 5.33 1.33 ;
      RECT  5.21 1.33 5.695 1.42 ;
      RECT  5.605 1.42 5.695 1.55 ;
      RECT  5.605 1.55 6.07 1.655 ;
      RECT  2.44 1.39 2.56 1.47 ;
      RECT  1.37 1.47 2.56 1.59 ;
      RECT  0.695 1.02 0.795 1.485 ;
      LAYER M2 ;
      RECT  3.71 0.35 5.135 0.45 ;
      RECT  0.655 1.15 3.03 1.25 ;
      LAYER V1 ;
      RECT  3.75 0.35 3.85 0.45 ;
      RECT  4.995 0.35 5.095 0.45 ;
      RECT  0.695 1.15 0.795 1.25 ;
      RECT  2.89 1.15 2.99 1.25 ;
  END
END SEN_FSDPMQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPMQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, 2-to-1 muxed data inputs, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D1&S&!SE)|(!S&(!SE&D0))|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPMQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDPMQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.585 0.585 5.675 0.83 ;
      RECT  5.585 0.83 5.695 0.92 ;
      RECT  5.605 0.92 5.695 1.21 ;
      RECT  4.815 0.71 5.05 0.9 ;
      RECT  4.95 0.9 5.05 0.98 ;
      RECT  4.95 0.98 5.25 1.08 ;
      RECT  5.15 1.08 5.25 1.21 ;
      RECT  5.15 1.21 5.695 1.3 ;
      RECT  5.345 1.3 5.45 1.57 ;
      RECT  5.345 1.57 5.98 1.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0747 ;
  END CK
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.075 0.71 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.115 0.91 ;
      RECT  1.95 0.91 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.22 0.51 7.355 0.69 ;
      RECT  7.265 0.69 7.355 1.11 ;
      RECT  7.15 1.11 7.355 1.49 ;
    END
    ANTENNADIFFAREA 0.139 ;
  END Q
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.65 ;
      RECT  0.27 0.65 0.45 0.82 ;
      RECT  1.11 0.35 1.45 0.45 ;
      RECT  1.34 0.45 1.45 0.71 ;
      RECT  1.34 0.71 1.86 0.91 ;
      RECT  1.75 0.51 1.86 0.71 ;
      RECT  1.34 0.91 1.45 1.09 ;
      LAYER M2 ;
      RECT  0.445 0.35 1.29 0.45 ;
      RECT  0.445 0.45 0.555 0.55 ;
      RECT  0.31 0.55 0.555 0.65 ;
      LAYER V1 ;
      RECT  0.35 0.55 0.45 0.65 ;
      RECT  1.15 0.35 1.25 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0915 ;
  END S
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.695 0.485 0.795 1.035 ;
      RECT  2.8 0.15 2.975 0.25 ;
      RECT  2.865 0.25 2.975 0.35 ;
      RECT  2.865 0.35 3.055 0.45 ;
      LAYER M2 ;
      RECT  1.41 0.35 3.055 0.45 ;
      RECT  1.41 0.45 1.51 0.55 ;
      RECT  0.655 0.55 1.51 0.65 ;
      LAYER V1 ;
      RECT  0.695 0.55 0.795 0.65 ;
      RECT  2.915 0.35 3.015 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.91 0.565 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.715 0.31 6.85 0.535 ;
      RECT  6.75 0.535 6.85 0.985 ;
      RECT  6.7 0.985 6.85 1.29 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.38 0.455 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  2.69 1.56 2.81 1.75 ;
      RECT  3.435 1.515 3.575 1.75 ;
      RECT  4.655 1.43 4.775 1.75 ;
      RECT  5.08 1.425 5.2 1.75 ;
      RECT  6.165 1.64 6.335 1.75 ;
      RECT  6.955 1.04 7.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  5.075 0.05 5.245 0.19 ;
      RECT  0.345 0.05 0.45 0.225 ;
      RECT  6.965 0.05 7.085 0.41 ;
      RECT  4.655 0.05 4.775 0.42 ;
      RECT  3.445 0.05 3.565 0.455 ;
      RECT  6.21 0.05 6.33 0.46 ;
      RECT  2.58 0.05 2.7 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  5.38 0.14 6.01 0.23 ;
      RECT  5.38 0.23 5.47 0.28 ;
      RECT  4.915 0.28 5.47 0.37 ;
      RECT  4.915 0.37 5.035 0.52 ;
      RECT  4.585 0.52 5.035 0.62 ;
      RECT  4.585 0.62 4.675 0.775 ;
      RECT  4.56 0.775 4.675 1.24 ;
      RECT  4.56 1.24 5.045 1.25 ;
      RECT  4.93 1.17 5.045 1.24 ;
      RECT  4.44 1.25 5.045 1.34 ;
      RECT  4.44 1.34 4.53 1.525 ;
      RECT  3.74 1.525 4.53 1.625 ;
      RECT  0.54 0.14 1.435 0.24 ;
      RECT  0.54 0.24 0.63 0.315 ;
      RECT  0.075 0.315 0.63 0.405 ;
      RECT  0.075 0.405 0.195 0.515 ;
      RECT  0.075 0.515 0.18 1.37 ;
      RECT  0.075 1.37 0.195 1.61 ;
      RECT  1.61 0.215 2.49 0.33 ;
      RECT  6.475 0.29 6.61 0.46 ;
      RECT  6.52 0.46 6.61 1.01 ;
      RECT  6.155 0.875 6.245 1.01 ;
      RECT  6.155 1.01 6.61 1.105 ;
      RECT  6.47 1.105 6.61 1.37 ;
      RECT  5.605 0.355 5.875 0.475 ;
      RECT  5.775 0.475 5.875 0.69 ;
      RECT  5.785 0.69 5.875 1.39 ;
      RECT  5.58 1.39 5.875 1.48 ;
      RECT  4.175 0.21 4.28 0.505 ;
      RECT  4.115 0.505 4.28 0.605 ;
      RECT  4.115 0.605 4.205 1.11 ;
      RECT  4.115 1.11 4.215 1.325 ;
      RECT  4.115 1.325 4.35 1.435 ;
      RECT  5.965 0.32 6.065 0.505 ;
      RECT  5.975 0.505 6.065 1.165 ;
      RECT  5.965 1.165 6.065 1.39 ;
      RECT  5.965 1.39 6.3 1.46 ;
      RECT  5.965 1.46 6.72 1.48 ;
      RECT  6.21 1.48 6.72 1.55 ;
      RECT  6.63 1.55 6.72 1.57 ;
      RECT  6.63 1.57 6.85 1.66 ;
      RECT  3.175 0.38 3.295 0.55 ;
      RECT  3.175 0.55 3.795 0.65 ;
      RECT  3.175 0.65 3.28 1.19 ;
      RECT  2.07 0.495 2.295 0.615 ;
      RECT  2.205 0.615 2.295 1.0 ;
      RECT  2.14 1.0 2.295 1.1 ;
      RECT  2.14 1.1 2.24 1.29 ;
      RECT  6.17 0.55 6.43 0.65 ;
      RECT  6.33 0.65 6.43 0.845 ;
      RECT  2.825 0.545 3.02 0.665 ;
      RECT  2.825 0.665 2.915 0.775 ;
      RECT  2.385 0.7 2.485 0.775 ;
      RECT  2.385 0.775 2.915 0.875 ;
      RECT  2.435 0.875 2.555 1.185 ;
      RECT  2.33 1.185 2.555 1.275 ;
      RECT  2.33 1.275 2.42 1.38 ;
      RECT  1.135 1.285 1.81 1.375 ;
      RECT  1.72 1.375 1.81 1.38 ;
      RECT  1.135 1.375 1.225 1.395 ;
      RECT  1.72 1.38 2.42 1.47 ;
      RECT  0.695 1.125 0.795 1.395 ;
      RECT  0.695 1.395 1.225 1.485 ;
      RECT  4.37 0.495 4.495 0.69 ;
      RECT  4.37 0.69 4.47 0.75 ;
      RECT  4.295 0.75 4.47 0.92 ;
      RECT  4.37 0.92 4.47 1.16 ;
      RECT  6.95 0.51 7.05 0.755 ;
      RECT  6.95 0.755 7.155 0.925 ;
      RECT  5.17 0.51 5.285 0.89 ;
      RECT  5.375 0.46 5.485 1.03 ;
      RECT  5.345 1.03 5.515 1.12 ;
      RECT  3.37 0.74 3.47 1.13 ;
      RECT  3.37 1.13 4.025 1.22 ;
      RECT  3.915 0.245 4.025 1.13 ;
      RECT  0.885 0.465 0.985 1.29 ;
      RECT  2.51 1.37 3.175 1.46 ;
      RECT  2.51 1.46 2.6 1.57 ;
      RECT  3.005 1.46 3.175 1.66 ;
      RECT  1.39 1.465 1.565 1.57 ;
      RECT  1.39 1.57 2.6 1.66 ;
      LAYER M2 ;
      RECT  3.61 0.55 5.31 0.65 ;
      RECT  5.735 0.55 7.09 0.65 ;
      RECT  0.845 1.15 4.26 1.25 ;
      LAYER V1 ;
      RECT  3.65 0.55 3.75 0.65 ;
      RECT  5.17 0.55 5.27 0.65 ;
      RECT  5.775 0.55 5.875 0.65 ;
      RECT  6.24 0.55 6.34 0.65 ;
      RECT  6.95 0.55 7.05 0.65 ;
      RECT  0.885 1.15 0.985 1.25 ;
      RECT  2.14 1.15 2.24 1.25 ;
      RECT  4.115 1.15 4.215 1.25 ;
  END
END SEN_FSDPMQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPMQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, 2-to-1 muxed data inputs, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D1&S&!SE)|(!S&(!SE&D0))|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPMQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDPMQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.8 0.74 7.205 0.84 ;
      RECT  6.8 0.84 6.9 1.25 ;
      RECT  6.2 0.71 6.45 0.89 ;
      RECT  6.35 0.89 6.45 1.25 ;
      RECT  6.35 1.25 6.9 1.295 ;
      RECT  6.35 1.295 7.16 1.34 ;
      RECT  6.8 1.34 7.16 1.385 ;
      RECT  7.07 1.385 7.16 1.56 ;
      RECT  7.07 1.56 8.015 1.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0957 ;
  END CK
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.12 0.875 1.385 1.07 ;
      LAYER M2 ;
      RECT  1.14 0.95 1.745 1.05 ;
      LAYER V1 ;
      RECT  1.23 0.95 1.33 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0816 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.885 0.69 2.985 0.845 ;
      RECT  2.71 0.845 2.985 0.955 ;
      LAYER M2 ;
      RECT  2.81 0.75 3.49 0.85 ;
      LAYER V1 ;
      RECT  2.885 0.75 2.985 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0816 ;
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.35 0.51 9.65 0.69 ;
      RECT  9.55 0.69 9.65 1.11 ;
      RECT  9.345 1.11 9.65 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.59 2.795 0.69 ;
      RECT  2.41 0.69 2.51 0.95 ;
      RECT  1.735 0.87 1.855 0.95 ;
      RECT  1.735 0.95 2.51 1.04 ;
      RECT  0.26 0.71 0.36 0.75 ;
      RECT  0.26 0.75 0.605 0.89 ;
      LAYER M2 ;
      RECT  0.425 0.75 2.55 0.85 ;
      LAYER V1 ;
      RECT  2.41 0.75 2.51 0.85 ;
      RECT  0.465 0.75 0.565 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1185 ;
  END S
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.125 0.51 4.225 1.035 ;
      RECT  3.7 1.035 4.225 1.14 ;
      RECT  0.43 0.55 0.79 0.65 ;
      RECT  0.695 0.65 0.79 0.775 ;
      LAYER M2 ;
      RECT  0.525 0.55 4.265 0.65 ;
      LAYER V1 ;
      RECT  4.125 0.55 4.225 0.65 ;
      RECT  0.565 0.55 0.665 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.087 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.09 0.65 1.29 ;
      RECT  0.55 1.29 0.65 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.85 0.51 9.05 0.665 ;
      RECT  8.95 0.665 9.05 1.02 ;
      RECT  8.835 1.02 9.05 1.11 ;
      RECT  8.835 1.11 8.96 1.31 ;
    END
    ANTENNADIFFAREA 0.11 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.39 0.445 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  3.34 1.61 3.51 1.75 ;
      RECT  3.97 1.23 4.09 1.75 ;
      RECT  5.485 1.43 5.605 1.75 ;
      RECT  6.28 1.43 6.45 1.75 ;
      RECT  6.81 1.475 6.98 1.75 ;
      RECT  8.2 1.535 8.345 1.75 ;
      RECT  8.525 1.475 8.675 1.75 ;
      RECT  9.085 1.195 9.205 1.75 ;
      RECT  9.595 1.41 9.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  3.7 0.05 3.87 0.2 ;
      RECT  4.05 0.05 4.22 0.2 ;
      RECT  6.375 0.05 6.53 0.24 ;
      RECT  6.92 0.05 7.07 0.24 ;
      RECT  8.125 0.05 8.295 0.26 ;
      RECT  0.335 0.05 0.455 0.28 ;
      RECT  9.595 0.05 9.735 0.39 ;
      RECT  5.865 0.05 5.97 0.41 ;
      RECT  9.075 0.05 9.215 0.41 ;
      RECT  5.35 0.05 5.52 0.515 ;
      RECT  8.64 0.05 8.76 0.655 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.715 0.14 2.305 0.2 ;
      RECT  1.11 0.2 2.305 0.26 ;
      RECT  1.11 0.26 1.805 0.32 ;
      RECT  2.185 0.26 2.305 0.32 ;
      RECT  7.305 0.155 7.95 0.255 ;
      RECT  7.305 0.255 7.395 0.33 ;
      RECT  6.125 0.33 7.395 0.42 ;
      RECT  6.125 0.42 6.245 0.485 ;
      RECT  6.02 0.485 6.245 0.575 ;
      RECT  6.02 0.575 6.11 0.785 ;
      RECT  5.51 0.785 6.11 0.885 ;
      RECT  5.99 0.885 6.11 1.2 ;
      RECT  2.405 0.175 3.11 0.265 ;
      RECT  2.405 0.265 2.59 0.32 ;
      RECT  2.93 0.265 3.11 0.32 ;
      RECT  3.62 0.29 4.76 0.38 ;
      RECT  4.64 0.38 4.76 0.525 ;
      RECT  3.62 0.38 3.71 0.64 ;
      RECT  4.64 0.525 4.78 0.625 ;
      RECT  4.675 0.625 4.78 1.225 ;
      RECT  3.075 0.61 3.395 0.64 ;
      RECT  3.075 0.64 3.71 0.73 ;
      RECT  3.075 0.73 3.165 1.045 ;
      RECT  2.64 1.045 3.165 1.135 ;
      RECT  0.885 0.59 1.585 0.68 ;
      RECT  0.885 0.68 1.03 0.785 ;
      RECT  1.48 0.68 1.585 1.135 ;
      RECT  0.94 0.785 1.03 1.44 ;
      RECT  1.48 1.135 2.81 1.225 ;
      RECT  0.835 1.44 1.03 1.495 ;
      RECT  0.835 1.495 1.51 1.61 ;
      RECT  0.065 0.37 0.985 0.41 ;
      RECT  0.065 0.41 1.785 0.46 ;
      RECT  0.88 0.46 1.785 0.5 ;
      RECT  0.065 0.46 0.17 1.515 ;
      RECT  1.695 0.5 1.785 0.645 ;
      RECT  1.695 0.645 2.23 0.745 ;
      RECT  1.925 0.35 2.03 0.41 ;
      RECT  1.925 0.41 3.53 0.5 ;
      RECT  2.68 0.37 2.85 0.41 ;
      RECT  3.42 0.19 3.53 0.41 ;
      RECT  1.925 0.5 2.03 0.52 ;
      RECT  4.87 0.405 5.025 0.585 ;
      RECT  4.87 0.585 4.96 1.04 ;
      RECT  4.87 1.04 5.035 1.13 ;
      RECT  4.925 1.13 5.035 1.315 ;
      RECT  4.495 0.745 4.585 1.315 ;
      RECT  4.495 1.315 5.035 1.405 ;
      RECT  5.635 0.445 5.755 0.605 ;
      RECT  5.125 0.605 5.755 0.695 ;
      RECT  5.125 0.695 5.215 0.73 ;
      RECT  5.05 0.73 5.215 0.9 ;
      RECT  5.125 0.9 5.215 0.99 ;
      RECT  5.125 0.99 5.875 1.16 ;
      RECT  6.59 0.515 7.535 0.635 ;
      RECT  6.59 0.635 6.71 1.035 ;
      RECT  7.43 0.635 7.535 1.225 ;
      RECT  6.54 1.035 6.71 1.16 ;
      RECT  8.23 0.53 8.55 0.65 ;
      RECT  8.23 0.65 8.34 0.815 ;
      RECT  8.065 0.815 8.34 0.985 ;
      RECT  8.215 0.985 8.34 1.17 ;
      RECT  3.8 0.535 4.035 0.705 ;
      RECT  3.8 0.705 3.89 0.845 ;
      RECT  3.255 0.845 3.89 0.945 ;
      RECT  3.255 0.945 3.36 1.225 ;
      RECT  3.13 1.225 3.36 1.33 ;
      RECT  8.655 0.785 8.86 0.89 ;
      RECT  8.655 0.89 8.745 1.26 ;
      RECT  7.875 0.415 7.995 0.61 ;
      RECT  7.875 0.61 7.975 1.115 ;
      RECT  7.875 1.115 8.02 1.215 ;
      RECT  7.92 1.215 8.02 1.26 ;
      RECT  7.92 1.26 8.745 1.35 ;
      RECT  7.92 1.35 8.09 1.445 ;
      RECT  9.145 0.785 9.44 0.895 ;
      RECT  9.145 0.895 9.245 1.09 ;
      RECT  8.44 0.75 8.565 1.115 ;
      RECT  0.74 0.895 0.85 1.3 ;
      RECT  7.625 0.42 7.74 1.305 ;
      RECT  7.625 1.305 7.83 1.335 ;
      RECT  7.095 1.095 7.34 1.205 ;
      RECT  7.25 1.205 7.34 1.335 ;
      RECT  7.25 1.335 7.83 1.425 ;
      RECT  1.12 1.2 1.225 1.315 ;
      RECT  1.12 1.315 2.055 1.405 ;
      RECT  2.925 1.31 3.04 1.315 ;
      RECT  2.355 1.315 3.04 1.405 ;
      RECT  2.925 1.405 3.04 1.48 ;
      RECT  5.295 1.25 5.805 1.34 ;
      RECT  5.295 1.34 5.395 1.495 ;
      RECT  5.715 1.34 5.805 1.54 ;
      RECT  4.315 0.47 4.51 0.64 ;
      RECT  4.315 0.64 4.405 1.4 ;
      RECT  4.2 1.4 4.405 1.495 ;
      RECT  4.2 1.495 5.395 1.52 ;
      RECT  4.315 1.52 5.395 1.585 ;
      RECT  5.715 1.54 6.08 1.64 ;
      RECT  3.135 1.42 3.855 1.52 ;
      RECT  3.135 1.52 3.225 1.57 ;
      RECT  1.6 1.495 2.82 1.57 ;
      RECT  1.6 1.57 3.225 1.6 ;
      RECT  2.715 1.6 3.225 1.66 ;
      LAYER M2 ;
      RECT  7.59 0.95 9.285 1.05 ;
      RECT  0.71 1.15 3.395 1.25 ;
      LAYER V1 ;
      RECT  7.63 0.95 7.73 1.05 ;
      RECT  8.44 0.95 8.54 1.05 ;
      RECT  9.145 0.95 9.245 1.05 ;
      RECT  0.75 1.15 0.85 1.25 ;
      RECT  3.255 1.15 3.355 1.25 ;
  END
END SEN_FSDPMQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPMQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, 2-to-1 muxed data inputs, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(D1&S&!SE)|(!S&(!SE&D0))|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPMQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDPMQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.33 0.71 7.65 0.89 ;
      RECT  7.55 0.89 7.65 1.245 ;
      RECT  7.55 1.245 8.45 1.335 ;
      RECT  8.35 1.335 8.45 1.355 ;
      RECT  8.35 1.355 8.575 1.525 ;
      RECT  8.485 1.525 8.575 1.56 ;
      RECT  8.485 1.56 9.495 1.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1245 ;
  END CK
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.12 0.875 1.385 1.07 ;
      LAYER M2 ;
      RECT  1.14 0.95 1.745 1.05 ;
      LAYER V1 ;
      RECT  1.23 0.95 1.33 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1062 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.745 3.13 1.03 ;
      LAYER M2 ;
      RECT  2.875 0.75 3.555 0.85 ;
      LAYER V1 ;
      RECT  2.99 0.75 3.09 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1062 ;
  END D1
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.75 0.51 11.47 0.69 ;
      RECT  11.35 0.69 11.47 1.11 ;
      RECT  10.835 1.11 11.47 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.735 0.87 1.855 0.95 ;
      RECT  1.735 0.95 2.72 1.04 ;
      RECT  2.62 0.61 2.72 0.95 ;
      RECT  0.26 0.71 0.36 0.75 ;
      RECT  0.26 0.75 0.605 0.89 ;
      LAYER M2 ;
      RECT  0.425 0.75 2.76 0.85 ;
      LAYER V1 ;
      RECT  2.62 0.75 2.72 0.85 ;
      RECT  0.465 0.75 0.565 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1545 ;
  END S
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.49 4.85 0.835 ;
      RECT  4.595 0.835 4.85 1.09 ;
      RECT  0.43 0.55 0.79 0.65 ;
      RECT  0.695 0.65 0.79 0.745 ;
      LAYER M2 ;
      RECT  0.525 0.55 4.89 0.65 ;
      LAYER V1 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  0.565 0.55 0.665 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1035 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.055 0.65 1.29 ;
      RECT  0.55 1.29 0.65 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.35 0.31 10.45 0.545 ;
      RECT  10.35 0.545 10.535 0.69 ;
      RECT  10.44 0.69 10.535 1.02 ;
      RECT  10.325 1.02 10.535 1.11 ;
      RECT  10.325 1.11 10.45 1.31 ;
    END
    ANTENNADIFFAREA 0.11 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  6.95 1.0 7.06 1.325 ;
      RECT  6.95 1.325 7.385 1.415 ;
      RECT  7.295 1.415 7.385 1.425 ;
      RECT  7.295 1.425 7.705 1.515 ;
      RECT  7.535 1.515 7.705 1.75 ;
      RECT  0.31 1.39 0.46 1.75 ;
      RECT  0.0 1.75 11.8 1.85 ;
      RECT  3.87 1.61 4.04 1.75 ;
      RECT  4.54 1.39 4.69 1.75 ;
      RECT  5.175 1.64 5.345 1.75 ;
      RECT  6.45 1.43 6.57 1.75 ;
      RECT  8.055 1.425 8.225 1.75 ;
      RECT  9.69 1.535 9.835 1.75 ;
      RECT  10.015 1.46 10.165 1.75 ;
      RECT  10.585 1.19 10.695 1.75 ;
      RECT  11.095 1.39 11.215 1.75 ;
      RECT  11.615 1.21 11.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.8 0.05 ;
      RECT  5.245 0.05 5.415 0.195 ;
      RECT  4.295 0.05 4.465 0.2 ;
      RECT  4.64 0.05 4.81 0.2 ;
      RECT  7.46 0.05 7.615 0.24 ;
      RECT  8.005 0.05 8.155 0.24 ;
      RECT  0.32 0.05 0.47 0.28 ;
      RECT  3.77 0.05 3.9 0.305 ;
      RECT  6.425 0.05 6.595 0.405 ;
      RECT  10.585 0.05 10.695 0.41 ;
      RECT  11.095 0.05 11.215 0.41 ;
      RECT  9.64 0.05 9.76 0.415 ;
      RECT  6.95 0.05 7.07 0.42 ;
      RECT  11.615 0.05 11.735 0.59 ;
      RECT  10.13 0.05 10.25 0.655 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.59 0.14 2.33 0.2 ;
      RECT  1.11 0.2 2.33 0.28 ;
      RECT  1.11 0.28 1.7 0.32 ;
      RECT  8.285 0.155 9.39 0.255 ;
      RECT  8.285 0.255 8.375 0.33 ;
      RECT  7.21 0.33 8.375 0.42 ;
      RECT  7.21 0.42 7.33 0.485 ;
      RECT  7.15 0.485 7.33 0.575 ;
      RECT  7.15 0.575 7.24 0.765 ;
      RECT  6.56 0.765 7.24 0.865 ;
      RECT  7.15 0.865 7.24 1.03 ;
      RECT  7.15 1.03 7.38 1.155 ;
      RECT  2.42 0.2 3.68 0.32 ;
      RECT  4.235 0.29 5.595 0.38 ;
      RECT  4.235 0.38 4.325 0.64 ;
      RECT  5.475 0.38 5.595 0.85 ;
      RECT  3.24 0.59 3.42 0.64 ;
      RECT  3.24 0.64 4.325 0.695 ;
      RECT  3.33 0.695 4.325 0.73 ;
      RECT  3.33 0.73 3.42 1.135 ;
      RECT  5.475 0.85 5.69 0.94 ;
      RECT  5.6 0.94 5.69 1.09 ;
      RECT  5.6 1.09 5.825 1.19 ;
      RECT  0.885 0.61 1.585 0.7 ;
      RECT  0.885 0.7 1.03 0.785 ;
      RECT  1.48 0.7 1.585 1.135 ;
      RECT  0.94 0.785 1.03 1.44 ;
      RECT  1.48 1.135 3.42 1.225 ;
      RECT  0.835 1.44 1.03 1.495 ;
      RECT  0.835 1.495 1.51 1.61 ;
      RECT  0.065 0.37 0.985 0.41 ;
      RECT  0.065 0.41 1.785 0.46 ;
      RECT  0.88 0.46 1.785 0.5 ;
      RECT  0.065 0.46 0.17 1.41 ;
      RECT  1.695 0.5 1.785 0.66 ;
      RECT  1.695 0.66 2.36 0.75 ;
      RECT  2.255 0.75 2.36 0.83 ;
      RECT  1.915 0.38 2.03 0.41 ;
      RECT  1.915 0.41 4.145 0.5 ;
      RECT  4.045 0.28 4.145 0.41 ;
      RECT  1.915 0.5 2.03 0.55 ;
      RECT  8.535 0.375 9.22 0.495 ;
      RECT  9.12 0.495 9.22 1.305 ;
      RECT  9.12 1.305 9.32 1.335 ;
      RECT  8.595 1.04 8.795 1.16 ;
      RECT  8.695 1.16 8.795 1.335 ;
      RECT  8.695 1.335 9.32 1.425 ;
      RECT  7.75 0.52 8.44 0.585 ;
      RECT  7.75 0.585 9.025 0.64 ;
      RECT  8.35 0.64 9.025 0.705 ;
      RECT  7.75 0.64 7.87 1.04 ;
      RECT  8.905 0.705 9.025 1.215 ;
      RECT  7.75 1.04 8.46 1.155 ;
      RECT  8.34 0.96 8.46 1.04 ;
      RECT  6.175 0.495 6.89 0.615 ;
      RECT  6.175 0.615 6.265 0.69 ;
      RECT  5.96 0.69 6.265 0.795 ;
      RECT  6.175 0.795 6.265 0.99 ;
      RECT  6.175 0.99 6.845 1.16 ;
      RECT  5.76 0.41 5.87 0.635 ;
      RECT  5.78 0.635 5.87 0.89 ;
      RECT  5.78 0.89 6.035 0.98 ;
      RECT  5.915 0.98 6.035 1.28 ;
      RECT  5.215 0.745 5.315 1.075 ;
      RECT  5.215 1.075 5.51 1.165 ;
      RECT  5.4 1.165 5.51 1.28 ;
      RECT  5.4 1.28 6.035 1.37 ;
      RECT  9.72 0.53 10.04 0.65 ;
      RECT  9.72 0.65 9.83 0.815 ;
      RECT  9.555 0.815 9.83 0.985 ;
      RECT  9.705 0.985 9.83 1.16 ;
      RECT  4.415 0.495 4.645 0.665 ;
      RECT  4.415 0.665 4.505 1.21 ;
      RECT  3.625 0.82 3.775 0.99 ;
      RECT  3.67 0.99 3.775 1.21 ;
      RECT  3.67 1.21 4.505 1.3 ;
      RECT  10.145 0.785 10.35 0.89 ;
      RECT  10.145 0.89 10.235 1.26 ;
      RECT  9.365 0.4 9.485 0.61 ;
      RECT  9.365 0.61 9.465 1.115 ;
      RECT  9.365 1.115 9.51 1.215 ;
      RECT  9.41 1.215 9.51 1.26 ;
      RECT  9.41 1.26 10.235 1.35 ;
      RECT  9.41 1.35 9.58 1.445 ;
      RECT  10.635 0.785 11.24 0.895 ;
      RECT  10.635 0.895 10.735 1.09 ;
      RECT  9.93 0.75 10.055 1.115 ;
      RECT  0.74 0.895 0.85 1.3 ;
      RECT  1.12 1.2 1.225 1.315 ;
      RECT  1.12 1.315 2.055 1.405 ;
      RECT  6.26 1.25 6.78 1.34 ;
      RECT  6.26 1.34 6.36 1.46 ;
      RECT  6.69 1.34 6.78 1.54 ;
      RECT  5.005 0.47 5.105 1.3 ;
      RECT  4.865 1.3 5.105 1.42 ;
      RECT  5.005 1.42 5.105 1.46 ;
      RECT  5.005 1.46 6.36 1.55 ;
      RECT  6.69 1.54 7.205 1.64 ;
      RECT  2.355 1.315 3.575 1.405 ;
      RECT  3.665 1.4 4.355 1.52 ;
      RECT  3.665 1.52 3.755 1.57 ;
      RECT  1.6 1.495 2.82 1.57 ;
      RECT  1.6 1.57 3.755 1.6 ;
      RECT  2.715 1.6 3.755 1.66 ;
      LAYER M2 ;
      RECT  9.08 0.95 10.775 1.05 ;
      RECT  0.71 1.15 3.81 1.25 ;
      LAYER V1 ;
      RECT  9.12 0.95 9.22 1.05 ;
      RECT  9.93 0.95 10.03 1.05 ;
      RECT  10.635 0.95 10.735 1.05 ;
      RECT  0.75 1.15 0.85 1.25 ;
      RECT  3.67 1.15 3.77 1.25 ;
  END
END SEN_FSDPMQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQ_DV1_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQ_DV1_1
  CLASS CORE ;
  FOREIGN SEN_FSDPQ_DV1_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.57 0.89 3.67 1.105 ;
      RECT  3.57 1.105 3.94 1.195 ;
      RECT  2.27 0.72 2.36 0.865 ;
      RECT  2.27 0.865 3.115 0.955 ;
      RECT  3.025 0.73 3.115 0.865 ;
      RECT  3.015 0.955 3.115 1.11 ;
      LAYER M2 ;
      RECT  2.93 0.95 3.71 1.05 ;
      LAYER V1 ;
      RECT  3.57 0.95 3.67 1.05 ;
      RECT  3.015 0.95 3.115 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.51 1.05 0.71 ;
      RECT  0.94 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.51 4.945 0.69 ;
      RECT  4.84 0.69 4.945 1.11 ;
      RECT  4.55 1.11 4.945 1.29 ;
    END
    ANTENNADIFFAREA 0.139 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.55 0.71 0.85 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.575 0.6 ;
      RECT  0.35 0.6 0.45 1.065 ;
      RECT  0.35 1.065 1.45 1.155 ;
      RECT  1.35 0.71 1.45 1.065 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.43 0.445 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.425 1.48 1.61 1.75 ;
      RECT  2.64 1.23 2.745 1.75 ;
      RECT  2.92 1.43 3.04 1.75 ;
      RECT  4.075 1.465 4.245 1.75 ;
      RECT  4.565 1.39 4.685 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  1.32 0.05 1.41 0.345 ;
      RECT  2.92 0.05 3.04 0.36 ;
      RECT  0.325 0.05 0.445 0.405 ;
      RECT  4.565 0.05 4.685 0.41 ;
      RECT  2.64 0.05 2.755 0.585 ;
      RECT  4.1 0.05 4.22 0.63 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.5 0.18 1.94 0.27 ;
      RECT  1.85 0.27 1.94 0.325 ;
      RECT  1.5 0.27 1.59 0.435 ;
      RECT  1.85 0.325 2.09 0.445 ;
      RECT  0.735 0.215 1.23 0.335 ;
      RECT  1.14 0.335 1.23 0.435 ;
      RECT  1.14 0.435 1.59 0.525 ;
      RECT  3.205 0.18 3.94 0.27 ;
      RECT  3.205 0.27 3.295 0.45 ;
      RECT  2.845 0.45 3.295 0.54 ;
      RECT  2.845 0.54 2.935 0.675 ;
      RECT  3.205 0.54 3.295 1.16 ;
      RECT  2.04 0.14 2.54 0.23 ;
      RECT  2.45 0.23 2.54 0.675 ;
      RECT  2.45 0.675 2.935 0.765 ;
      RECT  0.045 0.19 0.185 0.41 ;
      RECT  0.045 0.41 0.135 1.25 ;
      RECT  0.045 1.25 0.625 1.34 ;
      RECT  0.535 1.34 0.625 1.52 ;
      RECT  0.045 1.34 0.185 1.62 ;
      RECT  0.535 1.52 1.25 1.63 ;
      RECT  2.18 0.37 2.3 0.54 ;
      RECT  1.885 0.54 2.3 0.63 ;
      RECT  1.885 0.63 1.975 0.76 ;
      RECT  1.85 0.76 1.975 0.9 ;
      RECT  1.85 0.9 2.15 0.99 ;
      RECT  2.06 0.99 2.15 1.06 ;
      RECT  2.06 1.06 2.34 1.16 ;
      RECT  3.585 0.445 3.87 0.565 ;
      RECT  3.78 0.565 3.87 0.925 ;
      RECT  3.78 0.925 4.28 1.015 ;
      RECT  4.095 1.015 4.28 1.13 ;
      RECT  4.095 1.13 4.185 1.285 ;
      RECT  3.64 1.285 4.185 1.375 ;
      RECT  3.64 1.375 3.76 1.61 ;
      RECT  4.31 0.17 4.425 0.645 ;
      RECT  4.31 0.645 4.45 0.735 ;
      RECT  4.0 0.735 4.45 0.78 ;
      RECT  4.0 0.78 4.75 0.835 ;
      RECT  4.37 0.835 4.75 0.95 ;
      RECT  4.37 0.95 4.46 1.22 ;
      RECT  4.275 1.22 4.46 1.325 ;
      RECT  2.43 1.05 2.925 1.14 ;
      RECT  2.43 1.14 2.52 1.25 ;
      RECT  2.835 1.14 2.925 1.25 ;
      RECT  1.68 0.51 1.785 0.605 ;
      RECT  1.635 0.605 1.785 0.685 ;
      RECT  1.635 0.685 1.725 1.08 ;
      RECT  1.635 1.08 1.97 1.2 ;
      RECT  1.88 1.2 1.97 1.25 ;
      RECT  1.88 1.25 2.52 1.34 ;
      RECT  2.835 1.25 3.48 1.34 ;
      RECT  3.385 0.44 3.48 1.25 ;
      RECT  3.37 1.34 3.48 1.61 ;
      RECT  0.895 1.29 1.79 1.39 ;
      RECT  1.7 1.39 1.79 1.46 ;
      RECT  1.7 1.46 2.08 1.58 ;
  END
END SEN_FSDPQ_DV1_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQ_DV1_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQ_DV1_2
  CLASS CORE ;
  FOREIGN SEN_FSDPQ_DV1_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.57 0.89 3.67 1.105 ;
      RECT  3.57 1.105 3.94 1.195 ;
      RECT  2.26 0.72 2.36 0.865 ;
      RECT  2.26 0.865 3.115 0.955 ;
      RECT  3.025 0.7 3.115 0.865 ;
      RECT  3.015 0.955 3.115 1.11 ;
      LAYER M2 ;
      RECT  2.93 0.95 3.71 1.05 ;
      LAYER V1 ;
      RECT  3.57 0.95 3.67 1.05 ;
      RECT  3.015 0.95 3.115 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.51 1.05 0.71 ;
      RECT  0.94 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.82 0.51 5.05 0.69 ;
      RECT  4.95 0.69 5.05 1.11 ;
      RECT  4.845 1.11 5.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.55 0.71 0.85 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.505 0.575 0.605 ;
      RECT  0.35 0.605 0.45 1.065 ;
      RECT  0.35 1.065 1.45 1.155 ;
      RECT  1.35 0.71 1.45 1.065 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.43 0.445 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  1.425 1.48 1.61 1.75 ;
      RECT  2.64 1.23 2.745 1.75 ;
      RECT  2.92 1.43 3.04 1.75 ;
      RECT  4.075 1.465 4.245 1.75 ;
      RECT  4.585 1.19 4.705 1.75 ;
      RECT  5.14 1.21 5.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  1.32 0.05 1.41 0.345 ;
      RECT  2.92 0.05 3.04 0.36 ;
      RECT  0.325 0.05 0.445 0.405 ;
      RECT  2.64 0.05 2.755 0.585 ;
      RECT  4.1 0.05 4.22 0.59 ;
      RECT  5.14 0.05 5.26 0.59 ;
      RECT  4.585 0.05 4.705 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.5 0.18 1.94 0.27 ;
      RECT  1.85 0.27 1.94 0.325 ;
      RECT  1.5 0.27 1.59 0.435 ;
      RECT  1.85 0.325 2.09 0.445 ;
      RECT  0.735 0.215 1.23 0.335 ;
      RECT  1.14 0.335 1.23 0.435 ;
      RECT  1.14 0.435 1.59 0.525 ;
      RECT  3.19 0.18 3.94 0.27 ;
      RECT  3.19 0.27 3.295 0.45 ;
      RECT  2.845 0.45 3.295 0.54 ;
      RECT  2.845 0.54 2.935 0.675 ;
      RECT  3.205 0.54 3.295 1.16 ;
      RECT  2.04 0.14 2.54 0.23 ;
      RECT  2.45 0.23 2.54 0.675 ;
      RECT  2.45 0.675 2.935 0.765 ;
      RECT  0.045 0.19 0.185 0.41 ;
      RECT  0.045 0.41 0.135 1.25 ;
      RECT  0.045 1.25 0.625 1.34 ;
      RECT  0.535 1.34 0.625 1.52 ;
      RECT  0.045 1.34 0.185 1.61 ;
      RECT  0.535 1.52 1.25 1.63 ;
      RECT  2.18 0.37 2.3 0.54 ;
      RECT  1.885 0.54 2.3 0.63 ;
      RECT  1.885 0.63 1.975 0.76 ;
      RECT  1.85 0.76 1.975 0.9 ;
      RECT  1.85 0.9 2.15 0.99 ;
      RECT  2.06 0.99 2.15 1.06 ;
      RECT  2.06 1.06 2.34 1.165 ;
      RECT  3.585 0.445 3.87 0.565 ;
      RECT  3.78 0.565 3.87 0.885 ;
      RECT  3.78 0.885 4.28 0.975 ;
      RECT  4.12 0.975 4.28 1.13 ;
      RECT  4.12 1.13 4.21 1.285 ;
      RECT  3.64 1.285 4.21 1.375 ;
      RECT  3.64 1.375 3.76 1.61 ;
      RECT  4.325 0.17 4.445 0.695 ;
      RECT  4.0 0.695 4.47 0.79 ;
      RECT  4.0 0.79 4.86 0.795 ;
      RECT  4.38 0.795 4.86 0.89 ;
      RECT  4.38 0.89 4.47 1.255 ;
      RECT  4.3 1.255 4.47 1.36 ;
      RECT  2.43 1.05 2.925 1.14 ;
      RECT  2.835 1.14 2.925 1.25 ;
      RECT  2.43 1.14 2.52 1.255 ;
      RECT  2.835 1.25 3.48 1.34 ;
      RECT  3.385 0.415 3.48 1.25 ;
      RECT  1.68 0.51 1.785 0.605 ;
      RECT  1.635 0.605 1.785 0.685 ;
      RECT  1.635 0.685 1.725 1.08 ;
      RECT  1.635 1.08 1.97 1.2 ;
      RECT  1.88 1.2 1.97 1.255 ;
      RECT  1.88 1.255 2.52 1.345 ;
      RECT  3.37 1.34 3.48 1.61 ;
      RECT  0.895 1.29 1.79 1.39 ;
      RECT  1.7 1.39 1.79 1.46 ;
      RECT  1.7 1.46 2.08 1.58 ;
  END
END SEN_FSDPQ_DV1_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQ_DV1_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQ_DV1_4
  CLASS CORE ;
  FOREIGN SEN_FSDPQ_DV1_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.57 0.89 3.67 1.105 ;
      RECT  3.57 1.105 3.94 1.195 ;
      RECT  2.265 0.73 2.36 0.865 ;
      RECT  2.265 0.865 3.115 0.955 ;
      RECT  3.025 0.7 3.115 0.865 ;
      RECT  3.015 0.955 3.115 1.11 ;
      LAYER M2 ;
      RECT  2.93 0.95 3.71 1.05 ;
      LAYER V1 ;
      RECT  3.57 0.95 3.67 1.05 ;
      RECT  3.015 0.95 3.115 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.51 1.05 0.71 ;
      RECT  0.94 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.82 0.51 5.65 0.69 ;
      RECT  5.35 0.69 5.45 1.11 ;
      RECT  4.845 1.11 5.65 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.55 0.71 0.85 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.61 0.6 ;
      RECT  0.35 0.6 0.45 1.065 ;
      RECT  0.35 1.065 1.45 1.155 ;
      RECT  1.35 0.71 1.45 1.065 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.43 0.445 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  1.425 1.48 1.61 1.75 ;
      RECT  2.64 1.24 2.745 1.75 ;
      RECT  2.92 1.43 3.04 1.75 ;
      RECT  4.075 1.465 4.245 1.75 ;
      RECT  4.585 1.19 4.705 1.75 ;
      RECT  5.105 1.39 5.225 1.75 ;
      RECT  5.615 1.41 5.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  1.32 0.05 1.41 0.345 ;
      RECT  2.92 0.05 3.04 0.36 ;
      RECT  5.615 0.05 5.745 0.39 ;
      RECT  0.325 0.05 0.445 0.405 ;
      RECT  5.105 0.05 5.225 0.41 ;
      RECT  2.64 0.05 2.755 0.585 ;
      RECT  4.1 0.05 4.22 0.59 ;
      RECT  4.585 0.05 4.705 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.5 0.18 1.94 0.27 ;
      RECT  1.85 0.27 1.94 0.325 ;
      RECT  1.5 0.27 1.59 0.435 ;
      RECT  1.85 0.325 2.065 0.445 ;
      RECT  0.76 0.215 1.23 0.335 ;
      RECT  1.14 0.335 1.23 0.435 ;
      RECT  1.14 0.435 1.59 0.525 ;
      RECT  3.205 0.18 3.94 0.27 ;
      RECT  3.205 0.27 3.295 0.45 ;
      RECT  2.845 0.45 3.295 0.54 ;
      RECT  2.845 0.54 2.935 0.675 ;
      RECT  3.205 0.54 3.295 1.16 ;
      RECT  2.04 0.14 2.54 0.23 ;
      RECT  2.45 0.23 2.54 0.675 ;
      RECT  2.45 0.675 2.935 0.765 ;
      RECT  0.045 0.205 0.185 0.425 ;
      RECT  0.045 0.425 0.135 1.25 ;
      RECT  0.045 1.25 0.625 1.34 ;
      RECT  0.535 1.34 0.625 1.52 ;
      RECT  0.045 1.34 0.185 1.61 ;
      RECT  0.535 1.52 1.25 1.63 ;
      RECT  2.18 0.355 2.3 0.54 ;
      RECT  1.885 0.54 2.3 0.63 ;
      RECT  1.885 0.63 1.975 0.76 ;
      RECT  1.85 0.76 1.975 0.9 ;
      RECT  1.85 0.9 2.15 0.99 ;
      RECT  2.06 0.99 2.15 1.05 ;
      RECT  2.06 1.05 2.34 1.17 ;
      RECT  3.585 0.445 3.87 0.565 ;
      RECT  3.78 0.565 3.87 0.885 ;
      RECT  3.78 0.885 4.28 0.975 ;
      RECT  4.12 0.975 4.28 1.13 ;
      RECT  4.12 1.13 4.21 1.285 ;
      RECT  3.64 1.285 4.21 1.375 ;
      RECT  3.64 1.375 3.76 1.61 ;
      RECT  4.325 0.19 4.445 0.695 ;
      RECT  4.0 0.695 4.47 0.785 ;
      RECT  4.0 0.785 5.24 0.795 ;
      RECT  4.38 0.795 5.24 0.885 ;
      RECT  4.38 0.885 4.47 1.24 ;
      RECT  4.3 1.24 4.47 1.36 ;
      RECT  2.43 1.05 2.925 1.14 ;
      RECT  2.835 1.14 2.925 1.25 ;
      RECT  2.43 1.14 2.52 1.26 ;
      RECT  2.835 1.25 3.48 1.34 ;
      RECT  3.385 0.415 3.48 1.25 ;
      RECT  1.68 0.51 1.785 0.605 ;
      RECT  1.635 0.605 1.785 0.685 ;
      RECT  1.635 0.685 1.725 1.08 ;
      RECT  1.635 1.08 1.97 1.2 ;
      RECT  1.88 1.2 1.97 1.26 ;
      RECT  1.88 1.26 2.52 1.35 ;
      RECT  3.37 1.34 3.48 1.61 ;
      RECT  0.895 1.29 1.79 1.39 ;
      RECT  1.7 1.39 1.79 1.46 ;
      RECT  1.7 1.46 2.08 1.58 ;
  END
END SEN_FSDPQ_DV1_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQ_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDPQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.0 ;
      RECT  1.35 1.0 1.65 1.09 ;
      RECT  1.55 0.8 1.65 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.51 0.85 0.95 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.31 4.91 1.29 ;
    END
    ANTENNADIFFAREA 0.178 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.235 0.8 0.35 1.05 ;
      RECT  0.235 1.05 1.05 1.14 ;
      RECT  0.95 0.51 1.05 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.275 1.625 1.445 1.75 ;
      RECT  1.72 1.625 1.89 1.75 ;
      RECT  2.96 1.445 3.13 1.75 ;
      RECT  4.01 1.41 4.13 1.75 ;
      RECT  4.535 1.21 4.655 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  1.265 0.05 1.435 0.215 ;
      RECT  1.755 0.05 1.925 0.215 ;
      RECT  3.98 0.05 4.155 0.32 ;
      RECT  0.325 0.05 0.445 0.42 ;
      RECT  3.0 0.05 3.12 0.57 ;
      RECT  4.535 0.05 4.655 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.28 0.18 2.4 0.305 ;
      RECT  0.74 0.305 2.4 0.405 ;
      RECT  3.54 0.16 3.66 0.41 ;
      RECT  3.54 0.41 4.19 0.5 ;
      RECT  4.09 0.5 4.19 0.85 ;
      RECT  3.69 0.85 4.19 0.94 ;
      RECT  3.69 0.94 3.78 1.465 ;
      RECT  3.49 1.465 3.78 1.59 ;
      RECT  0.055 0.16 0.175 0.6 ;
      RECT  0.055 0.6 0.575 0.71 ;
      RECT  0.055 0.71 0.145 1.235 ;
      RECT  0.055 1.235 0.645 1.325 ;
      RECT  0.555 1.325 0.645 1.54 ;
      RECT  0.055 1.325 0.175 1.64 ;
      RECT  0.555 1.54 1.11 1.65 ;
      RECT  3.49 0.59 3.8 0.7 ;
      RECT  3.49 0.7 3.59 1.265 ;
      RECT  1.565 0.52 1.96 0.64 ;
      RECT  1.85 0.64 1.96 1.22 ;
      RECT  1.42 1.22 1.96 1.25 ;
      RECT  1.42 1.25 2.74 1.265 ;
      RECT  1.42 1.265 3.59 1.34 ;
      RECT  2.63 1.34 3.59 1.355 ;
      RECT  2.63 1.355 2.74 1.66 ;
      RECT  4.28 0.26 4.395 0.79 ;
      RECT  4.28 0.79 4.595 0.89 ;
      RECT  4.28 0.89 4.395 1.045 ;
      RECT  3.88 1.045 4.395 1.15 ;
      RECT  4.265 1.15 4.395 1.48 ;
      RECT  2.54 0.34 2.66 0.855 ;
      RECT  2.54 0.855 3.18 0.945 ;
      RECT  3.08 0.73 3.18 0.855 ;
      RECT  2.54 0.945 2.66 1.055 ;
      RECT  2.485 1.055 2.66 1.16 ;
      RECT  2.05 0.5 2.17 0.9 ;
      RECT  2.05 0.9 2.395 1.01 ;
      RECT  2.05 1.01 2.17 1.16 ;
      RECT  3.27 0.49 3.4 1.055 ;
      RECT  2.79 1.055 3.4 1.175 ;
      RECT  0.755 1.315 1.31 1.43 ;
      RECT  0.755 1.43 2.41 1.435 ;
      RECT  1.22 1.435 2.41 1.52 ;
  END
END SEN_FSDPQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQ_D_1P5
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQ_D_1P5
  CLASS CORE ;
  FOREIGN SEN_FSDPQ_D_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.18 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.3 5.255 1.5 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.235 0.65 0.475 ;
      RECT  0.405 0.475 0.65 0.595 ;
      RECT  0.55 0.595 0.65 1.08 ;
      RECT  0.55 1.08 1.46 1.17 ;
      RECT  1.365 1.0 1.46 1.08 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.4 1.44 0.52 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  1.59 1.63 1.76 1.75 ;
      RECT  1.91 1.63 2.08 1.75 ;
      RECT  3.29 1.48 3.46 1.75 ;
      RECT  4.38 1.21 4.5 1.75 ;
      RECT  4.89 1.19 5.01 1.75 ;
      RECT  5.415 1.21 5.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  1.945 0.05 2.115 0.2 ;
      RECT  1.24 0.05 1.41 0.36 ;
      RECT  0.325 0.05 0.445 0.375 ;
      RECT  4.34 0.05 4.48 0.39 ;
      RECT  5.41 0.05 5.54 0.39 ;
      RECT  4.89 0.05 5.01 0.565 ;
      RECT  3.25 0.05 3.37 0.57 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.81 0.215 4.17 0.335 ;
      RECT  4.08 0.335 4.17 0.71 ;
      RECT  4.08 0.71 4.59 0.72 ;
      RECT  4.05 0.72 4.59 0.8 ;
      RECT  4.5 0.8 4.59 0.94 ;
      RECT  4.05 0.8 4.14 1.48 ;
      RECT  3.83 1.48 4.14 1.595 ;
      RECT  3.52 0.19 3.72 0.36 ;
      RECT  3.63 0.36 3.72 1.08 ;
      RECT  3.165 0.855 3.255 1.08 ;
      RECT  3.165 1.08 3.72 1.21 ;
      RECT  1.5 0.3 2.69 0.42 ;
      RECT  1.5 0.42 1.59 0.45 ;
      RECT  0.795 0.165 0.915 0.45 ;
      RECT  0.795 0.45 1.59 0.54 ;
      RECT  4.64 0.245 4.77 0.465 ;
      RECT  4.68 0.465 4.77 0.77 ;
      RECT  4.68 0.77 5.06 0.94 ;
      RECT  4.68 0.94 4.77 1.03 ;
      RECT  4.23 0.89 4.32 1.03 ;
      RECT  4.23 1.03 4.77 1.12 ;
      RECT  4.64 1.12 4.77 1.41 ;
      RECT  1.68 0.51 2.08 0.61 ;
      RECT  1.99 0.61 2.08 0.795 ;
      RECT  1.99 0.795 2.25 0.965 ;
      RECT  1.99 0.965 2.08 1.27 ;
      RECT  1.67 1.27 2.08 1.36 ;
      RECT  3.82 0.48 3.99 0.65 ;
      RECT  3.82 0.65 3.91 1.3 ;
      RECT  3.055 1.3 3.91 1.39 ;
      RECT  3.055 1.39 3.145 1.565 ;
      RECT  2.61 0.67 2.7 0.855 ;
      RECT  2.61 0.855 2.76 0.945 ;
      RECT  2.67 0.945 2.76 1.565 ;
      RECT  2.67 1.565 3.145 1.66 ;
      RECT  2.79 0.39 2.9 0.675 ;
      RECT  2.79 0.675 3.51 0.765 ;
      RECT  3.42 0.765 3.51 0.985 ;
      RECT  2.85 0.765 2.94 1.465 ;
      RECT  2.2 0.56 2.52 0.68 ;
      RECT  2.43 0.68 2.52 1.1 ;
      RECT  2.22 1.1 2.52 1.19 ;
      RECT  2.22 1.19 2.34 1.35 ;
      RECT  0.065 0.165 0.185 1.26 ;
      RECT  0.065 1.26 0.805 1.35 ;
      RECT  0.715 1.35 0.805 1.545 ;
      RECT  0.065 1.35 0.185 1.63 ;
      RECT  0.715 1.545 1.275 1.66 ;
      RECT  0.895 1.305 1.465 1.425 ;
      RECT  1.365 1.425 1.465 1.45 ;
      RECT  1.365 1.45 2.58 1.54 ;
      RECT  2.475 1.28 2.58 1.45 ;
  END
END SEN_FSDPQ_D_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.0 ;
      RECT  1.35 1.0 1.65 1.09 ;
      RECT  1.55 0.8 1.65 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.51 0.85 0.95 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.31 4.86 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.235 0.8 0.35 1.05 ;
      RECT  0.235 1.05 1.05 1.14 ;
      RECT  0.95 0.51 1.05 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  1.275 1.625 1.445 1.75 ;
      RECT  1.72 1.625 1.89 1.75 ;
      RECT  2.96 1.445 3.13 1.75 ;
      RECT  4.005 1.41 4.135 1.75 ;
      RECT  4.48 1.41 4.61 1.75 ;
      RECT  5.015 1.21 5.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  1.265 0.05 1.435 0.215 ;
      RECT  1.755 0.05 1.925 0.215 ;
      RECT  3.98 0.05 4.155 0.32 ;
      RECT  4.48 0.05 4.61 0.39 ;
      RECT  0.32 0.05 0.45 0.4 ;
      RECT  2.995 0.05 3.125 0.57 ;
      RECT  5.015 0.05 5.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.28 0.18 2.4 0.305 ;
      RECT  0.74 0.305 2.4 0.405 ;
      RECT  3.54 0.17 3.66 0.41 ;
      RECT  3.54 0.41 4.19 0.5 ;
      RECT  4.09 0.5 4.19 0.79 ;
      RECT  3.69 0.79 4.19 0.88 ;
      RECT  3.69 0.88 3.78 1.465 ;
      RECT  3.5 1.465 3.78 1.59 ;
      RECT  0.055 0.17 0.175 0.6 ;
      RECT  0.055 0.6 0.605 0.71 ;
      RECT  0.055 0.71 0.145 1.235 ;
      RECT  0.055 1.235 0.645 1.325 ;
      RECT  0.555 1.325 0.645 1.54 ;
      RECT  0.055 1.325 0.175 1.63 ;
      RECT  0.555 1.54 1.1 1.65 ;
      RECT  3.49 0.59 3.82 0.7 ;
      RECT  3.49 0.7 3.59 1.265 ;
      RECT  1.55 0.52 1.96 0.64 ;
      RECT  1.85 0.64 1.96 1.22 ;
      RECT  1.42 1.22 1.96 1.25 ;
      RECT  1.42 1.25 2.74 1.265 ;
      RECT  1.42 1.265 3.59 1.34 ;
      RECT  2.63 1.34 3.59 1.355 ;
      RECT  2.63 1.355 2.74 1.66 ;
      RECT  4.28 0.39 4.39 0.785 ;
      RECT  4.28 0.785 4.64 0.895 ;
      RECT  4.28 0.895 4.39 0.985 ;
      RECT  3.87 0.985 4.39 1.09 ;
      RECT  4.27 1.09 4.39 1.35 ;
      RECT  2.54 0.34 2.66 0.855 ;
      RECT  2.54 0.855 3.18 0.945 ;
      RECT  3.08 0.775 3.18 0.855 ;
      RECT  2.54 0.945 2.66 1.055 ;
      RECT  2.485 1.055 2.66 1.16 ;
      RECT  2.05 0.5 2.17 0.9 ;
      RECT  2.05 0.9 2.395 1.01 ;
      RECT  2.05 1.01 2.17 1.16 ;
      RECT  3.27 0.49 3.4 1.055 ;
      RECT  2.83 1.055 3.4 1.175 ;
      RECT  0.75 1.315 1.31 1.43 ;
      RECT  0.75 1.43 2.41 1.435 ;
      RECT  1.22 1.435 2.41 1.52 ;
  END
END SEN_FSDPQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQ_D_3
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQ_D_3
  CLASS CORE ;
  FOREIGN SEN_FSDPQ_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.18 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.31 5.48 0.51 ;
      RECT  4.86 0.51 5.48 0.69 ;
      RECT  5.35 0.69 5.48 1.11 ;
      RECT  4.85 1.11 5.48 1.29 ;
    END
    ANTENNADIFFAREA 0.363 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.235 0.65 0.45 ;
      RECT  0.405 0.45 0.65 0.6 ;
      RECT  0.55 0.6 0.65 1.0 ;
      RECT  0.55 1.0 1.46 1.115 ;
      RECT  1.37 1.115 1.46 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.44 0.545 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  1.53 1.63 1.7 1.75 ;
      RECT  1.85 1.63 2.02 1.75 ;
      RECT  3.255 1.48 3.425 1.75 ;
      RECT  4.38 1.19 4.5 1.75 ;
      RECT  5.095 1.39 5.215 1.75 ;
      RECT  5.615 1.41 5.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  1.945 0.05 2.115 0.185 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  1.265 0.05 1.385 0.385 ;
      RECT  5.615 0.05 5.745 0.395 ;
      RECT  5.105 0.05 5.225 0.42 ;
      RECT  3.25 0.05 3.37 0.57 ;
      RECT  4.38 0.05 4.5 0.595 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.8 0.215 4.245 0.335 ;
      RECT  4.155 0.335 4.245 0.685 ;
      RECT  4.05 0.685 4.59 0.775 ;
      RECT  4.495 0.775 4.59 0.885 ;
      RECT  4.05 0.775 4.14 1.48 ;
      RECT  3.81 1.48 4.14 1.585 ;
      RECT  3.52 0.19 3.685 0.36 ;
      RECT  3.595 0.36 3.685 1.105 ;
      RECT  3.12 0.855 3.23 1.105 ;
      RECT  3.12 1.105 3.685 1.21 ;
      RECT  4.64 0.19 4.77 0.36 ;
      RECT  4.68 0.36 4.77 0.785 ;
      RECT  4.68 0.785 5.26 0.895 ;
      RECT  4.68 0.895 4.77 0.975 ;
      RECT  4.23 0.865 4.33 0.975 ;
      RECT  4.23 0.975 4.77 1.065 ;
      RECT  4.59 1.065 4.705 1.44 ;
      RECT  4.59 1.44 4.76 1.61 ;
      RECT  1.48 0.3 2.69 0.42 ;
      RECT  1.48 0.42 1.57 0.475 ;
      RECT  0.795 0.18 0.915 0.475 ;
      RECT  0.795 0.475 1.57 0.565 ;
      RECT  3.785 0.505 4.03 0.595 ;
      RECT  3.785 0.595 3.875 1.3 ;
      RECT  3.0 1.3 3.875 1.39 ;
      RECT  3.0 1.39 3.09 1.53 ;
      RECT  2.555 0.7 2.645 0.855 ;
      RECT  2.555 0.855 2.7 0.945 ;
      RECT  2.61 0.945 2.7 1.53 ;
      RECT  2.61 1.53 3.09 1.66 ;
      RECT  1.66 0.52 2.03 0.61 ;
      RECT  1.94 0.61 2.03 0.795 ;
      RECT  1.94 0.795 2.23 0.89 ;
      RECT  1.94 0.89 2.03 1.27 ;
      RECT  1.61 1.27 2.03 1.36 ;
      RECT  2.79 0.365 2.9 0.675 ;
      RECT  2.79 0.675 3.5 0.765 ;
      RECT  3.39 0.765 3.5 1.01 ;
      RECT  2.79 0.765 2.88 1.44 ;
      RECT  2.255 0.535 2.465 0.705 ;
      RECT  2.375 0.705 2.465 1.095 ;
      RECT  2.16 1.095 2.465 1.185 ;
      RECT  2.16 1.185 2.28 1.355 ;
      RECT  0.065 0.165 0.185 1.26 ;
      RECT  0.065 1.26 0.755 1.35 ;
      RECT  0.665 1.35 0.755 1.55 ;
      RECT  0.065 1.35 0.185 1.63 ;
      RECT  0.665 1.55 1.275 1.66 ;
      RECT  0.895 1.285 1.455 1.405 ;
      RECT  1.365 1.405 1.455 1.45 ;
      RECT  1.365 1.45 2.52 1.54 ;
      RECT  2.415 1.275 2.52 1.45 ;
  END
END SEN_FSDPQ_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQ_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDPQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.0 ;
      RECT  1.35 1.0 1.65 1.09 ;
      RECT  1.55 0.8 1.65 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.51 0.85 0.95 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.81 0.51 5.45 0.69 ;
      RECT  5.35 0.69 5.45 1.11 ;
      RECT  4.81 1.11 5.45 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.235 0.8 0.35 1.05 ;
      RECT  0.235 1.05 1.05 1.14 ;
      RECT  0.95 0.51 1.05 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  1.275 1.625 1.445 1.75 ;
      RECT  1.72 1.625 1.89 1.75 ;
      RECT  2.96 1.445 3.13 1.75 ;
      RECT  4.02 1.44 4.15 1.75 ;
      RECT  4.55 1.21 4.67 1.75 ;
      RECT  5.065 1.415 5.195 1.75 ;
      RECT  5.605 1.21 5.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  1.265 0.05 1.435 0.215 ;
      RECT  1.755 0.05 1.925 0.215 ;
      RECT  3.995 0.05 4.17 0.32 ;
      RECT  5.065 0.05 5.195 0.39 ;
      RECT  0.32 0.05 0.45 0.4 ;
      RECT  2.995 0.05 3.125 0.57 ;
      RECT  4.55 0.05 4.67 0.59 ;
      RECT  5.605 0.05 5.725 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.28 0.18 2.4 0.305 ;
      RECT  0.74 0.305 2.4 0.405 ;
      RECT  3.54 0.17 3.66 0.41 ;
      RECT  3.54 0.41 4.19 0.5 ;
      RECT  4.09 0.5 4.19 0.835 ;
      RECT  3.69 0.835 4.19 0.925 ;
      RECT  3.69 0.925 3.78 1.465 ;
      RECT  3.5 1.465 3.78 1.59 ;
      RECT  0.055 0.17 0.175 0.6 ;
      RECT  0.055 0.6 0.605 0.71 ;
      RECT  0.055 0.71 0.145 1.235 ;
      RECT  0.055 1.235 0.645 1.325 ;
      RECT  0.555 1.325 0.645 1.54 ;
      RECT  0.055 1.325 0.175 1.63 ;
      RECT  0.555 1.54 1.1 1.65 ;
      RECT  3.49 0.59 3.8 0.7 ;
      RECT  3.49 0.7 3.59 1.265 ;
      RECT  1.55 0.52 1.96 0.64 ;
      RECT  1.85 0.64 1.96 1.22 ;
      RECT  1.43 1.22 1.96 1.25 ;
      RECT  1.43 1.25 2.74 1.265 ;
      RECT  1.43 1.265 3.59 1.34 ;
      RECT  2.63 1.34 3.59 1.355 ;
      RECT  2.63 1.355 2.74 1.66 ;
      RECT  4.3 0.45 4.42 0.785 ;
      RECT  4.3 0.785 5.25 0.895 ;
      RECT  4.3 0.895 4.42 1.105 ;
      RECT  3.88 1.105 4.42 1.215 ;
      RECT  2.54 0.34 2.66 0.855 ;
      RECT  2.54 0.855 3.18 0.945 ;
      RECT  3.08 0.775 3.18 0.855 ;
      RECT  2.54 0.945 2.66 1.055 ;
      RECT  2.485 1.055 2.66 1.16 ;
      RECT  2.05 0.5 2.17 0.9 ;
      RECT  2.05 0.9 2.395 1.01 ;
      RECT  2.05 1.01 2.17 1.16 ;
      RECT  3.27 0.49 3.4 1.055 ;
      RECT  2.83 1.055 3.4 1.175 ;
      RECT  0.75 1.315 1.31 1.43 ;
      RECT  0.75 1.43 2.41 1.435 ;
      RECT  1.22 1.435 2.41 1.52 ;
  END
END SEN_FSDPQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_1
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.9 4.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.3 6.325 0.59 ;
      RECT  6.15 0.59 6.25 1.21 ;
      RECT  6.15 1.21 6.295 1.5 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.97 0.6 2.07 1.025 ;
      RECT  0.73 0.68 1.05 0.92 ;
      LAYER M2 ;
      RECT  0.86 0.75 2.11 0.85 ;
      LAYER V1 ;
      RECT  1.97 0.75 2.07 0.85 ;
      RECT  0.95 0.75 1.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.9 1.45 1.29 ;
      RECT  1.15 1.29 1.45 1.5 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.565 1.61 0.745 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  1.085 1.61 1.265 1.75 ;
      RECT  2.065 1.42 2.18 1.75 ;
      RECT  3.515 1.59 3.695 1.75 ;
      RECT  4.115 1.59 4.295 1.75 ;
      RECT  5.6 1.61 5.78 1.75 ;
      RECT  5.92 1.4 6.05 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  0.96 0.05 1.14 0.23 ;
      RECT  1.28 0.05 1.46 0.23 ;
      RECT  5.625 0.05 5.755 0.37 ;
      RECT  1.86 0.05 1.99 0.38 ;
      RECT  0.58 0.05 0.71 0.4 ;
      RECT  4.19 0.05 4.32 0.4 ;
      RECT  3.68 0.05 3.81 0.59 ;
      RECT  5.95 0.05 6.06 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.08 0.17 0.185 0.3 ;
      RECT  0.08 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 0.495 ;
      RECT  0.34 0.495 0.955 0.59 ;
      RECT  0.835 0.36 0.955 0.495 ;
      RECT  0.34 0.59 0.64 0.65 ;
      RECT  0.34 0.65 0.43 1.21 ;
      RECT  0.065 1.21 0.43 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  4.67 0.25 5.03 0.35 ;
      RECT  4.93 0.35 5.03 1.2 ;
      RECT  4.74 1.2 5.03 1.29 ;
      RECT  4.74 1.29 4.845 1.42 ;
      RECT  1.565 0.19 1.695 0.36 ;
      RECT  1.565 0.36 1.655 0.6 ;
      RECT  1.15 0.6 1.655 0.69 ;
      RECT  1.15 0.69 1.25 1.01 ;
      RECT  1.565 0.69 1.655 1.475 ;
      RECT  0.52 0.76 0.61 1.01 ;
      RECT  0.52 1.01 1.25 1.1 ;
      RECT  1.565 1.475 1.955 1.575 ;
      RECT  2.23 0.3 2.46 0.4 ;
      RECT  2.23 0.4 2.33 0.71 ;
      RECT  2.23 0.71 2.42 0.89 ;
      RECT  2.315 0.89 2.42 1.22 ;
      RECT  2.49 0.49 2.79 0.59 ;
      RECT  2.69 0.59 2.79 1.4 ;
      RECT  4.4 0.52 4.65 0.62 ;
      RECT  4.56 0.62 4.65 1.0 ;
      RECT  4.56 1.0 4.82 1.09 ;
      RECT  4.56 1.09 4.65 1.41 ;
      RECT  3.73 0.695 3.865 0.905 ;
      RECT  3.73 0.905 3.82 1.41 ;
      RECT  2.55 0.14 3.45 0.23 ;
      RECT  3.36 0.23 3.45 1.21 ;
      RECT  3.135 1.21 3.45 1.31 ;
      RECT  3.36 1.31 3.45 1.41 ;
      RECT  3.36 1.41 4.65 1.5 ;
      RECT  5.695 0.46 5.785 0.72 ;
      RECT  5.49 0.72 6.06 0.81 ;
      RECT  5.97 0.81 6.06 1.14 ;
      RECT  5.67 1.14 6.06 1.31 ;
      RECT  4.74 0.46 4.84 0.89 ;
      RECT  2.975 0.48 3.09 0.905 ;
      RECT  3.955 0.39 4.055 0.99 ;
      RECT  3.91 0.99 4.055 1.21 ;
      RECT  3.18 0.39 3.27 0.995 ;
      RECT  2.945 0.995 3.27 1.085 ;
      RECT  2.945 1.085 3.045 1.51 ;
      RECT  2.51 0.7 2.6 1.51 ;
      RECT  2.51 1.51 3.045 1.6 ;
      RECT  5.49 0.94 5.88 1.03 ;
      RECT  5.49 1.03 5.58 1.41 ;
      RECT  5.12 0.38 5.21 1.41 ;
      RECT  4.97 1.41 5.58 1.51 ;
      RECT  3.54 0.7 3.64 1.125 ;
      RECT  1.765 0.48 1.865 1.3 ;
      RECT  5.3 0.48 5.4 1.3 ;
      RECT  0.325 1.41 0.985 1.5 ;
      RECT  0.325 1.5 0.445 1.61 ;
      RECT  0.865 1.5 0.985 1.61 ;
      LAYER M2 ;
      RECT  0.42 0.55 2.83 0.65 ;
      RECT  2.95 0.55 5.5 0.65 ;
      RECT  2.23 0.75 5.11 0.85 ;
      LAYER V1 ;
      RECT  0.5 0.55 0.6 0.65 ;
      RECT  1.765 0.55 1.865 0.65 ;
      RECT  2.69 0.55 2.79 0.65 ;
      RECT  2.99 0.55 3.09 0.65 ;
      RECT  3.955 0.55 4.055 0.65 ;
      RECT  4.74 0.55 4.84 0.65 ;
      RECT  5.3 0.55 5.4 0.65 ;
      RECT  2.32 0.75 2.42 0.85 ;
      RECT  3.54 0.75 3.64 0.85 ;
      RECT  4.93 0.75 5.03 0.85 ;
  END
END SEN_FSDPQB_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_1P5
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_1P5
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.91 5.45 1.09 ;
      RECT  5.35 1.09 5.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0501 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 1.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0792 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.105 0.31 7.25 0.485 ;
      RECT  7.15 0.485 7.25 1.3 ;
      RECT  7.105 1.3 7.25 1.49 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.445 0.465 2.545 1.11 ;
      RECT  0.345 0.95 0.835 1.05 ;
      LAYER M2 ;
      RECT  0.455 0.95 2.585 1.05 ;
      LAYER V1 ;
      RECT  2.445 0.95 2.545 1.05 ;
      RECT  0.495 0.95 0.595 1.05 ;
      RECT  0.695 0.95 0.795 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0768 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 1.05 0.8 ;
      RECT  0.95 0.8 1.05 1.1 ;
      RECT  0.15 0.8 0.25 1.29 ;
      RECT  0.95 1.1 2.145 1.19 ;
      RECT  2.045 0.97 2.145 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.11 1.41 0.25 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  0.625 1.495 0.795 1.75 ;
      RECT  2.185 1.485 2.355 1.75 ;
      RECT  2.585 1.46 2.725 1.75 ;
      RECT  3.135 1.46 3.255 1.75 ;
      RECT  4.185 1.37 4.305 1.75 ;
      RECT  4.685 1.485 4.855 1.75 ;
      RECT  6.42 1.42 6.54 1.75 ;
      RECT  6.845 1.19 6.965 1.75 ;
      RECT  7.385 1.21 7.505 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  1.71 0.05 1.88 0.185 ;
      RECT  2.455 0.05 2.625 0.195 ;
      RECT  3.06 0.05 3.23 0.195 ;
      RECT  4.67 0.05 4.84 0.23 ;
      RECT  0.15 0.05 0.27 0.385 ;
      RECT  6.83 0.05 6.95 0.4 ;
      RECT  4.1 0.05 4.215 0.42 ;
      RECT  6.325 0.05 6.445 0.465 ;
      RECT  7.38 0.05 7.5 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.635 0.14 1.62 0.235 ;
      RECT  1.53 0.235 1.62 0.285 ;
      RECT  0.635 0.235 0.755 0.39 ;
      RECT  1.53 0.285 3.52 0.375 ;
      RECT  2.635 0.375 3.52 0.405 ;
      RECT  2.635 0.405 2.725 1.28 ;
      RECT  1.69 1.28 3.46 1.37 ;
      RECT  3.37 1.37 3.46 1.465 ;
      RECT  1.69 1.37 1.81 1.57 ;
      RECT  3.37 1.465 3.58 1.585 ;
      RECT  1.145 1.495 1.315 1.57 ;
      RECT  1.145 1.57 1.81 1.66 ;
      RECT  5.24 0.17 6.165 0.27 ;
      RECT  5.24 0.27 5.34 0.32 ;
      RECT  6.075 0.27 6.165 1.15 ;
      RECT  4.305 0.32 5.34 0.43 ;
      RECT  4.305 0.43 4.395 1.035 ;
      RECT  3.73 0.77 3.82 1.035 ;
      RECT  3.73 1.035 4.395 1.125 ;
      RECT  4.295 1.125 4.395 1.15 ;
      RECT  4.295 1.15 4.565 1.24 ;
      RECT  4.445 1.24 4.565 1.37 ;
      RECT  0.86 0.325 1.43 0.42 ;
      RECT  1.34 0.42 1.43 0.465 ;
      RECT  1.34 0.465 2.165 0.575 ;
      RECT  6.555 0.18 6.675 0.555 ;
      RECT  6.255 0.555 6.675 0.645 ;
      RECT  6.255 0.645 6.345 1.015 ;
      RECT  6.255 1.015 6.55 1.135 ;
      RECT  4.97 0.55 5.09 0.63 ;
      RECT  4.7 0.63 5.09 0.71 ;
      RECT  4.485 0.71 5.09 0.72 ;
      RECT  4.485 0.72 4.79 0.89 ;
      RECT  4.7 0.89 4.79 1.29 ;
      RECT  4.7 1.29 5.25 1.395 ;
      RECT  5.16 1.395 5.25 1.645 ;
      RECT  3.82 0.55 4.205 0.65 ;
      RECT  3.95 0.65 4.06 0.945 ;
      RECT  5.2 0.55 5.69 0.65 ;
      RECT  5.6 0.65 5.69 1.36 ;
      RECT  5.6 1.36 5.795 1.48 ;
      RECT  2.815 0.535 3.46 0.665 ;
      RECT  2.815 0.665 2.905 1.07 ;
      RECT  2.815 1.07 3.035 1.19 ;
      RECT  3.55 0.51 3.73 0.68 ;
      RECT  3.55 0.68 3.64 0.815 ;
      RECT  2.995 0.815 3.64 0.925 ;
      RECT  3.55 0.925 3.64 1.25 ;
      RECT  3.55 1.25 3.875 1.37 ;
      RECT  2.255 0.545 2.355 0.725 ;
      RECT  1.81 0.725 2.355 0.815 ;
      RECT  1.81 0.815 1.9 0.955 ;
      RECT  2.235 0.815 2.355 1.19 ;
      RECT  6.64 0.735 7.06 0.905 ;
      RECT  6.64 0.905 6.73 1.24 ;
      RECT  5.43 0.36 5.985 0.46 ;
      RECT  5.885 0.46 5.985 1.24 ;
      RECT  5.885 1.24 6.73 1.33 ;
      RECT  5.885 1.33 6.005 1.57 ;
      RECT  5.355 1.39 5.475 1.57 ;
      RECT  5.355 1.57 6.005 1.66 ;
      RECT  0.39 1.315 1.575 1.405 ;
      RECT  1.405 1.405 1.575 1.48 ;
      RECT  0.39 1.405 0.51 1.615 ;
      RECT  0.91 1.405 1.03 1.615 ;
      LAYER M2 ;
      RECT  3.08 0.55 5.58 0.65 ;
      LAYER V1 ;
      RECT  3.12 0.55 3.22 0.65 ;
      RECT  3.32 0.55 3.42 0.65 ;
      RECT  3.86 0.55 3.96 0.65 ;
      RECT  4.065 0.55 4.165 0.65 ;
      RECT  5.24 0.55 5.34 0.65 ;
      RECT  5.44 0.55 5.54 0.65 ;
  END
END SEN_FSDPQB_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_2
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.9 5.25 1.09 ;
      RECT  4.95 1.09 5.05 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0918 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.3 7.26 1.3 ;
    END
    ANTENNADIFFAREA 0.232 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.21 0.6 2.31 1.025 ;
      RECT  0.95 0.7 1.25 0.76 ;
      RECT  0.95 0.76 1.5 0.9 ;
      LAYER M2 ;
      RECT  0.84 0.75 2.4 0.85 ;
      LAYER V1 ;
      RECT  2.21 0.75 2.31 0.85 ;
      RECT  0.95 0.75 1.05 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.078 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 1.3 1.7 1.5 ;
      RECT  1.61 1.5 1.7 1.66 ;
      LAYER M2 ;
      RECT  1.28 1.35 1.92 1.45 ;
      LAYER V1 ;
      RECT  1.35 1.35 1.45 1.45 ;
      RECT  1.55 1.35 1.65 1.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.84 1.4 0.97 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  1.325 1.61 1.5 1.75 ;
      RECT  2.35 1.41 2.47 1.75 ;
      RECT  2.88 1.2 3.0 1.75 ;
      RECT  4.29 1.59 4.47 1.75 ;
      RECT  4.855 1.59 5.035 1.75 ;
      RECT  6.545 1.61 6.725 1.75 ;
      RECT  6.85 1.4 6.98 1.75 ;
      RECT  7.4 1.21 7.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  1.71 0.05 1.89 0.21 ;
      RECT  1.41 0.05 1.59 0.22 ;
      RECT  6.61 0.05 6.74 0.37 ;
      RECT  2.35 0.05 2.475 0.39 ;
      RECT  0.84 0.05 0.97 0.4 ;
      RECT  4.82 0.05 4.95 0.41 ;
      RECT  5.34 0.05 5.47 0.41 ;
      RECT  4.31 0.05 4.44 0.59 ;
      RECT  7.415 0.05 7.535 0.59 ;
      RECT  2.875 0.05 2.995 0.6 ;
      RECT  6.895 0.05 7.015 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.065 0.14 0.705 0.23 ;
      RECT  0.065 0.23 0.185 0.39 ;
      RECT  0.585 0.23 0.705 0.5 ;
      RECT  0.585 0.5 1.225 0.59 ;
      RECT  1.105 0.275 1.225 0.5 ;
      RECT  2.09 0.16 2.2 0.3 ;
      RECT  1.81 0.3 2.2 0.39 ;
      RECT  1.81 0.39 1.9 1.01 ;
      RECT  0.755 0.69 0.845 1.01 ;
      RECT  0.755 1.01 1.9 1.1 ;
      RECT  1.81 1.1 1.9 1.475 ;
      RECT  1.81 1.475 2.26 1.575 ;
      RECT  1.34 0.365 1.48 0.505 ;
      RECT  1.34 0.505 1.72 0.65 ;
      RECT  3.32 0.41 3.53 0.51 ;
      RECT  3.32 0.51 3.42 1.29 ;
      RECT  5.8 0.335 5.96 0.545 ;
      RECT  5.8 0.545 5.9 1.48 ;
      RECT  4.575 0.345 4.7 0.6 ;
      RECT  4.6 0.6 4.7 1.32 ;
      RECT  5.085 0.285 5.205 0.7 ;
      RECT  5.085 0.7 5.45 0.79 ;
      RECT  5.36 0.79 5.45 1.125 ;
      RECT  5.36 1.125 5.635 1.235 ;
      RECT  5.36 1.235 5.45 1.41 ;
      RECT  4.36 0.73 4.51 0.92 ;
      RECT  4.36 0.92 4.45 1.41 ;
      RECT  3.285 0.14 4.08 0.23 ;
      RECT  3.99 0.23 4.08 1.41 ;
      RECT  3.99 1.41 5.45 1.5 ;
      RECT  6.585 0.46 6.77 0.72 ;
      RECT  6.425 0.72 7.04 0.81 ;
      RECT  6.95 0.81 7.04 1.12 ;
      RECT  6.6 1.12 7.04 1.31 ;
      RECT  3.125 0.345 3.23 0.79 ;
      RECT  2.835 0.79 3.23 0.89 ;
      RECT  3.14 0.89 3.23 1.455 ;
      RECT  3.14 1.455 3.9 1.555 ;
      RECT  3.81 0.38 3.9 1.455 ;
      RECT  5.59 0.48 5.69 0.93 ;
      RECT  6.42 0.92 6.86 1.01 ;
      RECT  6.42 1.01 6.51 1.43 ;
      RECT  5.575 0.14 6.245 0.23 ;
      RECT  6.05 0.23 6.245 0.38 ;
      RECT  5.575 0.23 5.695 0.39 ;
      RECT  6.05 0.38 6.14 0.655 ;
      RECT  6.01 0.655 6.14 0.745 ;
      RECT  6.01 0.745 6.1 1.43 ;
      RECT  6.01 1.43 6.51 1.52 ;
      RECT  6.01 1.52 6.15 1.57 ;
      RECT  5.54 1.39 5.645 1.57 ;
      RECT  5.54 1.57 6.15 1.66 ;
      RECT  3.62 0.465 3.72 1.025 ;
      RECT  6.23 0.49 6.33 1.1 ;
      RECT  6.19 1.1 6.33 1.32 ;
      RECT  4.17 0.7 4.27 1.125 ;
      RECT  2.615 0.45 2.735 1.23 ;
      RECT  0.585 1.2 1.225 1.29 ;
      RECT  1.105 1.29 1.225 1.43 ;
      RECT  0.585 1.29 0.705 1.54 ;
      RECT  0.065 1.41 0.185 1.54 ;
      RECT  0.065 1.54 0.705 1.63 ;
      RECT  2.01 0.48 2.11 1.33 ;
      RECT  0.34 0.34 0.44 1.43 ;
      LAYER M2 ;
      RECT  0.195 0.55 3.46 0.65 ;
      RECT  3.58 0.55 6.4 0.65 ;
      RECT  2.555 0.75 6.0 0.85 ;
      LAYER V1 ;
      RECT  0.34 0.55 0.44 0.65 ;
      RECT  1.38 0.55 1.48 0.65 ;
      RECT  1.58 0.55 1.68 0.65 ;
      RECT  2.01 0.55 2.11 0.65 ;
      RECT  3.32 0.55 3.42 0.65 ;
      RECT  3.62 0.55 3.72 0.65 ;
      RECT  4.6 0.55 4.7 0.65 ;
      RECT  5.59 0.55 5.69 0.65 ;
      RECT  6.23 0.55 6.33 0.65 ;
      RECT  2.63 0.75 2.73 0.85 ;
      RECT  4.17 0.75 4.27 0.85 ;
      RECT  5.8 0.75 5.9 0.85 ;
  END
END SEN_FSDPQB_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_3
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_3
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.71 5.45 0.89 ;
      RECT  5.35 0.89 5.685 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0726 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.95 0.71 1.25 0.93 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1116 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.515 0.31 8.65 0.47 ;
      RECT  7.945 0.47 8.65 0.59 ;
      RECT  8.55 0.59 8.65 1.11 ;
      RECT  7.95 1.11 8.65 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.37 0.815 2.485 0.965 ;
      RECT  2.385 0.965 2.485 1.225 ;
      RECT  0.35 0.91 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.31 0.95 2.525 1.05 ;
      LAYER V1 ;
      RECT  2.385 0.95 2.485 1.05 ;
      RECT  0.35 0.95 0.45 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0999 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.85 0.8 ;
      RECT  0.15 0.8 0.25 0.89 ;
      RECT  0.75 0.8 0.85 1.055 ;
      RECT  0.75 1.055 2.095 1.145 ;
      RECT  2.005 1.145 2.095 1.225 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0345 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.35 0.19 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.565 1.495 0.735 1.75 ;
      RECT  2.145 1.495 2.315 1.75 ;
      RECT  2.58 1.495 2.75 1.75 ;
      RECT  3.1 1.495 3.27 1.75 ;
      RECT  4.655 1.425 4.775 1.75 ;
      RECT  5.21 1.48 5.38 1.75 ;
      RECT  5.83 1.48 5.95 1.75 ;
      RECT  7.345 1.475 7.515 1.75 ;
      RECT  7.735 1.19 7.855 1.75 ;
      RECT  8.255 1.405 8.375 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  2.41 0.05 2.58 0.17 ;
      RECT  2.98 0.05 3.15 0.17 ;
      RECT  1.63 0.05 1.8 0.175 ;
      RECT  5.06 0.05 5.23 0.2 ;
      RECT  5.6 0.05 5.77 0.2 ;
      RECT  8.255 0.05 8.375 0.38 ;
      RECT  0.07 0.05 0.21 0.39 ;
      RECT  4.565 0.05 4.695 0.42 ;
      RECT  7.235 0.05 7.355 0.485 ;
      RECT  7.735 0.05 7.855 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.55 0.14 1.54 0.23 ;
      RECT  1.445 0.23 1.54 0.265 ;
      RECT  0.55 0.23 0.67 0.395 ;
      RECT  1.445 0.265 3.96 0.37 ;
      RECT  1.445 0.37 2.53 0.385 ;
      RECT  3.79 0.37 3.96 0.42 ;
      RECT  2.44 0.385 2.53 0.635 ;
      RECT  2.44 0.635 2.665 0.725 ;
      RECT  2.575 0.725 2.665 1.305 ;
      RECT  2.575 1.305 3.56 1.315 ;
      RECT  1.645 1.315 3.56 1.405 ;
      RECT  3.47 1.405 3.56 1.48 ;
      RECT  1.645 1.405 1.765 1.495 ;
      RECT  3.47 1.48 4.075 1.6 ;
      RECT  1.06 1.495 1.765 1.6 ;
      RECT  5.905 0.155 7.095 0.265 ;
      RECT  5.905 0.265 5.995 0.29 ;
      RECT  7.005 0.265 7.095 1.165 ;
      RECT  4.785 0.29 5.995 0.38 ;
      RECT  4.825 0.38 4.915 1.11 ;
      RECT  4.085 1.03 4.175 1.11 ;
      RECT  4.085 1.11 4.915 1.2 ;
      RECT  4.825 1.2 4.915 1.26 ;
      RECT  4.825 1.26 5.025 1.35 ;
      RECT  4.915 1.35 5.025 1.6 ;
      RECT  0.76 0.32 1.3 0.42 ;
      RECT  1.205 0.42 1.3 0.475 ;
      RECT  1.205 0.475 2.085 0.595 ;
      RECT  3.555 0.46 3.675 0.51 ;
      RECT  3.555 0.51 4.245 0.64 ;
      RECT  3.555 0.64 3.675 0.805 ;
      RECT  2.945 0.805 3.74 0.915 ;
      RECT  3.65 0.915 3.74 1.29 ;
      RECT  3.65 1.29 4.285 1.39 ;
      RECT  4.165 1.39 4.285 1.51 ;
      RECT  2.695 0.46 3.175 0.55 ;
      RECT  2.755 0.55 3.465 0.565 ;
      RECT  3.085 0.565 3.465 0.65 ;
      RECT  2.755 0.565 2.845 1.07 ;
      RECT  2.755 1.07 3.53 1.19 ;
      RECT  7.465 0.165 7.585 0.575 ;
      RECT  7.185 0.575 7.585 0.695 ;
      RECT  7.185 0.695 7.44 0.745 ;
      RECT  7.335 0.745 7.44 1.16 ;
      RECT  5.115 0.47 5.5 0.59 ;
      RECT  5.115 0.59 5.205 0.895 ;
      RECT  5.005 0.895 5.205 1.065 ;
      RECT  5.115 1.065 5.205 1.285 ;
      RECT  5.115 1.285 6.16 1.39 ;
      RECT  6.065 1.39 6.16 1.545 ;
      RECT  6.065 1.545 6.775 1.66 ;
      RECT  5.615 0.55 6.62 0.65 ;
      RECT  6.53 0.65 6.62 1.06 ;
      RECT  6.53 1.06 6.715 1.165 ;
      RECT  4.435 0.51 4.735 0.69 ;
      RECT  4.47 0.69 4.57 1.0 ;
      RECT  2.175 0.52 2.28 0.825 ;
      RECT  1.66 0.825 2.28 0.935 ;
      RECT  2.185 0.935 2.28 1.015 ;
      RECT  2.185 1.015 2.295 1.2 ;
      RECT  7.53 0.785 8.385 0.895 ;
      RECT  7.53 0.895 7.635 1.255 ;
      RECT  6.085 0.355 6.895 0.46 ;
      RECT  6.805 0.46 6.895 1.255 ;
      RECT  6.295 1.165 6.415 1.255 ;
      RECT  6.295 1.255 7.635 1.385 ;
      RECT  0.28 1.285 1.515 1.405 ;
      LAYER M2 ;
      RECT  3.085 0.55 5.995 0.65 ;
      LAYER V1 ;
      RECT  3.125 0.55 3.225 0.65 ;
      RECT  3.325 0.55 3.425 0.65 ;
      RECT  4.435 0.55 4.535 0.65 ;
      RECT  4.635 0.55 4.735 0.65 ;
      RECT  5.655 0.55 5.755 0.65 ;
      RECT  5.855 0.55 5.955 0.65 ;
  END
END SEN_FSDPQB_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_4
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.7 5.45 0.9 ;
      RECT  5.35 0.9 5.85 1.1 ;
      LAYER M2 ;
      RECT  5.3 0.95 5.9 1.05 ;
      LAYER V1 ;
      RECT  5.45 0.95 5.55 1.05 ;
      RECT  5.65 0.95 5.75 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0756 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.51 8.45 0.69 ;
      RECT  8.35 0.69 8.45 1.11 ;
      RECT  7.75 1.11 8.45 1.29 ;
    END
    ANTENNADIFFAREA 0.46 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.26 0.6 2.36 1.19 ;
      RECT  0.95 0.7 1.325 0.92 ;
      LAYER M2 ;
      RECT  0.84 0.75 2.455 0.85 ;
      LAYER V1 ;
      RECT  2.26 0.75 2.36 0.85 ;
      RECT  0.95 0.75 1.05 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.099 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 1.3 1.74 1.5 ;
      RECT  1.65 1.5 1.74 1.66 ;
      LAYER M2 ;
      RECT  1.3 1.35 1.9 1.45 ;
      LAYER V1 ;
      RECT  1.395 1.35 1.495 1.45 ;
      RECT  1.595 1.35 1.695 1.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.845 1.4 0.965 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  1.345 1.61 1.525 1.75 ;
      RECT  2.415 1.41 2.545 1.75 ;
      RECT  2.94 1.21 3.06 1.75 ;
      RECT  3.46 1.21 3.58 1.75 ;
      RECT  4.81 1.48 4.99 1.75 ;
      RECT  5.33 1.48 5.51 1.75 ;
      RECT  5.84 1.48 6.02 1.75 ;
      RECT  7.195 1.61 7.375 1.75 ;
      RECT  7.51 1.41 7.64 1.75 ;
      RECT  8.04 1.41 8.17 1.75 ;
      RECT  8.6 1.21 8.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  1.745 0.05 1.925 0.21 ;
      RECT  1.425 0.05 1.605 0.23 ;
      RECT  7.16 0.05 7.29 0.37 ;
      RECT  2.35 0.05 2.48 0.39 ;
      RECT  8.035 0.05 8.165 0.39 ;
      RECT  0.84 0.05 0.97 0.41 ;
      RECT  4.84 0.05 4.97 0.59 ;
      RECT  8.6 0.05 8.72 0.59 ;
      RECT  2.875 0.05 2.995 0.6 ;
      RECT  3.395 0.05 3.515 0.6 ;
      RECT  5.355 0.05 5.475 0.6 ;
      RECT  5.875 0.05 5.995 0.6 ;
      RECT  7.48 0.05 7.6 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.065 0.14 0.705 0.23 ;
      RECT  0.065 0.23 0.185 0.39 ;
      RECT  0.585 0.23 0.705 0.5 ;
      RECT  0.585 0.5 1.225 0.59 ;
      RECT  1.105 0.37 1.225 0.5 ;
      RECT  2.095 0.16 2.215 0.3 ;
      RECT  1.85 0.3 2.215 0.39 ;
      RECT  1.85 0.39 1.94 1.01 ;
      RECT  0.75 0.69 0.84 1.01 ;
      RECT  0.75 1.01 1.94 1.1 ;
      RECT  1.85 1.1 1.94 1.525 ;
      RECT  1.85 1.525 2.285 1.635 ;
      RECT  2.16 1.42 2.285 1.525 ;
      RECT  1.37 0.365 1.475 0.5 ;
      RECT  1.37 0.5 1.72 0.6 ;
      RECT  1.42 0.6 1.72 0.7 ;
      RECT  5.09 0.38 5.23 0.6 ;
      RECT  5.13 0.6 5.23 0.99 ;
      RECT  5.1 0.99 5.23 1.19 ;
      RECT  7.075 0.555 7.35 0.655 ;
      RECT  7.075 0.655 7.175 1.025 ;
      RECT  7.075 1.025 7.41 1.125 ;
      RECT  3.84 0.4 4.01 0.7 ;
      RECT  3.91 0.7 4.01 1.28 ;
      RECT  3.91 1.28 4.14 1.38 ;
      RECT  5.615 0.44 5.735 0.7 ;
      RECT  5.615 0.7 6.03 0.79 ;
      RECT  5.94 0.79 6.03 1.035 ;
      RECT  5.94 1.035 6.095 1.27 ;
      RECT  5.94 1.27 6.03 1.28 ;
      RECT  4.92 0.715 5.04 0.92 ;
      RECT  4.92 0.92 5.01 1.28 ;
      RECT  3.845 0.14 4.6 0.23 ;
      RECT  4.51 0.23 4.6 1.28 ;
      RECT  4.51 1.28 6.03 1.37 ;
      RECT  5.61 1.37 5.725 1.51 ;
      RECT  2.615 0.46 2.735 0.71 ;
      RECT  2.615 0.71 3.335 0.89 ;
      RECT  3.135 0.46 3.255 0.71 ;
      RECT  2.68 0.89 2.8 1.23 ;
      RECT  3.2 0.89 3.32 1.23 ;
      RECT  3.66 0.44 3.75 0.755 ;
      RECT  3.445 0.755 3.75 0.795 ;
      RECT  3.445 0.795 3.815 0.925 ;
      RECT  3.725 0.925 3.815 1.47 ;
      RECT  3.725 1.47 4.42 1.57 ;
      RECT  4.33 0.5 4.42 1.47 ;
      RECT  7.52 0.79 8.24 0.89 ;
      RECT  7.52 0.89 7.62 1.23 ;
      RECT  7.075 1.23 7.62 1.32 ;
      RECT  7.075 1.32 7.165 1.41 ;
      RECT  6.125 0.14 6.75 0.23 ;
      RECT  6.125 0.23 6.245 0.41 ;
      RECT  6.655 0.23 6.75 1.41 ;
      RECT  6.655 1.41 7.165 1.5 ;
      RECT  6.655 1.5 6.75 1.57 ;
      RECT  6.12 1.36 6.24 1.57 ;
      RECT  6.12 1.57 6.75 1.66 ;
      RECT  6.14 0.5 6.24 0.93 ;
      RECT  4.69 0.685 4.81 1.05 ;
      RECT  6.84 0.48 6.94 1.115 ;
      RECT  6.84 1.115 6.985 1.32 ;
      RECT  4.14 0.475 4.24 1.125 ;
      RECT  0.585 1.2 1.225 1.29 ;
      RECT  1.105 1.29 1.225 1.42 ;
      RECT  0.585 1.29 0.705 1.54 ;
      RECT  0.065 1.41 0.185 1.54 ;
      RECT  0.065 1.54 0.705 1.63 ;
      RECT  2.05 0.48 2.15 1.32 ;
      RECT  0.34 0.44 0.44 1.41 ;
      RECT  6.39 0.44 6.5 1.46 ;
      LAYER M2 ;
      RECT  0.25 0.55 3.98 0.65 ;
      RECT  4.1 0.55 7.065 0.65 ;
      RECT  2.9 0.75 6.6 0.85 ;
      LAYER V1 ;
      RECT  0.34 0.55 0.44 0.65 ;
      RECT  1.42 0.55 1.52 0.65 ;
      RECT  1.62 0.55 1.72 0.65 ;
      RECT  2.05 0.55 2.15 0.65 ;
      RECT  3.84 0.55 3.94 0.65 ;
      RECT  4.14 0.55 4.24 0.65 ;
      RECT  5.13 0.55 5.23 0.65 ;
      RECT  6.14 0.55 6.24 0.65 ;
      RECT  6.84 0.55 6.94 0.65 ;
      RECT  3.035 0.75 3.135 0.85 ;
      RECT  3.235 0.75 3.335 0.85 ;
      RECT  4.69 0.75 4.79 0.85 ;
      RECT  6.395 0.75 6.495 0.85 ;
  END
END SEN_FSDPQB_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0417 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.31 5.06 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.235 0.65 0.43 ;
      RECT  0.435 0.43 0.65 0.6 ;
      RECT  0.55 0.6 0.65 1.01 ;
      RECT  0.55 1.01 1.425 1.1 ;
      RECT  1.335 1.1 1.425 1.195 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.38 1.44 0.52 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  1.41 1.615 1.58 1.75 ;
      RECT  1.92 1.615 2.09 1.75 ;
      RECT  3.335 1.44 3.455 1.75 ;
      RECT  4.375 1.465 4.545 1.75 ;
      RECT  4.695 1.44 4.815 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  1.98 0.05 2.15 0.17 ;
      RECT  0.29 0.05 0.46 0.34 ;
      RECT  1.3 0.05 1.42 0.36 ;
      RECT  4.375 0.05 4.495 0.385 ;
      RECT  3.335 0.05 3.455 0.425 ;
      RECT  4.695 0.05 4.815 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.51 0.26 2.745 0.35 ;
      RECT  1.51 0.35 1.6 0.45 ;
      RECT  0.785 0.19 0.91 0.45 ;
      RECT  0.785 0.45 1.6 0.54 ;
      RECT  3.84 0.24 4.275 0.36 ;
      RECT  4.185 0.36 4.275 1.26 ;
      RECT  4.045 1.26 4.725 1.35 ;
      RECT  4.635 0.725 4.725 1.26 ;
      RECT  4.045 1.35 4.135 1.465 ;
      RECT  3.85 1.465 4.135 1.585 ;
      RECT  2.28 0.44 2.57 0.545 ;
      RECT  2.47 0.545 2.57 1.095 ;
      RECT  2.215 1.095 2.57 1.185 ;
      RECT  2.215 1.185 2.335 1.345 ;
      RECT  1.69 0.465 2.085 0.585 ;
      RECT  1.995 0.585 2.085 0.73 ;
      RECT  1.995 0.73 2.36 0.84 ;
      RECT  1.995 0.84 2.085 1.255 ;
      RECT  1.63 1.255 2.085 1.345 ;
      RECT  2.84 0.19 2.955 0.675 ;
      RECT  2.84 0.675 3.52 0.765 ;
      RECT  3.43 0.765 3.52 0.98 ;
      RECT  2.84 0.765 2.945 1.44 ;
      RECT  4.435 0.475 4.545 0.76 ;
      RECT  4.365 0.76 4.545 0.93 ;
      RECT  4.435 0.93 4.545 1.17 ;
      RECT  3.8 0.485 3.9 0.905 ;
      RECT  4.005 0.475 4.095 1.0 ;
      RECT  3.84 1.0 4.095 1.09 ;
      RECT  3.84 1.09 3.93 1.26 ;
      RECT  3.07 1.26 3.93 1.35 ;
      RECT  3.07 1.35 3.16 1.565 ;
      RECT  2.66 0.67 2.75 1.565 ;
      RECT  2.66 1.565 3.16 1.66 ;
      RECT  3.185 0.855 3.275 1.08 ;
      RECT  3.185 1.08 3.71 1.17 ;
      RECT  3.61 0.27 3.71 1.08 ;
      RECT  0.055 0.185 0.175 1.26 ;
      RECT  0.055 1.26 0.835 1.35 ;
      RECT  0.745 1.35 0.835 1.555 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.745 1.555 1.245 1.66 ;
      RECT  0.925 1.285 1.425 1.405 ;
      RECT  1.335 1.405 1.425 1.435 ;
      RECT  1.335 1.435 2.57 1.525 ;
      RECT  2.465 1.275 2.57 1.435 ;
      LAYER M2 ;
      RECT  2.43 0.55 3.94 0.65 ;
      LAYER V1 ;
      RECT  2.47 0.55 2.57 0.65 ;
      RECT  3.8 0.55 3.9 0.65 ;
  END
END SEN_FSDPQB_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_D_1P5
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_D_1P5
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_D_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0417 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.3 5.06 0.51 ;
      RECT  4.95 0.51 5.25 0.6 ;
      RECT  5.15 0.6 5.25 1.11 ;
      RECT  4.93 1.11 5.25 1.29 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.235 0.65 0.43 ;
      RECT  0.435 0.43 0.65 0.6 ;
      RECT  0.55 0.6 0.65 1.01 ;
      RECT  0.55 1.01 1.425 1.1 ;
      RECT  1.335 1.1 1.425 1.195 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.38 1.44 0.52 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  1.41 1.615 1.58 1.75 ;
      RECT  1.91 1.615 2.08 1.75 ;
      RECT  3.325 1.44 3.445 1.75 ;
      RECT  4.355 1.465 4.525 1.75 ;
      RECT  4.685 1.44 4.805 1.75 ;
      RECT  5.205 1.41 5.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  1.97 0.05 2.14 0.17 ;
      RECT  0.29 0.05 0.46 0.34 ;
      RECT  1.29 0.05 1.41 0.36 ;
      RECT  4.365 0.05 4.485 0.385 ;
      RECT  5.205 0.05 5.34 0.39 ;
      RECT  3.325 0.05 3.445 0.57 ;
      RECT  4.695 0.05 4.815 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.5 0.26 2.735 0.35 ;
      RECT  1.5 0.35 1.59 0.45 ;
      RECT  0.785 0.19 0.905 0.45 ;
      RECT  0.785 0.45 1.59 0.54 ;
      RECT  2.27 0.44 2.56 0.545 ;
      RECT  2.46 0.545 2.56 1.095 ;
      RECT  2.205 1.095 2.56 1.185 ;
      RECT  2.205 1.185 2.325 1.345 ;
      RECT  1.68 0.465 2.075 0.585 ;
      RECT  1.985 0.585 2.075 0.73 ;
      RECT  1.985 0.73 2.34 0.84 ;
      RECT  1.985 0.84 2.075 1.255 ;
      RECT  1.615 1.255 2.075 1.345 ;
      RECT  2.83 0.19 2.945 0.675 ;
      RECT  2.83 0.675 3.51 0.765 ;
      RECT  3.42 0.765 3.51 0.93 ;
      RECT  2.83 0.765 2.935 1.465 ;
      RECT  4.425 0.475 4.535 0.755 ;
      RECT  4.355 0.755 4.535 0.925 ;
      RECT  4.425 0.925 4.535 1.17 ;
      RECT  4.635 0.775 5.055 0.895 ;
      RECT  4.635 0.895 4.725 1.26 ;
      RECT  3.83 0.24 4.265 0.36 ;
      RECT  4.175 0.36 4.265 1.26 ;
      RECT  4.035 1.26 4.725 1.35 ;
      RECT  4.035 1.35 4.125 1.465 ;
      RECT  3.84 1.465 4.125 1.585 ;
      RECT  3.79 0.485 3.89 0.93 ;
      RECT  3.995 0.475 4.085 1.025 ;
      RECT  3.83 1.025 4.085 1.115 ;
      RECT  3.83 1.115 3.92 1.26 ;
      RECT  3.06 1.26 3.92 1.35 ;
      RECT  3.06 1.35 3.15 1.565 ;
      RECT  2.65 0.67 2.74 1.565 ;
      RECT  2.65 1.565 3.15 1.66 ;
      RECT  3.175 0.855 3.265 1.08 ;
      RECT  3.175 1.08 3.7 1.17 ;
      RECT  3.6 0.27 3.7 1.08 ;
      RECT  0.055 0.165 0.175 1.26 ;
      RECT  0.055 1.26 0.82 1.35 ;
      RECT  0.73 1.35 0.82 1.555 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.73 1.555 1.25 1.66 ;
      RECT  0.91 1.29 1.43 1.405 ;
      RECT  1.34 1.405 1.43 1.435 ;
      RECT  1.34 1.435 2.56 1.525 ;
      RECT  2.455 1.29 2.56 1.435 ;
      LAYER M2 ;
      RECT  2.42 0.55 3.93 0.65 ;
      LAYER V1 ;
      RECT  2.46 0.55 2.56 0.65 ;
      RECT  3.79 0.55 3.89 0.65 ;
  END
END SEN_FSDPQB_D_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0417 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.905 0.455 5.25 0.575 ;
      RECT  5.15 0.575 5.25 1.11 ;
      RECT  4.95 1.11 5.25 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.235 0.65 0.43 ;
      RECT  0.435 0.43 0.65 0.6 ;
      RECT  0.55 0.6 0.65 1.03 ;
      RECT  0.55 1.03 1.425 1.12 ;
      RECT  1.335 1.025 1.425 1.03 ;
      RECT  1.335 1.12 1.425 1.195 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.38 1.44 0.52 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  1.41 1.615 1.58 1.75 ;
      RECT  1.92 1.615 2.09 1.75 ;
      RECT  3.335 1.44 3.455 1.75 ;
      RECT  4.375 1.455 4.545 1.75 ;
      RECT  4.695 1.44 4.815 1.75 ;
      RECT  5.205 1.41 5.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  1.98 0.05 2.15 0.17 ;
      RECT  0.29 0.05 0.46 0.34 ;
      RECT  1.3 0.05 1.42 0.36 ;
      RECT  5.215 0.05 5.335 0.365 ;
      RECT  4.385 0.05 4.505 0.385 ;
      RECT  3.335 0.05 3.455 0.585 ;
      RECT  4.695 0.05 4.815 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.51 0.26 2.745 0.35 ;
      RECT  1.51 0.35 1.6 0.45 ;
      RECT  0.785 0.19 0.905 0.45 ;
      RECT  0.785 0.45 1.6 0.54 ;
      RECT  2.28 0.44 2.57 0.545 ;
      RECT  2.47 0.545 2.57 1.095 ;
      RECT  2.215 1.095 2.57 1.185 ;
      RECT  2.215 1.185 2.335 1.315 ;
      RECT  1.69 0.465 2.085 0.585 ;
      RECT  1.995 0.585 2.085 0.73 ;
      RECT  1.995 0.73 2.35 0.84 ;
      RECT  1.995 0.84 2.085 1.255 ;
      RECT  1.625 1.255 2.085 1.345 ;
      RECT  2.84 0.19 2.955 0.675 ;
      RECT  2.84 0.675 3.52 0.765 ;
      RECT  3.43 0.765 3.52 0.93 ;
      RECT  2.84 0.765 2.945 1.44 ;
      RECT  4.425 0.475 4.545 0.755 ;
      RECT  4.365 0.755 4.545 0.925 ;
      RECT  4.425 0.925 4.545 1.17 ;
      RECT  4.635 0.785 5.055 0.895 ;
      RECT  4.635 0.895 4.725 1.26 ;
      RECT  3.84 0.24 4.275 0.36 ;
      RECT  4.185 0.36 4.275 1.26 ;
      RECT  4.045 1.26 4.725 1.35 ;
      RECT  4.045 1.35 4.135 1.465 ;
      RECT  3.85 1.465 4.135 1.585 ;
      RECT  3.8 0.485 3.9 0.93 ;
      RECT  4.005 0.475 4.095 1.025 ;
      RECT  3.84 1.025 4.095 1.115 ;
      RECT  3.84 1.115 3.93 1.26 ;
      RECT  3.07 1.26 3.93 1.35 ;
      RECT  3.07 1.35 3.16 1.565 ;
      RECT  2.66 0.67 2.75 1.565 ;
      RECT  2.66 1.565 3.16 1.66 ;
      RECT  3.185 0.855 3.275 1.08 ;
      RECT  3.185 1.08 3.71 1.17 ;
      RECT  3.61 0.27 3.71 1.08 ;
      RECT  0.055 0.165 0.175 1.26 ;
      RECT  0.055 1.26 0.82 1.35 ;
      RECT  0.73 1.35 0.82 1.555 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.73 1.555 1.25 1.66 ;
      RECT  0.91 1.285 1.43 1.405 ;
      RECT  1.34 1.405 1.43 1.435 ;
      RECT  1.34 1.435 2.57 1.525 ;
      RECT  2.465 1.29 2.57 1.435 ;
      LAYER M2 ;
      RECT  2.43 0.55 3.94 0.65 ;
      LAYER V1 ;
      RECT  2.47 0.55 2.57 0.65 ;
      RECT  3.8 0.55 3.9 0.65 ;
  END
END SEN_FSDPQB_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_D_3
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_D_3
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0417 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.51 5.65 0.69 ;
      RECT  5.55 0.69 5.65 1.11 ;
      RECT  4.95 1.11 5.65 1.29 ;
    END
    ANTENNADIFFAREA 0.391 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.235 0.65 0.43 ;
      RECT  0.435 0.43 0.65 0.6 ;
      RECT  0.55 0.6 0.65 1.0 ;
      RECT  0.55 1.0 1.435 1.09 ;
      RECT  1.345 1.09 1.435 1.18 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.38 1.44 0.52 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  1.42 1.615 1.59 1.75 ;
      RECT  1.93 1.615 2.1 1.75 ;
      RECT  3.345 1.44 3.465 1.75 ;
      RECT  4.385 1.465 4.555 1.75 ;
      RECT  4.735 1.44 4.855 1.75 ;
      RECT  5.255 1.415 5.375 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  1.99 0.05 2.16 0.17 ;
      RECT  0.29 0.05 0.46 0.34 ;
      RECT  1.31 0.05 1.43 0.36 ;
      RECT  4.395 0.05 4.515 0.385 ;
      RECT  5.245 0.05 5.385 0.41 ;
      RECT  3.345 0.05 3.465 0.585 ;
      RECT  4.735 0.05 4.855 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.52 0.26 2.755 0.35 ;
      RECT  1.52 0.35 1.61 0.45 ;
      RECT  0.785 0.19 0.905 0.45 ;
      RECT  0.785 0.45 1.61 0.54 ;
      RECT  2.29 0.44 2.58 0.545 ;
      RECT  2.48 0.545 2.58 1.095 ;
      RECT  2.225 1.095 2.58 1.185 ;
      RECT  2.225 1.185 2.345 1.315 ;
      RECT  1.7 0.465 2.095 0.585 ;
      RECT  2.005 0.585 2.095 0.73 ;
      RECT  2.005 0.73 2.36 0.84 ;
      RECT  2.005 0.84 2.095 1.255 ;
      RECT  1.635 1.255 2.095 1.345 ;
      RECT  2.85 0.19 2.965 0.675 ;
      RECT  2.85 0.675 3.53 0.765 ;
      RECT  3.44 0.765 3.53 0.93 ;
      RECT  2.85 0.765 2.955 1.44 ;
      RECT  4.465 0.475 4.575 0.755 ;
      RECT  4.375 0.755 4.575 0.925 ;
      RECT  4.465 0.925 4.575 1.17 ;
      RECT  4.75 0.785 5.44 0.895 ;
      RECT  4.75 0.895 4.84 1.26 ;
      RECT  3.85 0.24 4.285 0.36 ;
      RECT  4.195 0.36 4.285 1.26 ;
      RECT  4.055 1.26 4.84 1.35 ;
      RECT  4.055 1.35 4.145 1.465 ;
      RECT  3.86 1.465 4.145 1.585 ;
      RECT  3.8 0.485 3.9 0.93 ;
      RECT  4.015 0.475 4.105 1.025 ;
      RECT  3.85 1.025 4.105 1.115 ;
      RECT  3.85 1.115 3.94 1.26 ;
      RECT  3.08 1.26 3.94 1.35 ;
      RECT  3.08 1.35 3.17 1.565 ;
      RECT  2.67 0.67 2.76 1.565 ;
      RECT  2.67 1.565 3.17 1.66 ;
      RECT  3.195 0.855 3.285 1.08 ;
      RECT  3.195 1.08 3.75 1.17 ;
      RECT  3.62 0.27 3.71 1.08 ;
      RECT  0.055 0.19 0.175 1.26 ;
      RECT  0.055 1.26 0.845 1.35 ;
      RECT  0.755 1.35 0.845 1.555 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.755 1.555 1.27 1.66 ;
      RECT  0.935 1.285 1.45 1.405 ;
      RECT  1.36 1.405 1.45 1.435 ;
      RECT  1.36 1.435 2.58 1.525 ;
      RECT  2.475 1.29 2.58 1.435 ;
      LAYER M2 ;
      RECT  2.44 0.55 3.94 0.65 ;
      LAYER V1 ;
      RECT  2.48 0.55 2.58 0.65 ;
      RECT  3.8 0.55 3.9 0.65 ;
  END
END SEN_FSDPQB_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQB_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, qn-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):QN=iqn
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQB_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDPQB_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0417 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN QN
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.945 0.44 5.66 0.56 ;
      RECT  5.55 0.56 5.66 1.11 ;
      RECT  4.95 1.11 5.66 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END QN
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.235 0.65 0.465 ;
      RECT  0.395 0.465 0.65 0.565 ;
      RECT  0.55 0.565 0.65 1.03 ;
      RECT  0.55 1.03 1.435 1.12 ;
      RECT  1.345 1.025 1.435 1.03 ;
      RECT  1.345 1.12 1.435 1.195 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.38 1.44 0.52 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  1.42 1.615 1.59 1.75 ;
      RECT  1.93 1.615 2.1 1.75 ;
      RECT  3.345 1.44 3.465 1.75 ;
      RECT  4.395 1.465 4.565 1.75 ;
      RECT  4.735 1.44 4.855 1.75 ;
      RECT  5.255 1.39 5.375 1.75 ;
      RECT  5.79 1.21 5.91 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  1.99 0.05 2.16 0.17 ;
      RECT  0.29 0.05 0.46 0.34 ;
      RECT  5.255 0.05 5.375 0.35 ;
      RECT  1.255 0.05 1.375 0.36 ;
      RECT  4.385 0.05 4.505 0.385 ;
      RECT  4.735 0.05 4.855 0.565 ;
      RECT  3.345 0.05 3.465 0.585 ;
      RECT  5.79 0.05 5.91 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.49 0.26 2.755 0.35 ;
      RECT  1.49 0.35 1.58 0.45 ;
      RECT  0.785 0.19 0.905 0.45 ;
      RECT  0.785 0.45 1.58 0.54 ;
      RECT  2.29 0.44 2.58 0.545 ;
      RECT  2.48 0.545 2.58 1.095 ;
      RECT  2.225 1.095 2.58 1.185 ;
      RECT  2.225 1.185 2.345 1.315 ;
      RECT  1.7 0.465 2.095 0.585 ;
      RECT  2.005 0.585 2.095 0.73 ;
      RECT  2.005 0.73 2.36 0.84 ;
      RECT  2.005 0.84 2.095 1.255 ;
      RECT  1.635 1.255 2.095 1.345 ;
      RECT  2.85 0.19 2.965 0.675 ;
      RECT  2.85 0.675 3.53 0.765 ;
      RECT  3.44 0.765 3.53 0.93 ;
      RECT  2.85 0.765 2.955 1.465 ;
      RECT  4.455 0.475 4.575 0.755 ;
      RECT  4.375 0.755 4.575 0.925 ;
      RECT  4.455 0.925 4.575 1.17 ;
      RECT  4.75 0.785 5.42 0.895 ;
      RECT  4.75 0.895 4.84 1.26 ;
      RECT  3.85 0.24 4.285 0.36 ;
      RECT  4.195 0.36 4.285 1.26 ;
      RECT  4.055 1.26 4.84 1.35 ;
      RECT  4.055 1.35 4.145 1.465 ;
      RECT  3.86 1.465 4.145 1.585 ;
      RECT  3.8 0.485 3.9 0.93 ;
      RECT  4.015 0.475 4.105 1.025 ;
      RECT  3.85 1.025 4.105 1.115 ;
      RECT  3.85 1.115 3.94 1.26 ;
      RECT  3.08 1.26 3.94 1.35 ;
      RECT  3.08 1.35 3.17 1.565 ;
      RECT  2.67 0.67 2.76 1.565 ;
      RECT  2.67 1.565 3.17 1.66 ;
      RECT  3.195 0.855 3.285 1.08 ;
      RECT  3.195 1.08 3.71 1.17 ;
      RECT  3.62 0.27 3.71 1.08 ;
      RECT  0.055 0.19 0.175 1.26 ;
      RECT  0.055 1.26 0.845 1.35 ;
      RECT  0.755 1.35 0.845 1.555 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.755 1.555 1.27 1.66 ;
      RECT  0.935 1.285 1.45 1.405 ;
      RECT  1.36 1.405 1.45 1.435 ;
      RECT  1.36 1.435 2.58 1.525 ;
      RECT  2.475 1.29 2.58 1.435 ;
      LAYER M2 ;
      RECT  2.44 0.55 3.94 0.65 ;
      LAYER V1 ;
      RECT  2.48 0.55 2.58 0.65 ;
      RECT  3.8 0.55 3.9 0.65 ;
  END
END SEN_FSDPQB_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDPQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 4.45 0.75 ;
      RECT  4.25 0.75 4.45 0.91 ;
      RECT  4.25 0.91 4.85 0.92 ;
      RECT  4.35 0.92 4.85 1.105 ;
      RECT  3.045 0.69 3.145 0.82 ;
      RECT  3.045 0.82 3.785 0.99 ;
      LAYER M2 ;
      RECT  3.005 0.75 4.49 0.85 ;
      LAYER V1 ;
      RECT  4.35 0.75 4.45 0.85 ;
      RECT  3.045 0.75 3.145 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0765 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.85 0.845 ;
      RECT  0.75 0.845 1.17 0.945 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.31 6.45 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.29 0.69 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0714 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.99 ;
      RECT  1.35 0.99 1.575 1.07 ;
      RECT  0.45 0.495 0.65 0.595 ;
      RECT  0.55 0.595 0.65 1.07 ;
      RECT  0.55 1.07 1.575 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.815 0.415 5.935 1.02 ;
      RECT  5.75 1.02 5.935 1.11 ;
      RECT  5.75 1.11 5.85 1.49 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.44 1.43 0.58 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.635 1.51 1.755 1.75 ;
      RECT  3.015 1.515 3.185 1.75 ;
      RECT  3.845 1.415 3.965 1.75 ;
      RECT  5.135 1.6 5.305 1.75 ;
      RECT  5.425 1.6 5.595 1.75 ;
      RECT  5.995 1.215 6.115 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  4.965 0.05 5.135 0.23 ;
      RECT  5.52 0.05 5.69 0.23 ;
      RECT  2.965 0.05 3.135 0.31 ;
      RECT  1.475 0.05 1.58 0.36 ;
      RECT  0.385 0.05 0.505 0.405 ;
      RECT  3.845 0.05 3.965 0.405 ;
      RECT  6.065 0.05 6.19 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.245 0.155 4.68 0.245 ;
      RECT  4.245 0.245 4.335 0.35 ;
      RECT  4.09 0.35 4.335 0.45 ;
      RECT  1.67 0.18 2.31 0.27 ;
      RECT  1.67 0.27 1.76 0.45 ;
      RECT  2.19 0.27 2.31 0.48 ;
      RECT  0.955 0.19 1.075 0.45 ;
      RECT  0.955 0.45 1.76 0.54 ;
      RECT  1.67 0.54 1.76 1.25 ;
      RECT  1.035 1.25 1.76 1.33 ;
      RECT  1.035 1.33 2.13 1.42 ;
      RECT  2.04 1.42 2.13 1.495 ;
      RECT  2.04 1.495 2.34 1.625 ;
      RECT  3.325 0.275 3.445 0.4 ;
      RECT  2.865 0.4 3.445 0.49 ;
      RECT  2.865 0.49 2.955 0.705 ;
      RECT  2.58 0.705 2.955 0.875 ;
      RECT  2.865 0.875 2.955 1.155 ;
      RECT  2.865 1.155 3.47 1.245 ;
      RECT  3.3 1.09 3.47 1.155 ;
      RECT  2.4 0.24 2.57 0.41 ;
      RECT  2.4 0.41 2.49 0.78 ;
      RECT  2.1 0.78 2.49 0.95 ;
      RECT  2.4 0.95 2.49 1.055 ;
      RECT  2.4 1.055 2.545 1.225 ;
      RECT  4.72 0.33 5.66 0.42 ;
      RECT  4.72 0.42 4.84 0.55 ;
      RECT  5.57 0.42 5.66 0.755 ;
      RECT  5.57 0.755 5.72 0.925 ;
      RECT  5.57 0.925 5.66 1.42 ;
      RECT  4.825 1.42 5.66 1.51 ;
      RECT  3.59 0.29 3.74 0.59 ;
      RECT  3.235 0.59 3.965 0.7 ;
      RECT  3.875 0.7 3.965 1.12 ;
      RECT  3.57 1.12 3.965 1.29 ;
      RECT  5.12 0.51 5.445 0.62 ;
      RECT  5.12 0.62 5.22 0.975 ;
      RECT  5.12 0.975 5.285 1.145 ;
      RECT  4.065 0.54 4.285 0.645 ;
      RECT  4.065 0.645 4.155 1.24 ;
      RECT  4.065 1.24 4.475 1.35 ;
      RECT  4.355 1.35 4.475 1.46 ;
      RECT  5.35 0.71 5.465 0.89 ;
      RECT  5.375 0.89 5.465 1.24 ;
      RECT  4.425 0.4 4.63 0.52 ;
      RECT  4.54 0.52 4.63 0.72 ;
      RECT  4.54 0.72 5.03 0.81 ;
      RECT  4.94 0.81 5.03 1.24 ;
      RECT  4.615 1.24 5.465 1.33 ;
      RECT  4.615 1.33 4.735 1.6 ;
      RECT  1.85 0.36 2.01 1.1 ;
      RECT  1.85 1.1 2.31 1.19 ;
      RECT  2.22 1.19 2.31 1.315 ;
      RECT  2.22 1.315 2.695 1.335 ;
      RECT  2.22 1.335 3.49 1.405 ;
      RECT  2.635 1.405 3.49 1.425 ;
      RECT  3.4 1.425 3.49 1.545 ;
      RECT  2.825 1.425 2.915 1.59 ;
      RECT  3.4 1.545 3.65 1.655 ;
      RECT  6.045 0.53 6.15 1.125 ;
      RECT  0.065 0.19 0.185 1.25 ;
      RECT  0.065 1.25 0.945 1.34 ;
      RECT  0.855 1.34 0.945 1.54 ;
      RECT  0.065 1.34 0.185 1.61 ;
      RECT  0.855 1.54 1.34 1.65 ;
      LAYER M2 ;
      RECT  3.6 0.35 4.29 0.45 ;
      RECT  5.31 0.75 6.19 0.85 ;
      LAYER V1 ;
      RECT  3.64 0.35 3.74 0.45 ;
      RECT  4.15 0.35 4.25 0.45 ;
      RECT  5.35 0.75 5.45 0.85 ;
      RECT  6.05 0.75 6.15 0.85 ;
  END
END SEN_FSDPQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDPQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.51 6.65 0.725 ;
      RECT  6.44 0.725 6.65 0.895 ;
      RECT  5.67 0.71 5.955 0.9 ;
      RECT  4.825 0.715 5.09 0.895 ;
      LAYER M2 ;
      RECT  4.91 0.75 6.69 0.85 ;
      LAYER V1 ;
      RECT  6.55 0.75 6.65 0.85 ;
      RECT  5.75 0.75 5.85 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0987 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.335 0.71 2.45 0.855 ;
      RECT  2.35 0.855 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0816 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.05 0.31 8.17 0.45 ;
      RECT  8.05 0.45 8.45 0.54 ;
      RECT  8.35 0.54 8.45 1.05 ;
      RECT  8.05 1.05 8.45 1.14 ;
      RECT  8.05 1.14 8.17 1.25 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.5 0.71 0.65 1.025 ;
      RECT  0.5 1.025 0.795 1.115 ;
      RECT  0.705 1.115 0.795 1.225 ;
      RECT  0.705 1.225 1.6 1.33 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.084 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.615 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.28 0.29 7.4 0.445 ;
      RECT  7.28 0.445 7.45 0.535 ;
      RECT  7.35 0.535 7.45 1.045 ;
      RECT  7.25 1.045 7.45 1.165 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.625 0.5 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  1.44 1.42 1.56 1.75 ;
      RECT  2.465 1.46 2.635 1.75 ;
      RECT  3.945 1.495 4.115 1.75 ;
      RECT  4.515 1.495 4.685 1.75 ;
      RECT  5.31 1.605 5.48 1.75 ;
      RECT  6.97 1.62 7.14 1.75 ;
      RECT  7.705 1.625 7.875 1.75 ;
      RECT  8.33 1.23 8.45 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  5.31 0.05 5.48 0.185 ;
      RECT  1.925 0.05 2.095 0.195 ;
      RECT  8.335 0.05 8.455 0.36 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  3.99 0.05 4.11 0.41 ;
      RECT  7.79 0.05 7.91 0.415 ;
      RECT  6.995 0.05 7.115 0.455 ;
      RECT  2.71 0.05 2.83 0.465 ;
      RECT  4.54 0.05 4.66 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.65 0.14 1.58 0.23 ;
      RECT  0.65 0.23 0.77 0.505 ;
      RECT  0.65 0.505 0.975 0.595 ;
      RECT  0.885 0.595 0.975 0.96 ;
      RECT  0.885 0.96 2.1 1.05 ;
      RECT  0.885 1.05 1.055 1.135 ;
      RECT  2.01 1.05 2.1 1.25 ;
      RECT  2.01 1.25 3.325 1.37 ;
      RECT  3.22 0.195 3.325 1.25 ;
      RECT  2.01 1.37 2.1 1.465 ;
      RECT  1.915 1.465 2.1 1.585 ;
      RECT  2.465 0.19 2.555 0.32 ;
      RECT  0.86 0.32 2.555 0.415 ;
      RECT  6.565 0.26 6.85 0.38 ;
      RECT  6.75 0.38 6.85 0.725 ;
      RECT  6.75 0.725 7.24 0.835 ;
      RECT  6.75 0.835 6.85 1.01 ;
      RECT  6.63 1.01 6.85 1.13 ;
      RECT  0.32 0.19 0.45 0.41 ;
      RECT  0.32 0.41 0.41 1.15 ;
      RECT  0.22 1.15 0.41 1.25 ;
      RECT  5.03 0.275 5.815 0.445 ;
      RECT  5.695 0.445 5.815 0.45 ;
      RECT  5.695 0.45 6.135 0.54 ;
      RECT  6.045 0.54 6.135 1.29 ;
      RECT  5.605 1.29 6.27 1.38 ;
      RECT  5.605 1.38 5.71 1.395 ;
      RECT  6.1 1.38 6.27 1.415 ;
      RECT  5.015 1.395 5.71 1.515 ;
      RECT  4.8 0.165 4.92 0.535 ;
      RECT  4.8 0.535 5.505 0.625 ;
      RECT  5.415 0.625 5.505 1.02 ;
      RECT  5.415 1.02 5.945 1.12 ;
      RECT  5.415 1.12 5.515 1.165 ;
      RECT  4.8 1.165 5.515 1.255 ;
      RECT  4.8 1.255 4.92 1.315 ;
      RECT  3.61 1.18 3.7 1.315 ;
      RECT  3.61 1.315 4.92 1.405 ;
      RECT  4.8 1.405 4.92 1.495 ;
      RECT  3.61 1.405 3.7 1.52 ;
      RECT  2.725 1.52 3.7 1.63 ;
      RECT  3.76 0.505 4.43 0.61 ;
      RECT  4.33 0.61 4.43 0.985 ;
      RECT  4.33 0.985 5.325 1.075 ;
      RECT  5.225 0.73 5.325 0.985 ;
      RECT  4.33 1.075 4.43 1.12 ;
      RECT  4.2 1.12 4.43 1.225 ;
      RECT  1.09 0.515 2.39 0.62 ;
      RECT  3.48 0.19 3.6 0.735 ;
      RECT  3.48 0.735 4.215 0.82 ;
      RECT  3.415 0.82 4.215 0.905 ;
      RECT  3.415 0.905 3.52 1.26 ;
      RECT  7.73 0.785 8.21 0.895 ;
      RECT  7.73 0.895 7.82 1.44 ;
      RECT  5.955 0.19 6.46 0.36 ;
      RECT  6.26 0.36 6.46 0.405 ;
      RECT  6.26 0.405 6.35 0.985 ;
      RECT  6.26 0.985 6.54 1.155 ;
      RECT  6.425 1.155 6.54 1.44 ;
      RECT  6.425 1.44 7.82 1.53 ;
      RECT  6.425 1.53 6.54 1.555 ;
      RECT  5.84 1.47 6.01 1.555 ;
      RECT  5.84 1.555 6.54 1.66 ;
      RECT  2.97 0.24 3.085 1.03 ;
      RECT  2.75 1.03 3.085 1.15 ;
      RECT  7.54 0.19 7.64 1.255 ;
      RECT  6.76 1.255 7.64 1.35 ;
      RECT  1.71 1.15 1.92 1.295 ;
      RECT  1.71 1.295 1.82 1.62 ;
      RECT  0.07 1.335 0.19 1.435 ;
      RECT  0.07 1.435 1.325 1.535 ;
      RECT  1.155 1.535 1.325 1.58 ;
      LAYER M2 ;
      RECT  0.22 1.15 1.89 1.25 ;
      LAYER V1 ;
      RECT  0.26 1.15 0.36 1.25 ;
      RECT  1.75 1.15 1.85 1.25 ;
  END
END SEN_FSDPQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDPQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.91 0.63 7.09 0.89 ;
      RECT  6.115 0.66 6.255 0.75 ;
      RECT  5.97 0.75 6.255 0.9 ;
      RECT  4.75 0.66 4.855 0.75 ;
      RECT  4.75 0.75 5.19 0.85 ;
      RECT  4.75 0.85 4.855 0.89 ;
      LAYER M2 ;
      RECT  5.01 0.75 7.09 0.85 ;
      LAYER V1 ;
      RECT  6.95 0.75 7.05 0.85 ;
      RECT  6.125 0.75 6.225 0.85 ;
      RECT  5.05 0.75 5.15 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1275 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.45 0.75 ;
      RECT  1.405 0.75 2.45 0.855 ;
      RECT  2.35 0.855 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.35 0.31 8.48 0.475 ;
      RECT  8.35 0.475 9.05 0.595 ;
      RECT  8.95 0.595 9.05 1.11 ;
      RECT  8.33 1.11 9.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.675 0.52 1.25 ;
      RECT  0.35 1.25 1.585 1.36 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0993 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.555 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.55 0.29 7.715 0.51 ;
      RECT  7.55 0.51 7.85 0.615 ;
      RECT  7.65 0.615 7.85 0.89 ;
      RECT  7.65 0.89 7.74 0.97 ;
      RECT  7.57 0.97 7.74 1.075 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.63 0.5 1.75 ;
      RECT  0.0 1.75 9.4 1.85 ;
      RECT  1.415 1.45 1.585 1.75 ;
      RECT  2.485 1.39 2.59 1.75 ;
      RECT  4.055 1.445 4.175 1.75 ;
      RECT  4.595 1.445 4.715 1.75 ;
      RECT  5.135 1.395 5.255 1.75 ;
      RECT  5.68 1.575 5.795 1.75 ;
      RECT  7.285 1.62 7.455 1.75 ;
      RECT  8.055 1.525 8.175 1.75 ;
      RECT  8.635 1.39 8.755 1.75 ;
      RECT  9.18 1.21 9.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      RECT  1.905 0.05 2.075 0.19 ;
      RECT  5.68 0.05 5.85 0.31 ;
      RECT  4.04 0.05 4.21 0.325 ;
      RECT  5.135 0.05 5.255 0.36 ;
      RECT  7.315 0.05 7.435 0.37 ;
      RECT  8.635 0.05 8.755 0.385 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  2.795 0.05 2.915 0.41 ;
      RECT  4.595 0.05 4.715 0.57 ;
      RECT  9.18 0.05 9.3 0.59 ;
      RECT  8.12 0.05 8.23 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.61 0.15 1.545 0.26 ;
      RECT  0.61 0.26 0.715 0.945 ;
      RECT  0.61 0.945 2.13 1.035 ;
      RECT  0.885 1.035 1.055 1.16 ;
      RECT  2.04 1.035 2.13 1.21 ;
      RECT  2.04 1.21 3.425 1.3 ;
      RECT  3.32 0.39 3.425 1.21 ;
      RECT  2.04 1.3 2.13 1.475 ;
      RECT  1.93 1.475 2.13 1.6 ;
      RECT  7.805 0.215 8.03 0.335 ;
      RECT  7.94 0.335 8.03 1.015 ;
      RECT  7.86 1.015 8.03 1.165 ;
      RECT  7.36 1.165 8.03 1.255 ;
      RECT  7.36 1.255 7.45 1.26 ;
      RECT  7.095 1.26 7.45 1.35 ;
      RECT  2.535 0.22 2.655 0.35 ;
      RECT  0.805 0.35 2.655 0.44 ;
      RECT  3.53 0.24 3.735 0.36 ;
      RECT  3.53 0.36 3.62 0.715 ;
      RECT  3.53 0.715 4.315 0.885 ;
      RECT  3.53 0.885 3.62 1.39 ;
      RECT  2.925 1.39 3.62 1.48 ;
      RECT  6.485 0.32 6.605 0.4 ;
      RECT  5.46 0.4 6.605 0.5 ;
      RECT  5.46 0.5 5.565 0.62 ;
      RECT  6.4 0.5 6.49 1.285 ;
      RECT  5.965 1.285 6.64 1.375 ;
      RECT  5.965 1.375 6.085 1.395 ;
      RECT  6.47 1.375 6.64 1.405 ;
      RECT  5.395 1.395 6.085 1.485 ;
      RECT  5.395 1.485 5.515 1.615 ;
      RECT  7.025 0.21 7.145 0.45 ;
      RECT  7.025 0.45 7.27 0.54 ;
      RECT  7.18 0.54 7.27 0.705 ;
      RECT  7.18 0.705 7.535 0.805 ;
      RECT  7.18 0.805 7.27 0.99 ;
      RECT  7.04 0.99 7.27 1.16 ;
      RECT  0.33 0.19 0.45 0.485 ;
      RECT  0.15 0.485 0.45 0.575 ;
      RECT  0.15 0.575 0.25 1.29 ;
      RECT  3.875 0.415 4.495 0.535 ;
      RECT  3.875 0.535 4.045 0.625 ;
      RECT  4.405 0.535 4.495 1.005 ;
      RECT  4.3 1.005 4.495 1.01 ;
      RECT  4.3 1.01 5.105 1.1 ;
      RECT  4.935 0.97 5.105 1.01 ;
      RECT  4.3 1.1 4.47 1.135 ;
      RECT  4.825 0.45 5.37 0.57 ;
      RECT  5.28 0.57 5.37 0.99 ;
      RECT  5.28 0.99 6.305 1.1 ;
      RECT  5.28 1.1 5.37 1.215 ;
      RECT  4.955 1.215 5.37 1.225 ;
      RECT  3.735 1.185 3.825 1.225 ;
      RECT  3.735 1.225 5.37 1.305 ;
      RECT  3.735 1.305 5.0 1.355 ;
      RECT  3.735 1.355 3.825 1.57 ;
      RECT  2.68 1.57 3.825 1.66 ;
      RECT  1.055 0.53 2.36 0.62 ;
      RECT  8.12 0.79 8.84 0.9 ;
      RECT  8.12 0.9 8.21 1.345 ;
      RECT  7.54 1.345 8.21 1.435 ;
      RECT  7.54 1.435 7.63 1.44 ;
      RECT  6.2 0.14 6.885 0.23 ;
      RECT  6.2 0.23 6.37 0.31 ;
      RECT  6.73 0.23 6.885 0.36 ;
      RECT  6.73 0.36 6.82 1.0 ;
      RECT  6.73 1.0 6.87 1.17 ;
      RECT  6.77 1.17 6.87 1.44 ;
      RECT  6.77 1.44 7.63 1.53 ;
      RECT  6.21 1.465 6.38 1.53 ;
      RECT  6.21 1.53 6.875 1.62 ;
      RECT  3.055 0.27 3.16 1.015 ;
      RECT  3.055 1.015 3.225 1.03 ;
      RECT  2.77 1.03 3.225 1.12 ;
      RECT  1.715 1.15 1.95 1.265 ;
      RECT  1.715 1.265 1.83 1.62 ;
      RECT  0.07 1.38 0.19 1.45 ;
      RECT  0.07 1.45 1.325 1.54 ;
      RECT  1.155 1.54 1.325 1.58 ;
      RECT  0.07 1.54 0.185 1.6 ;
      LAYER M2 ;
      RECT  0.11 1.15 1.895 1.25 ;
      LAYER V1 ;
      RECT  0.15 1.15 0.25 1.25 ;
      RECT  1.755 1.15 1.855 1.25 ;
  END
END SEN_FSDPQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQO_6
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQO_6
  CLASS CORE ;
  FOREIGN SEN_FSDPQO_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.145 0.69 8.25 1.21 ;
      RECT  8.145 1.21 8.335 1.345 ;
      RECT  7.42 0.7 7.66 0.745 ;
      RECT  7.42 0.745 7.8 0.85 ;
      RECT  5.485 0.75 5.865 0.92 ;
      LAYER M2 ;
      RECT  5.485 0.75 8.29 0.85 ;
      LAYER V1 ;
      RECT  8.15 0.75 8.25 0.85 ;
      RECT  7.66 0.75 7.76 0.85 ;
      RECT  5.525 0.75 5.625 0.85 ;
      RECT  5.725 0.75 5.825 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1488 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.91 0.71 1.45 0.955 ;
      LAYER M2 ;
      RECT  0.425 0.75 1.29 0.85 ;
      LAYER V1 ;
      RECT  0.95 0.75 1.05 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.845 0.51 11.05 0.69 ;
      RECT  10.72 0.69 10.85 1.11 ;
      RECT  9.75 1.11 11.05 1.29 ;
    END
    ANTENNADIFFAREA 0.656 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.45 2.51 0.905 ;
      RECT  0.42 0.55 0.66 0.65 ;
      RECT  0.51 0.65 0.66 0.89 ;
      LAYER M2 ;
      RECT  0.42 0.55 2.55 0.65 ;
      LAYER V1 ;
      RECT  2.41 0.55 2.51 0.65 ;
      RECT  0.46 0.55 0.56 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1116 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.065 ;
      RECT  0.15 1.065 2.095 1.155 ;
      RECT  2.005 0.985 2.095 1.065 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.95 0.51 9.09 1.325 ;
    END
    ANTENNADIFFAREA 0.151 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.39 0.185 1.75 ;
      RECT  0.0 1.75 11.4 1.85 ;
      RECT  0.56 1.48 0.73 1.75 ;
      RECT  2.095 1.44 2.215 1.75 ;
      RECT  2.595 1.44 2.715 1.75 ;
      RECT  3.12 1.44 3.24 1.75 ;
      RECT  4.78 1.54 4.905 1.75 ;
      RECT  5.28 1.525 5.45 1.75 ;
      RECT  5.835 1.495 6.005 1.75 ;
      RECT  6.365 1.44 6.51 1.75 ;
      RECT  6.885 1.44 7.035 1.75 ;
      RECT  8.665 1.615 8.835 1.75 ;
      RECT  9.535 1.44 9.655 1.75 ;
      RECT  10.055 1.39 10.175 1.75 ;
      RECT  10.61 1.39 10.73 1.75 ;
      RECT  11.18 1.21 11.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.4 0.05 ;
      RECT  1.64 0.05 1.81 0.17 ;
      RECT  2.475 0.05 2.645 0.17 ;
      RECT  3.045 0.05 3.215 0.17 ;
      RECT  4.745 0.05 4.915 0.185 ;
      RECT  8.665 0.05 8.835 0.22 ;
      RECT  6.355 0.05 6.525 0.32 ;
      RECT  6.875 0.05 7.045 0.32 ;
      RECT  0.1 0.05 0.24 0.39 ;
      RECT  5.33 0.05 5.45 0.41 ;
      RECT  10.105 0.05 10.225 0.41 ;
      RECT  10.625 0.05 10.745 0.41 ;
      RECT  11.18 0.05 11.3 0.59 ;
      RECT  9.585 0.05 9.705 0.61 ;
      RECT  5.855 0.05 5.975 0.615 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.42 0.165 4.03 0.26 ;
      RECT  0.55 0.26 4.03 0.28 ;
      RECT  0.55 0.28 3.51 0.36 ;
      RECT  2.6 0.36 3.51 0.365 ;
      RECT  2.6 0.365 2.71 1.26 ;
      RECT  1.625 1.26 3.42 1.35 ;
      RECT  1.625 1.35 1.745 1.48 ;
      RECT  3.33 1.35 3.42 1.54 ;
      RECT  1.055 1.48 1.745 1.6 ;
      RECT  3.33 1.54 4.12 1.66 ;
      RECT  8.405 0.14 8.575 0.31 ;
      RECT  8.405 0.31 9.37 0.4 ;
      RECT  9.25 0.165 9.37 0.31 ;
      RECT  9.265 0.4 9.37 1.17 ;
      RECT  4.335 0.275 5.225 0.365 ;
      RECT  4.785 0.365 5.225 0.395 ;
      RECT  4.335 0.365 4.425 0.685 ;
      RECT  4.785 0.395 4.875 1.07 ;
      RECT  4.205 0.685 4.425 0.795 ;
      RECT  4.785 1.07 5.2 1.185 ;
      RECT  7.665 0.355 7.835 0.41 ;
      RECT  6.07 0.41 7.835 0.53 ;
      RECT  6.81 0.53 6.9 1.23 ;
      RECT  6.135 1.13 6.24 1.23 ;
      RECT  6.135 1.23 7.825 1.35 ;
      RECT  3.6 0.39 4.245 0.48 ;
      RECT  4.135 0.48 4.245 0.56 ;
      RECT  3.6 0.48 3.705 0.76 ;
      RECT  3.6 0.76 3.78 0.79 ;
      RECT  2.985 0.79 3.78 0.9 ;
      RECT  3.69 0.9 3.78 1.165 ;
      RECT  3.69 1.165 4.385 1.27 ;
      RECT  0.81 0.465 2.12 0.585 ;
      RECT  5.3 0.54 5.735 0.66 ;
      RECT  5.3 0.66 5.395 0.805 ;
      RECT  4.965 0.805 5.395 0.925 ;
      RECT  5.295 0.925 5.395 1.08 ;
      RECT  5.295 1.08 5.745 1.2 ;
      RECT  8.395 0.49 8.555 0.66 ;
      RECT  8.465 0.66 8.555 1.025 ;
      RECT  8.385 1.025 8.555 1.045 ;
      RECT  8.385 1.045 8.86 1.135 ;
      RECT  8.755 0.735 8.86 1.045 ;
      RECT  2.215 0.535 2.32 0.8 ;
      RECT  1.745 0.8 2.32 0.89 ;
      RECT  1.745 0.89 1.835 0.97 ;
      RECT  2.23 0.89 2.32 1.025 ;
      RECT  2.23 1.025 2.495 1.145 ;
      RECT  3.905 0.69 4.075 0.8 ;
      RECT  3.985 0.8 4.075 0.95 ;
      RECT  3.985 0.95 4.49 1.05 ;
      RECT  9.46 0.78 10.61 0.895 ;
      RECT  9.46 0.895 9.55 1.26 ;
      RECT  9.355 1.26 9.55 1.35 ;
      RECT  9.355 1.35 9.445 1.435 ;
      RECT  7.405 0.175 8.055 0.265 ;
      RECT  7.405 0.265 7.575 0.32 ;
      RECT  7.95 0.265 8.055 0.675 ;
      RECT  7.915 0.675 8.055 0.78 ;
      RECT  7.915 0.78 8.005 1.435 ;
      RECT  7.915 1.435 9.445 1.44 ;
      RECT  7.37 1.44 9.445 1.525 ;
      RECT  7.37 1.525 8.135 1.56 ;
      RECT  5.955 0.795 6.67 0.91 ;
      RECT  5.955 0.91 6.045 1.315 ;
      RECT  4.605 0.57 4.695 1.315 ;
      RECT  4.605 1.315 6.045 1.36 ;
      RECT  2.8 0.48 3.51 0.6 ;
      RECT  2.8 0.6 2.89 1.025 ;
      RECT  2.8 1.025 3.6 1.145 ;
      RECT  3.51 1.145 3.6 1.36 ;
      RECT  3.51 1.36 6.045 1.405 ;
      RECT  3.51 1.405 4.685 1.45 ;
      RECT  6.99 0.94 7.56 1.07 ;
      RECT  0.275 1.27 1.535 1.39 ;
      LAYER M2 ;
      RECT  4.31 0.95 7.2 1.05 ;
      LAYER V1 ;
      RECT  4.35 0.95 4.45 1.05 ;
      RECT  5.295 0.95 5.395 1.05 ;
      RECT  7.06 0.95 7.16 1.05 ;
  END
END SEN_FSDPQO_6
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPQO_8
#      Description : "D-Flip Flop w/scan, pos-edge triggered, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI)):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPQO_8
  CLASS CORE ;
  FOREIGN SEN_FSDPQO_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.095 0.75 8.275 0.93 ;
      RECT  8.095 0.93 8.185 1.225 ;
      RECT  8.095 1.225 8.285 1.345 ;
      RECT  7.555 0.675 7.8 0.775 ;
      RECT  7.555 0.775 7.665 0.97 ;
      RECT  5.385 0.75 5.78 0.92 ;
      LAYER M2 ;
      RECT  5.385 0.75 8.275 0.85 ;
      LAYER V1 ;
      RECT  8.135 0.75 8.235 0.85 ;
      RECT  7.555 0.75 7.655 0.85 ;
      RECT  5.425 0.75 5.525 0.85 ;
      RECT  5.625 0.75 5.725 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1611 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.75 1.45 0.855 ;
      RECT  0.945 0.855 1.45 0.945 ;
      LAYER M2 ;
      RECT  0.485 0.75 1.29 0.85 ;
      LAYER V1 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.75 0.51 11.45 0.69 ;
      RECT  11.08 0.69 11.25 1.11 ;
      RECT  9.75 1.11 11.45 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.4 0.51 2.515 0.905 ;
      RECT  0.485 0.55 0.69 0.65 ;
      RECT  0.485 0.65 0.605 0.965 ;
      LAYER M2 ;
      RECT  0.51 0.55 2.54 0.65 ;
      LAYER V1 ;
      RECT  2.4 0.55 2.5 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1188 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.055 ;
      RECT  0.15 1.055 2.13 1.145 ;
      RECT  2.04 0.935 2.13 1.055 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0474 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.94 0.51 9.06 1.34 ;
    END
    ANTENNADIFFAREA 0.142 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.235 0.185 1.75 ;
      RECT  0.0 1.75 11.8 1.85 ;
      RECT  0.56 1.485 0.73 1.75 ;
      RECT  2.1 1.435 2.22 1.75 ;
      RECT  2.6 1.435 2.72 1.75 ;
      RECT  3.13 1.435 3.245 1.75 ;
      RECT  4.73 1.51 4.85 1.75 ;
      RECT  5.265 1.495 5.385 1.75 ;
      RECT  5.795 1.495 5.965 1.75 ;
      RECT  6.34 1.44 6.46 1.75 ;
      RECT  6.86 1.44 6.98 1.75 ;
      RECT  8.63 1.615 8.8 1.75 ;
      RECT  9.495 1.435 9.615 1.75 ;
      RECT  10.0 1.39 10.145 1.75 ;
      RECT  10.52 1.39 10.665 1.75 ;
      RECT  11.04 1.39 11.185 1.75 ;
      RECT  11.59 1.21 11.71 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.8 0.05 ;
      RECT  2.46 0.05 2.63 0.175 ;
      RECT  3.03 0.05 3.2 0.175 ;
      RECT  4.69 0.05 4.86 0.175 ;
      RECT  1.625 0.05 1.795 0.19 ;
      RECT  8.63 0.05 8.8 0.22 ;
      RECT  6.835 0.05 7.005 0.32 ;
      RECT  0.09 0.05 0.23 0.39 ;
      RECT  10.015 0.05 10.135 0.395 ;
      RECT  10.535 0.05 10.655 0.395 ;
      RECT  11.055 0.05 11.175 0.395 ;
      RECT  5.29 0.05 5.43 0.41 ;
      RECT  9.495 0.05 9.61 0.425 ;
      RECT  6.34 0.05 6.46 0.43 ;
      RECT  11.59 0.05 11.71 0.59 ;
      RECT  5.82 0.05 5.94 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.395 0.14 3.98 0.23 ;
      RECT  3.395 0.23 3.5 0.28 ;
      RECT  3.86 0.23 3.98 0.33 ;
      RECT  0.545 0.28 3.5 0.37 ;
      RECT  0.545 0.37 2.695 0.4 ;
      RECT  2.605 0.4 2.695 1.255 ;
      RECT  1.63 1.255 3.425 1.345 ;
      RECT  1.63 1.345 1.75 1.48 ;
      RECT  3.335 1.345 3.425 1.54 ;
      RECT  1.055 1.48 1.75 1.6 ;
      RECT  3.335 1.54 4.12 1.66 ;
      RECT  8.37 0.14 8.54 0.31 ;
      RECT  8.37 0.31 9.345 0.4 ;
      RECT  9.225 0.205 9.345 0.31 ;
      RECT  9.225 0.4 9.345 1.165 ;
      RECT  4.325 0.265 5.17 0.355 ;
      RECT  4.76 0.355 5.17 0.385 ;
      RECT  4.325 0.355 4.415 0.63 ;
      RECT  4.76 0.385 4.85 1.05 ;
      RECT  4.26 0.63 4.415 0.805 ;
      RECT  4.76 1.05 5.105 1.22 ;
      RECT  7.12 0.26 7.24 0.41 ;
      RECT  7.03 0.41 7.785 0.505 ;
      RECT  7.615 0.38 7.785 0.41 ;
      RECT  7.03 0.505 7.13 0.545 ;
      RECT  6.03 0.545 7.13 0.665 ;
      RECT  7.04 0.665 7.13 1.23 ;
      RECT  6.05 1.23 7.825 1.35 ;
      RECT  4.13 0.29 4.235 0.42 ;
      RECT  3.59 0.42 4.235 0.51 ;
      RECT  3.59 0.51 3.705 0.735 ;
      RECT  3.59 0.735 3.785 0.79 ;
      RECT  3.0 0.79 3.785 0.895 ;
      RECT  3.695 0.895 3.785 1.18 ;
      RECT  3.695 1.18 4.39 1.27 ;
      RECT  0.795 0.51 2.105 0.615 ;
      RECT  5.205 0.54 5.73 0.66 ;
      RECT  5.205 0.66 5.295 0.77 ;
      RECT  4.94 0.77 5.295 0.88 ;
      RECT  5.195 0.88 5.295 1.08 ;
      RECT  5.195 1.08 5.68 1.19 ;
      RECT  8.36 0.49 8.505 0.66 ;
      RECT  8.415 0.66 8.505 1.0 ;
      RECT  8.335 1.0 8.505 1.06 ;
      RECT  8.335 1.06 8.81 1.15 ;
      RECT  8.72 0.735 8.81 1.06 ;
      RECT  2.2 0.5 2.31 0.735 ;
      RECT  1.72 0.735 2.31 0.825 ;
      RECT  1.72 0.825 1.81 0.955 ;
      RECT  2.22 0.825 2.31 0.995 ;
      RECT  2.22 0.995 2.435 1.165 ;
      RECT  3.91 0.72 4.08 0.81 ;
      RECT  3.99 0.81 4.08 0.99 ;
      RECT  3.99 0.99 4.49 1.09 ;
      RECT  4.31 0.95 4.49 0.99 ;
      RECT  5.87 0.78 6.72 0.895 ;
      RECT  5.87 0.895 5.96 1.315 ;
      RECT  4.58 0.59 4.67 1.315 ;
      RECT  4.58 1.315 5.96 1.36 ;
      RECT  2.785 0.51 3.5 0.625 ;
      RECT  2.785 0.625 2.89 1.025 ;
      RECT  2.785 1.025 3.605 1.13 ;
      RECT  3.515 1.13 3.605 1.36 ;
      RECT  3.515 1.36 5.96 1.405 ;
      RECT  3.515 1.405 4.66 1.45 ;
      RECT  9.52 0.785 10.97 0.895 ;
      RECT  9.52 0.895 9.61 1.255 ;
      RECT  9.225 1.255 9.61 1.345 ;
      RECT  9.225 1.345 9.315 1.435 ;
      RECT  7.355 0.175 8.005 0.265 ;
      RECT  7.355 0.265 7.525 0.305 ;
      RECT  7.915 0.265 8.005 1.435 ;
      RECT  7.915 1.435 9.315 1.465 ;
      RECT  7.37 1.465 9.315 1.525 ;
      RECT  7.37 1.525 8.135 1.58 ;
      RECT  7.22 0.835 7.45 1.13 ;
      RECT  0.275 1.26 1.54 1.38 ;
      LAYER M2 ;
      RECT  4.31 0.95 7.36 1.05 ;
      LAYER V1 ;
      RECT  4.35 0.95 4.45 1.05 ;
      RECT  5.195 0.95 5.295 1.05 ;
      RECT  7.22 0.95 7.32 1.05 ;
  END
END SEN_FSDPQO_8
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQ_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.5 6.05 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.43 0.29 5.53 0.89 ;
      RECT  3.385 0.24 3.685 0.49 ;
      LAYER M2 ;
      RECT  3.545 0.35 5.57 0.45 ;
      LAYER V1 ;
      RECT  5.43 0.35 5.53 0.45 ;
      RECT  3.585 0.35 3.685 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.042 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.485 ;
      RECT  0.365 0.485 0.65 0.585 ;
      RECT  0.55 0.585 0.65 1.08 ;
      RECT  0.55 1.08 1.445 1.17 ;
      RECT  1.355 1.0 1.445 1.08 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.39 1.44 0.52 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  1.43 1.615 1.6 1.75 ;
      RECT  1.94 1.615 2.11 1.75 ;
      RECT  3.58 1.495 3.71 1.75 ;
      RECT  3.845 1.5 4.015 1.75 ;
      RECT  4.965 1.22 5.085 1.75 ;
      RECT  5.595 1.44 5.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  2.085 0.05 2.255 0.18 ;
      RECT  1.365 0.05 1.495 0.36 ;
      RECT  4.855 0.05 4.975 0.39 ;
      RECT  0.31 0.05 0.44 0.395 ;
      RECT  3.8 0.05 3.92 0.56 ;
      RECT  5.68 0.05 5.8 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.34 0.215 4.745 0.305 ;
      RECT  4.655 0.305 4.745 0.65 ;
      RECT  4.655 0.65 5.16 0.675 ;
      RECT  4.63 0.675 5.16 0.74 ;
      RECT  5.055 0.74 5.16 0.82 ;
      RECT  4.63 0.74 4.72 1.495 ;
      RECT  4.39 1.495 4.72 1.585 ;
      RECT  1.615 0.28 2.805 0.4 ;
      RECT  1.615 0.4 1.705 0.45 ;
      RECT  0.785 0.18 0.905 0.45 ;
      RECT  0.785 0.45 1.705 0.54 ;
      RECT  4.07 0.3 4.19 0.43 ;
      RECT  4.07 0.43 4.285 0.52 ;
      RECT  4.195 0.52 4.285 1.13 ;
      RECT  3.325 0.865 3.84 0.965 ;
      RECT  3.75 0.965 3.84 1.13 ;
      RECT  3.75 1.13 4.285 1.225 ;
      RECT  4.375 0.43 4.565 0.6 ;
      RECT  4.375 0.6 4.465 1.315 ;
      RECT  3.38 1.315 4.465 1.405 ;
      RECT  3.38 1.405 3.47 1.57 ;
      RECT  2.695 0.66 2.785 1.57 ;
      RECT  2.695 1.57 3.47 1.66 ;
      RECT  1.8 0.49 2.13 0.61 ;
      RECT  2.04 0.61 2.13 0.775 ;
      RECT  2.04 0.775 2.37 0.885 ;
      RECT  2.04 0.885 2.13 1.225 ;
      RECT  1.64 1.225 2.13 1.345 ;
      RECT  2.34 0.51 2.59 0.63 ;
      RECT  2.5 0.63 2.59 1.09 ;
      RECT  2.235 1.09 2.59 1.19 ;
      RECT  2.92 0.41 3.04 0.65 ;
      RECT  2.92 0.65 4.06 0.655 ;
      RECT  2.885 0.655 4.06 0.74 ;
      RECT  3.97 0.74 4.06 1.04 ;
      RECT  2.885 0.74 3.005 1.475 ;
      RECT  5.62 0.785 5.86 0.895 ;
      RECT  5.62 0.895 5.71 1.205 ;
      RECT  5.065 0.3 5.34 0.42 ;
      RECT  5.25 0.42 5.34 0.91 ;
      RECT  4.81 0.83 4.905 0.91 ;
      RECT  4.81 0.91 5.34 1.0 ;
      RECT  5.25 1.0 5.34 1.205 ;
      RECT  5.25 1.205 5.71 1.31 ;
      RECT  5.25 1.31 5.375 1.59 ;
      RECT  3.145 1.115 3.66 1.225 ;
      RECT  3.145 1.225 3.265 1.48 ;
      RECT  0.055 0.17 0.175 1.26 ;
      RECT  0.055 1.26 0.82 1.35 ;
      RECT  0.73 1.35 0.82 1.57 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.73 1.57 1.28 1.66 ;
      RECT  0.92 1.295 1.46 1.415 ;
      RECT  1.37 1.415 1.46 1.435 ;
      RECT  1.37 1.435 2.605 1.525 ;
      RECT  2.485 1.29 2.605 1.435 ;
  END
END SEN_FSDPRBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQ_D_1P5
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQ_D_1P5
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQ_D_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.895 0.3 6.05 0.5 ;
      RECT  5.895 0.5 6.25 0.59 ;
      RECT  6.15 0.59 6.25 1.11 ;
      RECT  5.845 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.43 0.29 5.53 0.99 ;
      RECT  3.385 0.24 3.685 0.49 ;
      LAYER M2 ;
      RECT  3.545 0.35 5.57 0.45 ;
      LAYER V1 ;
      RECT  5.43 0.35 5.53 0.45 ;
      RECT  3.585 0.35 3.685 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.485 ;
      RECT  0.365 0.485 0.65 0.585 ;
      RECT  0.55 0.585 0.65 1.08 ;
      RECT  0.55 1.08 1.445 1.17 ;
      RECT  1.355 1.0 1.445 1.08 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.385 1.44 0.525 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  1.43 1.615 1.6 1.75 ;
      RECT  1.94 1.615 2.11 1.75 ;
      RECT  3.585 1.495 3.705 1.75 ;
      RECT  3.855 1.495 4.025 1.75 ;
      RECT  4.965 1.24 5.085 1.75 ;
      RECT  5.585 1.44 5.705 1.75 ;
      RECT  6.175 1.44 6.295 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  2.085 0.05 2.255 0.18 ;
      RECT  0.315 0.05 0.435 0.36 ;
      RECT  1.37 0.05 1.49 0.36 ;
      RECT  4.86 0.05 4.98 0.37 ;
      RECT  6.165 0.05 6.305 0.39 ;
      RECT  5.635 0.05 5.755 0.545 ;
      RECT  3.8 0.05 3.92 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.315 0.215 4.745 0.305 ;
      RECT  4.655 0.305 4.745 0.65 ;
      RECT  4.655 0.65 5.135 0.675 ;
      RECT  4.63 0.675 5.135 0.74 ;
      RECT  5.045 0.74 5.135 0.92 ;
      RECT  4.63 0.74 4.72 1.495 ;
      RECT  4.44 1.495 4.72 1.585 ;
      RECT  1.605 0.28 2.83 0.4 ;
      RECT  1.605 0.4 1.695 0.45 ;
      RECT  0.785 0.18 0.905 0.45 ;
      RECT  0.785 0.45 1.695 0.54 ;
      RECT  4.07 0.295 4.19 0.43 ;
      RECT  4.07 0.43 4.285 0.52 ;
      RECT  4.195 0.52 4.285 1.13 ;
      RECT  3.295 0.865 3.87 0.965 ;
      RECT  3.78 0.965 3.87 1.13 ;
      RECT  3.78 1.13 4.285 1.225 ;
      RECT  4.375 0.43 4.565 0.6 ;
      RECT  4.375 0.6 4.465 1.315 ;
      RECT  3.38 1.315 4.465 1.405 ;
      RECT  3.38 1.405 3.47 1.57 ;
      RECT  2.695 0.685 2.785 1.57 ;
      RECT  2.695 1.57 3.47 1.66 ;
      RECT  1.79 0.49 2.13 0.61 ;
      RECT  2.04 0.61 2.13 0.745 ;
      RECT  2.04 0.745 2.39 0.855 ;
      RECT  2.04 0.855 2.13 1.225 ;
      RECT  1.64 1.225 2.13 1.345 ;
      RECT  2.345 0.51 2.59 0.63 ;
      RECT  2.5 0.63 2.59 1.095 ;
      RECT  2.235 1.095 2.59 1.185 ;
      RECT  2.235 1.185 2.355 1.32 ;
      RECT  2.96 0.44 3.08 0.65 ;
      RECT  2.96 0.65 4.06 0.655 ;
      RECT  2.885 0.655 4.06 0.74 ;
      RECT  3.97 0.74 4.06 1.04 ;
      RECT  2.885 0.74 3.005 1.475 ;
      RECT  5.62 0.785 6.04 0.895 ;
      RECT  5.62 0.895 5.71 1.2 ;
      RECT  5.065 0.4 5.315 0.52 ;
      RECT  5.225 0.52 5.315 1.01 ;
      RECT  4.81 0.87 4.905 1.01 ;
      RECT  4.81 1.01 5.315 1.1 ;
      RECT  5.225 1.1 5.315 1.2 ;
      RECT  5.225 1.2 5.71 1.32 ;
      RECT  3.145 1.115 3.69 1.225 ;
      RECT  3.145 1.225 3.265 1.48 ;
      RECT  0.055 0.175 0.175 1.26 ;
      RECT  0.055 1.26 0.82 1.35 ;
      RECT  0.73 1.35 0.82 1.57 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.73 1.57 1.28 1.66 ;
      RECT  0.925 1.295 1.53 1.415 ;
      RECT  1.44 1.415 1.53 1.435 ;
      RECT  1.44 1.435 2.605 1.525 ;
      RECT  2.485 1.3 2.605 1.435 ;
  END
END SEN_FSDPRBQ_D_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.895 0.51 6.25 0.69 ;
      RECT  6.15 0.69 6.25 1.11 ;
      RECT  5.87 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.43 0.31 5.53 0.88 ;
      RECT  3.385 0.24 3.685 0.49 ;
      LAYER M2 ;
      RECT  3.545 0.35 5.57 0.45 ;
      LAYER V1 ;
      RECT  5.43 0.35 5.53 0.45 ;
      RECT  3.585 0.35 3.685 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.68 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.485 ;
      RECT  0.365 0.485 0.65 0.585 ;
      RECT  0.55 0.585 0.65 1.08 ;
      RECT  0.55 1.08 1.445 1.17 ;
      RECT  1.355 1.0 1.445 1.08 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.39 1.44 0.52 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  1.43 1.615 1.6 1.75 ;
      RECT  1.94 1.615 2.11 1.75 ;
      RECT  3.58 1.495 3.71 1.75 ;
      RECT  3.845 1.5 4.015 1.75 ;
      RECT  4.965 1.21 5.085 1.75 ;
      RECT  5.58 1.44 5.71 1.75 ;
      RECT  6.175 1.41 6.305 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  2.085 0.05 2.255 0.18 ;
      RECT  1.365 0.05 1.495 0.36 ;
      RECT  0.31 0.05 0.44 0.39 ;
      RECT  4.855 0.05 4.975 0.39 ;
      RECT  6.175 0.05 6.305 0.39 ;
      RECT  3.795 0.05 3.925 0.56 ;
      RECT  5.635 0.05 5.755 0.57 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.34 0.215 4.745 0.305 ;
      RECT  4.655 0.305 4.745 0.65 ;
      RECT  4.655 0.65 5.16 0.675 ;
      RECT  4.63 0.675 5.16 0.74 ;
      RECT  5.055 0.74 5.16 0.82 ;
      RECT  4.63 0.74 4.72 1.495 ;
      RECT  4.39 1.495 4.72 1.585 ;
      RECT  1.6 0.28 2.81 0.4 ;
      RECT  1.6 0.4 1.7 0.45 ;
      RECT  0.785 0.18 0.905 0.45 ;
      RECT  0.785 0.45 1.7 0.54 ;
      RECT  4.07 0.3 4.19 0.43 ;
      RECT  4.07 0.43 4.285 0.52 ;
      RECT  4.195 0.52 4.285 1.13 ;
      RECT  3.29 0.865 3.84 0.965 ;
      RECT  3.75 0.965 3.84 1.13 ;
      RECT  3.75 1.13 4.285 1.225 ;
      RECT  4.375 0.43 4.565 0.6 ;
      RECT  4.375 0.6 4.465 1.315 ;
      RECT  3.38 1.315 4.465 1.405 ;
      RECT  3.38 1.405 3.47 1.57 ;
      RECT  2.695 0.69 2.785 1.57 ;
      RECT  2.695 1.57 3.47 1.66 ;
      RECT  1.8 0.49 2.13 0.61 ;
      RECT  2.04 0.61 2.13 0.775 ;
      RECT  2.04 0.775 2.365 0.885 ;
      RECT  2.04 0.885 2.13 1.225 ;
      RECT  1.64 1.225 2.13 1.345 ;
      RECT  2.34 0.51 2.59 0.63 ;
      RECT  2.5 0.63 2.59 1.09 ;
      RECT  2.235 1.09 2.59 1.19 ;
      RECT  2.92 0.39 3.04 0.65 ;
      RECT  2.92 0.65 4.06 0.655 ;
      RECT  2.885 0.655 4.06 0.74 ;
      RECT  3.97 0.74 4.06 1.04 ;
      RECT  2.885 0.74 3.005 1.475 ;
      RECT  5.62 0.785 6.055 0.895 ;
      RECT  5.62 0.895 5.71 1.205 ;
      RECT  5.065 0.37 5.34 0.49 ;
      RECT  5.25 0.49 5.34 0.91 ;
      RECT  4.81 0.83 4.905 0.91 ;
      RECT  4.81 0.91 5.34 1.0 ;
      RECT  5.23 1.0 5.34 1.205 ;
      RECT  5.23 1.205 5.71 1.31 ;
      RECT  3.145 1.115 3.66 1.225 ;
      RECT  3.145 1.225 3.265 1.48 ;
      RECT  0.055 0.17 0.175 1.26 ;
      RECT  0.055 1.26 0.79 1.35 ;
      RECT  0.7 1.35 0.79 1.57 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.7 1.57 1.275 1.66 ;
      RECT  0.92 1.295 1.455 1.415 ;
      RECT  1.365 1.415 1.455 1.435 ;
      RECT  1.365 1.435 2.605 1.525 ;
      RECT  2.485 1.3 2.605 1.435 ;
  END
END SEN_FSDPRBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQ_D_3
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQ_D_3
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQ_D_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.895 0.51 6.535 0.69 ;
      RECT  6.35 0.69 6.45 1.11 ;
      RECT  5.87 1.11 6.535 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.43 0.29 5.53 0.91 ;
      RECT  3.385 0.24 3.685 0.49 ;
      LAYER M2 ;
      RECT  3.545 0.35 5.57 0.45 ;
      LAYER V1 ;
      RECT  5.43 0.35 5.53 0.45 ;
      RECT  3.585 0.35 3.685 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0663 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.485 ;
      RECT  0.36 0.485 0.65 0.585 ;
      RECT  0.55 0.585 0.65 1.08 ;
      RECT  0.55 1.08 1.445 1.17 ;
      RECT  1.355 1.0 1.445 1.08 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.385 1.44 0.525 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.43 1.615 1.6 1.75 ;
      RECT  1.94 1.615 2.11 1.75 ;
      RECT  3.585 1.495 3.705 1.75 ;
      RECT  3.855 1.495 4.025 1.75 ;
      RECT  4.965 1.24 5.085 1.75 ;
      RECT  5.585 1.385 5.705 1.75 ;
      RECT  6.155 1.44 6.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  2.085 0.05 2.255 0.18 ;
      RECT  0.315 0.05 0.435 0.36 ;
      RECT  1.37 0.05 1.49 0.36 ;
      RECT  4.86 0.05 4.98 0.36 ;
      RECT  6.155 0.05 6.275 0.37 ;
      RECT  3.8 0.05 3.92 0.56 ;
      RECT  5.635 0.05 5.755 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.34 0.22 4.745 0.34 ;
      RECT  4.655 0.34 4.745 0.65 ;
      RECT  4.655 0.65 5.135 0.675 ;
      RECT  4.63 0.675 5.135 0.74 ;
      RECT  5.045 0.74 5.135 0.85 ;
      RECT  4.63 0.74 4.72 1.495 ;
      RECT  4.415 1.495 4.72 1.6 ;
      RECT  1.605 0.28 2.83 0.4 ;
      RECT  1.605 0.4 1.695 0.45 ;
      RECT  0.785 0.19 0.905 0.45 ;
      RECT  0.785 0.45 1.695 0.54 ;
      RECT  4.07 0.295 4.19 0.43 ;
      RECT  4.07 0.43 4.285 0.52 ;
      RECT  4.195 0.52 4.285 1.13 ;
      RECT  3.295 0.865 3.865 0.965 ;
      RECT  3.775 0.965 3.865 1.13 ;
      RECT  3.775 1.13 4.285 1.225 ;
      RECT  4.375 0.43 4.565 0.6 ;
      RECT  4.375 0.6 4.465 1.315 ;
      RECT  3.38 1.315 4.465 1.405 ;
      RECT  3.38 1.405 3.47 1.57 ;
      RECT  2.695 0.685 2.785 1.57 ;
      RECT  2.695 1.57 3.47 1.66 ;
      RECT  1.79 0.49 2.13 0.61 ;
      RECT  2.04 0.61 2.13 0.745 ;
      RECT  2.04 0.745 2.38 0.855 ;
      RECT  2.04 0.855 2.13 1.225 ;
      RECT  1.645 1.225 2.13 1.345 ;
      RECT  2.34 0.51 2.59 0.63 ;
      RECT  2.5 0.63 2.59 1.095 ;
      RECT  2.235 1.095 2.59 1.185 ;
      RECT  2.235 1.185 2.355 1.31 ;
      RECT  2.92 0.41 3.04 0.65 ;
      RECT  2.92 0.65 4.06 0.655 ;
      RECT  2.885 0.655 4.06 0.74 ;
      RECT  3.97 0.74 4.06 1.04 ;
      RECT  2.885 0.74 3.005 1.475 ;
      RECT  5.62 0.795 6.24 0.905 ;
      RECT  5.62 0.905 5.71 1.16 ;
      RECT  5.045 0.44 5.315 0.56 ;
      RECT  5.225 0.56 5.315 0.94 ;
      RECT  4.81 0.83 4.905 0.94 ;
      RECT  4.81 0.94 5.315 1.03 ;
      RECT  5.225 1.03 5.315 1.16 ;
      RECT  5.225 1.16 5.71 1.28 ;
      RECT  3.145 1.115 3.685 1.225 ;
      RECT  3.145 1.225 3.265 1.48 ;
      RECT  0.055 0.18 0.175 1.26 ;
      RECT  0.055 1.26 0.82 1.35 ;
      RECT  0.73 1.35 0.82 1.57 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.73 1.57 1.28 1.66 ;
      RECT  0.925 1.295 1.46 1.415 ;
      RECT  1.37 1.415 1.46 1.435 ;
      RECT  1.37 1.435 2.605 1.525 ;
      RECT  2.485 1.305 2.605 1.435 ;
  END
END SEN_FSDPRBQ_D_3
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQ_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.845 0.51 6.485 0.69 ;
      RECT  6.35 0.69 6.45 1.11 ;
      RECT  5.82 1.11 6.485 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.4 0.3 5.5 0.745 ;
      RECT  5.4 0.745 5.53 0.915 ;
      RECT  3.385 0.24 3.685 0.49 ;
      LAYER M2 ;
      RECT  3.545 0.35 5.54 0.45 ;
      LAYER V1 ;
      RECT  5.4 0.35 5.5 0.45 ;
      RECT  3.585 0.35 3.685 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.485 ;
      RECT  0.36 0.485 0.65 0.585 ;
      RECT  0.55 0.585 0.65 1.08 ;
      RECT  0.55 1.08 1.445 1.17 ;
      RECT  1.355 1.0 1.445 1.08 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.39 1.44 0.52 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.43 1.615 1.6 1.75 ;
      RECT  1.94 1.615 2.11 1.75 ;
      RECT  3.58 1.495 3.71 1.75 ;
      RECT  3.845 1.5 4.015 1.75 ;
      RECT  4.965 1.21 5.085 1.75 ;
      RECT  5.58 1.41 5.71 1.75 ;
      RECT  6.1 1.41 6.23 1.75 ;
      RECT  6.62 1.41 6.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  2.085 0.05 2.255 0.18 ;
      RECT  1.365 0.05 1.495 0.36 ;
      RECT  4.855 0.05 4.985 0.375 ;
      RECT  0.31 0.05 0.44 0.39 ;
      RECT  6.1 0.05 6.23 0.39 ;
      RECT  6.62 0.05 6.74 0.39 ;
      RECT  3.795 0.05 3.925 0.56 ;
      RECT  5.59 0.05 5.705 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.34 0.215 4.745 0.305 ;
      RECT  4.655 0.305 4.745 0.65 ;
      RECT  4.655 0.65 5.13 0.675 ;
      RECT  4.63 0.675 5.13 0.74 ;
      RECT  5.025 0.74 5.13 0.82 ;
      RECT  4.63 0.74 4.72 1.495 ;
      RECT  4.39 1.495 4.72 1.585 ;
      RECT  1.595 0.28 2.83 0.4 ;
      RECT  1.595 0.4 1.695 0.45 ;
      RECT  0.785 0.18 0.905 0.45 ;
      RECT  0.785 0.45 1.695 0.54 ;
      RECT  4.07 0.29 4.19 0.43 ;
      RECT  4.07 0.43 4.285 0.52 ;
      RECT  4.195 0.52 4.285 1.13 ;
      RECT  3.285 0.865 3.84 0.965 ;
      RECT  3.75 0.965 3.84 1.13 ;
      RECT  3.75 1.13 4.285 1.225 ;
      RECT  4.375 0.43 4.565 0.6 ;
      RECT  4.375 0.6 4.465 1.315 ;
      RECT  3.38 1.315 4.465 1.405 ;
      RECT  3.38 1.405 3.47 1.57 ;
      RECT  2.695 0.66 2.785 1.57 ;
      RECT  2.695 1.57 3.47 1.66 ;
      RECT  1.79 0.49 2.13 0.61 ;
      RECT  2.04 0.61 2.13 0.775 ;
      RECT  2.04 0.775 2.365 0.885 ;
      RECT  2.04 0.885 2.13 1.225 ;
      RECT  1.65 1.225 2.13 1.345 ;
      RECT  2.34 0.51 2.59 0.63 ;
      RECT  2.5 0.63 2.59 1.09 ;
      RECT  2.22 1.09 2.59 1.19 ;
      RECT  2.92 0.41 3.04 0.65 ;
      RECT  2.92 0.65 4.06 0.655 ;
      RECT  2.885 0.655 4.06 0.74 ;
      RECT  3.97 0.74 4.06 1.04 ;
      RECT  2.885 0.74 3.005 1.475 ;
      RECT  5.62 0.785 6.25 0.895 ;
      RECT  5.62 0.895 5.71 1.14 ;
      RECT  5.05 0.44 5.31 0.56 ;
      RECT  5.22 0.56 5.31 0.91 ;
      RECT  4.81 0.875 4.905 0.91 ;
      RECT  4.81 0.91 5.31 1.045 ;
      RECT  5.2 1.045 5.31 1.14 ;
      RECT  5.2 1.14 5.71 1.26 ;
      RECT  3.145 1.115 3.66 1.225 ;
      RECT  3.145 1.225 3.265 1.48 ;
      RECT  0.055 0.17 0.175 1.26 ;
      RECT  0.055 1.26 0.8 1.35 ;
      RECT  0.71 1.35 0.8 1.57 ;
      RECT  0.055 1.35 0.175 1.63 ;
      RECT  0.71 1.57 1.275 1.66 ;
      RECT  0.93 1.295 1.465 1.415 ;
      RECT  1.365 1.415 1.465 1.435 ;
      RECT  1.365 1.435 2.605 1.525 ;
      RECT  2.485 1.3 2.605 1.435 ;
  END
END SEN_FSDPRBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.285 0.97 ;
      RECT  4.15 0.97 4.65 1.06 ;
      RECT  4.55 1.06 4.65 1.23 ;
      RECT  4.55 1.23 5.455 1.32 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0756 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.925 ;
      RECT  0.95 0.925 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0579 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.31 7.46 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.955 0.675 6.065 1.12 ;
      RECT  2.64 0.77 3.305 0.865 ;
      RECT  2.64 0.865 2.73 0.895 ;
      RECT  2.245 0.895 2.73 0.985 ;
      RECT  2.245 0.985 2.425 1.165 ;
      RECT  1.55 0.705 1.71 0.95 ;
      RECT  1.55 0.95 1.73 1.05 ;
      LAYER M2 ;
      RECT  1.55 0.95 6.095 1.05 ;
      LAYER V1 ;
      RECT  5.955 0.95 6.055 1.05 ;
      RECT  2.285 0.95 2.385 1.05 ;
      RECT  1.59 0.95 1.69 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.078 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0669 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.25 ;
      RECT  0.55 1.25 1.685 1.34 ;
      RECT  1.575 1.17 1.685 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.325 0.675 6.65 0.79 ;
      RECT  6.54 0.79 6.65 1.365 ;
      RECT  6.54 1.365 6.74 1.48 ;
    END
    ANTENNADIFFAREA 0.136 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.485 1.465 0.655 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  1.665 1.615 1.835 1.75 ;
      RECT  2.215 1.615 2.385 1.75 ;
      RECT  3.05 1.61 3.22 1.75 ;
      RECT  4.03 1.595 4.2 1.75 ;
      RECT  4.6 1.415 4.72 1.75 ;
      RECT  6.0 1.615 6.17 1.75 ;
      RECT  7.075 1.445 7.195 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  1.76 0.05 1.93 0.18 ;
      RECT  6.06 0.05 6.18 0.225 ;
      RECT  7.02 0.05 7.19 0.225 ;
      RECT  3.27 0.05 3.44 0.3 ;
      RECT  4.155 0.05 4.275 0.36 ;
      RECT  0.065 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.555 0.14 1.655 0.23 ;
      RECT  0.555 0.23 0.675 0.4 ;
      RECT  6.27 0.14 6.93 0.23 ;
      RECT  6.27 0.23 6.36 0.315 ;
      RECT  6.84 0.23 6.93 0.315 ;
      RECT  4.99 0.14 5.905 0.23 ;
      RECT  5.815 0.23 5.905 0.315 ;
      RECT  5.815 0.315 6.36 0.405 ;
      RECT  6.84 0.315 7.155 0.405 ;
      RECT  7.065 0.405 7.155 1.26 ;
      RECT  6.83 1.26 7.155 1.35 ;
      RECT  6.83 1.35 6.92 1.57 ;
      RECT  5.11 1.435 6.415 1.525 ;
      RECT  5.11 1.525 5.305 1.555 ;
      RECT  6.325 1.525 6.415 1.57 ;
      RECT  6.325 1.57 6.92 1.66 ;
      RECT  1.805 0.27 2.43 0.32 ;
      RECT  0.965 0.32 2.43 0.36 ;
      RECT  0.965 0.36 1.91 0.41 ;
      RECT  2.305 0.36 2.43 0.465 ;
      RECT  1.82 0.41 1.91 1.435 ;
      RECT  1.16 1.435 2.975 1.525 ;
      RECT  1.16 1.525 1.355 1.555 ;
      RECT  4.515 0.165 4.645 0.36 ;
      RECT  4.555 0.36 4.645 0.53 ;
      RECT  4.555 0.53 5.44 0.62 ;
      RECT  5.335 0.5 5.44 0.53 ;
      RECT  5.175 0.62 5.44 0.67 ;
      RECT  5.175 0.67 5.265 1.05 ;
      RECT  4.82 1.05 5.265 1.14 ;
      RECT  2.765 0.21 2.865 0.39 ;
      RECT  2.765 0.39 3.69 0.48 ;
      RECT  3.575 0.48 3.69 0.97 ;
      RECT  3.575 0.97 3.785 1.06 ;
      RECT  3.695 1.06 3.785 1.15 ;
      RECT  3.695 1.15 3.88 1.24 ;
      RECT  3.79 1.24 3.88 1.32 ;
      RECT  4.74 0.32 5.635 0.41 ;
      RECT  4.74 0.41 4.91 0.44 ;
      RECT  5.545 0.41 5.635 0.475 ;
      RECT  5.545 0.475 5.685 0.645 ;
      RECT  5.545 0.645 5.635 0.76 ;
      RECT  5.355 0.76 5.635 0.85 ;
      RECT  5.355 0.85 5.445 1.05 ;
      RECT  5.355 1.05 5.635 1.14 ;
      RECT  5.545 1.14 5.635 1.215 ;
      RECT  5.545 1.215 6.295 1.345 ;
      RECT  6.185 0.875 6.295 1.215 ;
      RECT  3.795 0.19 3.915 0.45 ;
      RECT  3.795 0.45 4.465 0.54 ;
      RECT  4.375 0.54 4.465 0.79 ;
      RECT  3.97 0.54 4.06 0.94 ;
      RECT  4.375 0.79 5.085 0.88 ;
      RECT  3.965 0.94 4.06 1.11 ;
      RECT  3.97 1.11 4.06 1.2 ;
      RECT  3.97 1.2 4.445 1.32 ;
      RECT  4.325 1.15 4.445 1.2 ;
      RECT  6.575 0.32 6.745 0.495 ;
      RECT  5.775 0.495 6.91 0.585 ;
      RECT  5.775 0.585 5.865 0.755 ;
      RECT  6.79 0.585 6.91 1.16 ;
      RECT  5.725 0.755 5.865 0.925 ;
      RECT  0.34 0.165 0.445 0.53 ;
      RECT  0.34 0.53 1.455 0.62 ;
      RECT  1.365 0.62 1.455 1.12 ;
      RECT  0.34 0.62 0.445 1.285 ;
      RECT  0.065 1.285 0.445 1.375 ;
      RECT  0.065 1.375 0.185 1.61 ;
      RECT  2.57 0.425 2.675 0.575 ;
      RECT  2.28 0.575 3.485 0.665 ;
      RECT  2.28 0.665 2.37 0.705 ;
      RECT  3.395 0.665 3.485 0.955 ;
      RECT  2.2 0.705 2.37 0.805 ;
      RECT  2.82 0.955 3.485 1.045 ;
      RECT  2.82 1.045 2.91 1.075 ;
      RECT  3.395 1.045 3.485 1.15 ;
      RECT  2.515 1.075 2.91 1.165 ;
      RECT  3.395 1.15 3.605 1.24 ;
      RECT  3.515 1.24 3.605 1.39 ;
      RECT  3.515 1.39 3.69 1.48 ;
      RECT  3.785 1.415 4.51 1.505 ;
      RECT  3.785 1.505 3.875 1.57 ;
      RECT  4.405 1.505 4.51 1.65 ;
      RECT  2.0 0.45 2.16 0.62 ;
      RECT  2.0 0.62 2.09 1.16 ;
      RECT  2.0 1.16 2.13 1.255 ;
      RECT  2.0 1.255 3.17 1.345 ;
      RECT  3.05 1.16 3.17 1.255 ;
      RECT  3.08 1.345 3.17 1.41 ;
      RECT  3.08 1.41 3.405 1.5 ;
      RECT  3.315 1.5 3.405 1.57 ;
      RECT  3.315 1.57 3.875 1.66 ;
  END
END SEN_FSDPRBQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.725 0.71 5.85 1.14 ;
      RECT  5.28 0.71 5.45 1.09 ;
      RECT  4.25 0.6 4.35 1.11 ;
      LAYER M2 ;
      RECT  4.21 0.95 5.865 1.05 ;
      LAYER V1 ;
      RECT  5.725 0.95 5.825 1.05 ;
      RECT  5.31 0.95 5.41 1.05 ;
      RECT  4.25 0.95 4.35 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.7 1.26 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.345 0.31 7.46 1.29 ;
    END
    ANTENNADIFFAREA 0.22 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.675 6.275 0.87 ;
      RECT  6.15 0.87 6.455 0.96 ;
      RECT  6.355 0.96 6.455 1.295 ;
      RECT  3.275 0.78 3.375 1.29 ;
      RECT  0.15 0.62 0.405 0.73 ;
      RECT  0.15 0.73 0.25 1.15 ;
      RECT  0.15 1.15 0.33 1.25 ;
      LAYER M2 ;
      RECT  0.15 1.15 6.495 1.25 ;
      LAYER V1 ;
      RECT  6.355 1.15 6.455 1.25 ;
      RECT  3.275 1.15 3.375 1.25 ;
      RECT  0.19 1.15 0.29 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.087 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.915 0.51 1.45 0.61 ;
      RECT  1.35 0.61 1.45 0.71 ;
      RECT  0.915 0.61 1.05 0.89 ;
      RECT  1.35 0.71 1.735 0.8 ;
      RECT  1.64 0.8 1.735 0.945 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0762 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.59 0.79 0.76 ;
      RECT  0.55 0.76 0.65 1.095 ;
      RECT  0.42 1.095 0.65 1.195 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.595 0.47 6.705 0.655 ;
      RECT  6.595 0.655 6.85 0.75 ;
      RECT  6.75 0.75 6.85 0.88 ;
      RECT  6.645 0.88 6.85 0.895 ;
      RECT  6.55 0.895 6.85 0.98 ;
      RECT  6.55 0.98 6.675 1.23 ;
      RECT  6.55 1.23 6.78 1.34 ;
    END
    ANTENNADIFFAREA 0.12 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.285 1.48 4.455 1.745 ;
      RECT  4.285 1.745 4.95 1.75 ;
      RECT  4.83 1.415 4.95 1.745 ;
      RECT  0.33 1.57 0.5 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  1.825 1.615 1.995 1.75 ;
      RECT  2.9 1.595 3.07 1.75 ;
      RECT  4.0 1.48 4.175 1.75 ;
      RECT  6.17 1.615 6.345 1.75 ;
      RECT  7.09 1.455 7.21 1.75 ;
      RECT  7.61 1.21 7.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  6.28 0.05 6.45 0.195 ;
      RECT  1.9 0.05 2.05 0.225 ;
      RECT  3.36 0.05 3.53 0.295 ;
      RECT  0.29 0.05 0.46 0.32 ;
      RECT  4.38 0.05 4.55 0.32 ;
      RECT  3.86 0.05 4.03 0.325 ;
      RECT  4.925 0.05 5.045 0.385 ;
      RECT  7.08 0.05 7.2 0.385 ;
      RECT  7.61 0.05 7.73 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  5.8 0.14 6.14 0.23 ;
      RECT  6.05 0.23 6.14 0.29 ;
      RECT  6.05 0.29 6.94 0.38 ;
      RECT  6.82 0.205 6.94 0.29 ;
      RECT  6.835 0.38 6.94 0.475 ;
      RECT  6.835 0.475 7.05 0.565 ;
      RECT  6.96 0.565 7.05 1.07 ;
      RECT  6.84 1.07 7.05 1.16 ;
      RECT  0.575 0.14 1.71 0.24 ;
      RECT  0.575 0.24 0.695 0.41 ;
      RECT  0.055 0.305 0.175 0.41 ;
      RECT  0.055 0.41 0.695 0.5 ;
      RECT  4.64 0.2 4.815 0.315 ;
      RECT  4.725 0.315 4.815 0.49 ;
      RECT  4.725 0.49 5.26 0.6 ;
      RECT  4.725 0.6 5.19 0.605 ;
      RECT  5.1 0.605 5.19 1.195 ;
      RECT  5.1 1.195 5.45 1.225 ;
      RECT  4.625 1.225 5.45 1.315 ;
      RECT  5.34 1.315 5.45 1.37 ;
      RECT  4.625 1.315 4.715 1.48 ;
      RECT  4.545 1.48 4.715 1.6 ;
      RECT  2.385 0.23 2.505 0.33 ;
      RECT  0.98 0.33 2.505 0.42 ;
      RECT  2.005 0.42 2.505 0.43 ;
      RECT  2.005 0.43 2.095 1.435 ;
      RECT  1.38 1.435 2.27 1.525 ;
      RECT  1.38 1.525 1.5 1.545 ;
      RECT  2.18 1.525 2.27 1.57 ;
      RECT  0.775 1.545 1.5 1.655 ;
      RECT  2.18 1.57 2.585 1.66 ;
      RECT  2.805 0.21 2.915 0.395 ;
      RECT  2.805 0.395 3.8 0.485 ;
      RECT  3.665 0.485 3.8 0.5 ;
      RECT  3.665 0.5 3.755 1.08 ;
      RECT  3.665 1.08 3.93 1.2 ;
      RECT  5.66 0.335 5.96 0.435 ;
      RECT  5.87 0.435 5.96 0.495 ;
      RECT  5.87 0.495 6.5 0.585 ;
      RECT  6.405 0.585 6.5 0.78 ;
      RECT  5.94 0.585 6.03 1.07 ;
      RECT  5.94 1.07 6.265 1.185 ;
      RECT  5.94 1.185 6.04 1.23 ;
      RECT  6.16 1.185 6.265 1.265 ;
      RECT  5.82 1.23 6.04 1.33 ;
      RECT  4.065 0.41 4.635 0.51 ;
      RECT  4.545 0.51 4.635 0.72 ;
      RECT  4.065 0.51 4.16 0.79 ;
      RECT  4.545 0.72 5.01 0.81 ;
      RECT  3.855 0.79 4.16 0.965 ;
      RECT  4.915 0.81 5.01 1.07 ;
      RECT  4.045 0.965 4.16 1.125 ;
      RECT  1.65 0.51 1.915 0.62 ;
      RECT  1.825 0.62 1.915 1.16 ;
      RECT  1.405 0.89 1.505 1.16 ;
      RECT  1.405 1.16 1.915 1.185 ;
      RECT  0.74 1.05 0.84 1.185 ;
      RECT  0.74 1.185 1.915 1.275 ;
      RECT  1.585 1.275 1.755 1.335 ;
      RECT  2.62 0.575 3.555 0.67 ;
      RECT  2.62 0.67 2.71 0.88 ;
      RECT  3.465 0.67 3.555 1.375 ;
      RECT  2.365 0.88 2.71 0.97 ;
      RECT  2.365 0.97 2.465 1.1 ;
      RECT  2.62 0.97 2.71 1.185 ;
      RECT  2.62 1.185 2.88 1.29 ;
      RECT  3.465 1.375 3.695 1.48 ;
      RECT  4.44 0.94 4.75 1.03 ;
      RECT  4.44 1.03 4.53 1.3 ;
      RECT  3.8 1.3 4.53 1.39 ;
      RECT  3.8 1.39 3.89 1.57 ;
      RECT  2.95 0.77 3.155 0.87 ;
      RECT  3.065 0.87 3.155 1.39 ;
      RECT  2.185 0.52 2.32 0.69 ;
      RECT  2.185 0.69 2.275 1.24 ;
      RECT  2.185 1.24 2.45 1.345 ;
      RECT  2.36 1.345 2.45 1.39 ;
      RECT  2.36 1.39 3.25 1.48 ;
      RECT  3.16 1.48 3.25 1.57 ;
      RECT  3.16 1.57 3.89 1.66 ;
      RECT  7.14 0.725 7.255 1.275 ;
      RECT  6.875 1.275 7.255 1.365 ;
      RECT  6.875 1.365 6.965 1.435 ;
      RECT  5.37 0.3 5.49 0.525 ;
      RECT  5.37 0.525 5.635 0.615 ;
      RECT  5.54 0.615 5.635 1.435 ;
      RECT  5.54 1.435 6.965 1.495 ;
      RECT  5.08 1.415 5.2 1.495 ;
      RECT  5.08 1.495 6.965 1.525 ;
      RECT  5.08 1.525 5.63 1.585 ;
      RECT  0.055 1.365 1.27 1.455 ;
      RECT  0.055 1.455 0.175 1.61 ;
  END
END SEN_FSDPRBQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.92 0.89 7.025 1.15 ;
      RECT  6.845 1.15 7.025 1.25 ;
      RECT  5.15 0.695 5.325 0.8 ;
      RECT  5.15 0.8 5.25 1.29 ;
      LAYER M2 ;
      RECT  5.11 1.15 7.05 1.25 ;
      LAYER V1 ;
      RECT  6.885 1.15 6.985 1.25 ;
      RECT  5.15 1.15 5.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1257 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.705 ;
      RECT  0.75 0.705 1.57 0.795 ;
      RECT  0.75 0.795 0.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0978 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.785 0.465 9.475 0.585 ;
      RECT  9.35 0.585 9.475 0.68 ;
      RECT  9.35 0.68 9.45 1.11 ;
      RECT  8.75 1.11 9.45 1.12 ;
      RECT  8.75 1.12 9.475 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.51 0.8 7.655 1.125 ;
      RECT  4.515 0.6 4.645 0.77 ;
      RECT  4.515 0.77 4.615 1.11 ;
      RECT  3.175 0.915 3.39 1.125 ;
      RECT  0.21 0.685 0.45 0.795 ;
      RECT  0.35 0.795 0.45 1.11 ;
      LAYER M2 ;
      RECT  0.31 0.95 7.655 1.05 ;
      LAYER V1 ;
      RECT  7.515 0.95 7.615 1.05 ;
      RECT  4.515 0.95 4.615 1.05 ;
      RECT  3.215 0.95 3.315 1.05 ;
      RECT  0.35 0.95 0.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0978 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.89 ;
      RECT  1.75 0.89 2.42 0.9 ;
      RECT  0.955 0.9 2.42 1.01 ;
      RECT  0.955 1.01 1.85 1.015 ;
      RECT  1.75 1.015 1.85 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0921 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 1.1 2.155 1.2 ;
      RECT  1.95 1.2 2.05 1.39 ;
      RECT  0.55 0.71 0.65 1.115 ;
      RECT  0.55 1.115 1.66 1.205 ;
      RECT  1.57 1.205 1.66 1.39 ;
      RECT  1.57 1.39 2.05 1.48 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.915 0.635 8.085 0.75 ;
      RECT  7.95 0.75 8.05 1.185 ;
      RECT  7.95 1.185 8.215 1.29 ;
    END
    ANTENNADIFFAREA 0.122 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  0.82 1.48 0.99 1.75 ;
      RECT  2.495 1.49 2.665 1.75 ;
      RECT  3.155 1.63 3.325 1.75 ;
      RECT  4.42 1.47 4.54 1.75 ;
      RECT  5.205 1.56 5.375 1.75 ;
      RECT  5.79 1.425 5.91 1.75 ;
      RECT  7.295 1.575 7.465 1.75 ;
      RECT  7.775 1.605 7.945 1.75 ;
      RECT  8.51 1.575 8.68 1.75 ;
      RECT  9.095 1.4 9.215 1.75 ;
      RECT  9.615 1.21 9.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  2.815 0.05 2.985 0.17 ;
      RECT  7.645 0.05 7.815 0.185 ;
      RECT  8.51 0.05 8.68 0.185 ;
      RECT  4.65 0.05 4.82 0.2 ;
      RECT  5.69 0.05 5.86 0.235 ;
      RECT  6.24 0.05 6.41 0.235 ;
      RECT  5.155 0.05 5.325 0.36 ;
      RECT  0.325 0.05 0.465 0.365 ;
      RECT  9.095 0.05 9.215 0.375 ;
      RECT  9.615 0.05 9.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.57 0.14 2.255 0.23 ;
      RECT  0.57 0.23 0.725 0.39 ;
      RECT  0.57 0.39 0.66 0.455 ;
      RECT  0.065 0.32 0.185 0.455 ;
      RECT  0.065 0.455 0.66 0.545 ;
      RECT  6.605 0.155 7.1 0.245 ;
      RECT  6.605 0.245 6.695 0.34 ;
      RECT  5.53 0.34 6.695 0.43 ;
      RECT  5.53 0.43 5.625 0.47 ;
      RECT  4.915 0.47 5.625 0.58 ;
      RECT  5.53 0.58 5.625 0.775 ;
      RECT  4.915 0.58 5.005 1.07 ;
      RECT  5.53 0.775 6.27 0.865 ;
      RECT  6.18 0.865 6.27 0.945 ;
      RECT  6.18 0.945 6.44 1.065 ;
      RECT  4.915 1.07 5.045 1.275 ;
      RECT  3.115 0.21 3.825 0.26 ;
      RECT  2.775 0.26 3.825 0.32 ;
      RECT  1.015 0.32 3.825 0.33 ;
      RECT  1.015 0.33 3.205 0.35 ;
      RECT  1.015 0.35 2.88 0.41 ;
      RECT  2.79 0.41 2.88 0.875 ;
      RECT  2.69 0.875 2.88 0.965 ;
      RECT  2.69 0.965 2.78 1.31 ;
      RECT  2.315 1.31 2.85 1.4 ;
      RECT  2.76 1.4 2.85 1.45 ;
      RECT  2.315 1.4 2.405 1.57 ;
      RECT  2.76 1.45 3.945 1.54 ;
      RECT  1.08 1.48 1.25 1.57 ;
      RECT  1.08 1.57 2.405 1.66 ;
      RECT  4.945 0.18 5.05 0.29 ;
      RECT  4.115 0.29 5.05 0.38 ;
      RECT  4.115 0.38 4.22 0.655 ;
      RECT  4.735 0.38 4.825 1.025 ;
      RECT  3.675 0.655 4.22 0.745 ;
      RECT  3.675 0.745 3.775 0.985 ;
      RECT  4.705 1.025 4.825 1.195 ;
      RECT  7.2 0.275 8.61 0.34 ;
      RECT  6.79 0.34 8.61 0.365 ;
      RECT  6.79 0.365 7.29 0.43 ;
      RECT  8.52 0.365 8.61 0.78 ;
      RECT  6.79 0.43 6.915 0.67 ;
      RECT  8.52 0.78 9.24 0.9 ;
      RECT  8.52 0.9 8.61 1.395 ;
      RECT  6.92 1.395 8.61 1.46 ;
      RECT  6.26 1.46 8.61 1.485 ;
      RECT  6.26 1.485 7.01 1.55 ;
      RECT  3.915 0.32 4.025 0.425 ;
      RECT  3.37 0.425 4.025 0.515 ;
      RECT  3.37 0.515 3.46 0.735 ;
      RECT  3.195 0.735 3.57 0.825 ;
      RECT  3.48 0.825 3.57 1.075 ;
      RECT  3.48 1.075 4.12 1.165 ;
      RECT  7.415 0.455 8.405 0.545 ;
      RECT  7.415 0.545 7.505 0.57 ;
      RECT  8.315 0.545 8.405 1.255 ;
      RECT  7.3 0.57 7.505 0.66 ;
      RECT  7.3 0.66 7.39 0.77 ;
      RECT  1.245 0.5 2.505 0.605 ;
      RECT  5.96 0.52 6.68 0.62 ;
      RECT  6.53 0.62 6.62 1.235 ;
      RECT  5.545 1.235 6.62 1.28 ;
      RECT  5.545 1.28 6.715 1.335 ;
      RECT  6.545 1.335 6.715 1.37 ;
      RECT  5.545 1.335 5.65 1.46 ;
      RECT  7.03 0.52 7.21 0.635 ;
      RECT  7.115 0.635 7.21 1.215 ;
      RECT  7.115 1.215 7.85 1.305 ;
      RECT  7.745 0.87 7.85 1.215 ;
      RECT  2.595 0.5 2.7 0.695 ;
      RECT  1.96 0.695 2.7 0.785 ;
      RECT  1.96 0.785 2.6 0.8 ;
      RECT  2.51 0.8 2.6 1.105 ;
      RECT  2.32 1.105 2.6 1.195 ;
      RECT  5.58 0.955 6.04 1.035 ;
      RECT  5.365 1.035 6.04 1.055 ;
      RECT  5.365 1.055 5.71 1.125 ;
      RECT  5.365 1.125 5.455 1.38 ;
      RECT  2.995 0.44 3.27 0.61 ;
      RECT  2.995 0.61 3.085 1.05 ;
      RECT  2.91 1.05 3.085 1.22 ;
      RECT  2.995 1.22 3.085 1.26 ;
      RECT  2.995 1.26 4.425 1.285 ;
      RECT  4.32 0.805 4.425 1.26 ;
      RECT  2.995 1.285 4.755 1.35 ;
      RECT  4.335 1.35 4.755 1.375 ;
      RECT  4.665 1.375 4.755 1.38 ;
      RECT  4.665 1.38 5.455 1.47 ;
      RECT  0.065 1.3 1.48 1.39 ;
      RECT  0.56 1.39 0.73 1.45 ;
      RECT  1.36 1.39 1.48 1.48 ;
      RECT  0.065 1.39 0.185 1.56 ;
  END
END SEN_FSDPRBQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQO_6
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQO_6
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQO_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.125 0.685 7.295 0.775 ;
      RECT  7.125 0.775 7.25 1.135 ;
      RECT  7.125 1.135 7.72 1.225 ;
      RECT  7.54 1.225 7.72 1.305 ;
      RECT  2.52 0.77 2.7 1.25 ;
      LAYER M2 ;
      RECT  2.52 1.15 7.72 1.25 ;
      LAYER V1 ;
      RECT  7.58 1.15 7.68 1.25 ;
      RECT  2.56 1.15 2.66 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1476 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1146 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.11 0.31 9.25 0.51 ;
      RECT  9.11 0.51 10.25 0.69 ;
      RECT  10.12 0.69 10.25 1.11 ;
      RECT  8.95 1.11 10.25 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.805 0.195 8.085 0.285 ;
      RECT  7.805 0.285 7.99 0.45 ;
      RECT  4.455 0.14 4.675 0.45 ;
      LAYER M2 ;
      RECT  4.485 0.35 7.99 0.45 ;
      LAYER V1 ;
      RECT  7.85 0.35 7.95 0.45 ;
      RECT  4.525 0.35 4.625 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1062 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.625 1.56 0.735 ;
      RECT  0.75 0.735 0.85 0.95 ;
      RECT  0.75 0.95 0.99 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.825 ;
      RECT  1.11 0.825 1.85 0.93 ;
      RECT  1.75 0.93 1.85 1.09 ;
      RECT  1.11 0.93 1.21 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.425 0.47 8.535 0.68 ;
      RECT  8.425 0.68 8.65 0.77 ;
      RECT  8.55 0.77 8.65 1.045 ;
      RECT  8.37 1.045 8.65 1.165 ;
    END
    ANTENNADIFFAREA 0.109 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.405 0.48 1.75 ;
      RECT  0.0 1.75 10.6 1.85 ;
      RECT  0.945 1.58 1.115 1.75 ;
      RECT  2.555 1.54 2.675 1.75 ;
      RECT  4.235 1.495 4.405 1.75 ;
      RECT  4.815 1.54 4.935 1.75 ;
      RECT  5.38 1.39 5.5 1.75 ;
      RECT  5.9 1.39 6.02 1.75 ;
      RECT  6.425 1.405 6.53 1.75 ;
      RECT  8.065 1.48 8.185 1.75 ;
      RECT  8.81 1.475 8.99 1.75 ;
      RECT  9.365 1.39 9.485 1.75 ;
      RECT  9.885 1.39 10.005 1.75 ;
      RECT  10.405 1.21 10.525 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.6 0.05 ;
      RECT  2.28 0.05 2.405 0.225 ;
      RECT  2.875 0.05 2.995 0.225 ;
      RECT  4.765 0.05 4.89 0.39 ;
      RECT  8.845 0.05 8.965 0.395 ;
      RECT  8.175 0.05 8.265 0.405 ;
      RECT  9.36 0.05 9.49 0.41 ;
      RECT  9.885 0.05 10.005 0.41 ;
      RECT  6.335 0.05 6.44 0.43 ;
      RECT  5.81 0.05 5.93 0.445 ;
      RECT  5.28 0.05 5.4 0.59 ;
      RECT  10.405 0.05 10.525 0.59 ;
      RECT  0.065 0.05 0.185 0.68 ;
      RECT  8.095 0.405 8.265 0.495 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  8.495 0.14 8.755 0.23 ;
      RECT  8.665 0.23 8.755 0.485 ;
      RECT  8.665 0.485 8.83 0.575 ;
      RECT  8.74 0.575 8.83 1.295 ;
      RECT  7.76 0.775 8.155 0.865 ;
      RECT  8.065 0.865 8.155 1.295 ;
      RECT  8.065 1.295 8.83 1.385 ;
      RECT  8.065 1.385 8.68 1.39 ;
      RECT  8.59 1.39 8.68 1.635 ;
      RECT  1.44 0.19 2.18 0.315 ;
      RECT  1.44 0.315 3.865 0.32 ;
      RECT  3.17 0.24 3.865 0.315 ;
      RECT  1.97 0.32 3.865 0.36 ;
      RECT  1.97 0.36 3.265 0.42 ;
      RECT  1.97 0.42 2.06 1.27 ;
      RECT  1.97 1.27 2.155 1.285 ;
      RECT  1.48 1.285 2.155 1.36 ;
      RECT  1.48 1.36 3.76 1.395 ;
      RECT  3.64 1.28 3.76 1.36 ;
      RECT  2.035 1.395 3.76 1.45 ;
      RECT  0.525 0.205 1.215 0.32 ;
      RECT  0.525 0.32 0.625 0.49 ;
      RECT  6.53 0.215 7.315 0.335 ;
      RECT  6.53 0.335 6.62 0.635 ;
      RECT  6.02 0.635 6.62 0.755 ;
      RECT  6.53 0.755 6.62 1.115 ;
      RECT  6.53 1.115 6.725 1.135 ;
      RECT  5.615 1.135 6.725 1.26 ;
      RECT  6.62 1.26 6.725 1.495 ;
      RECT  6.62 1.495 7.27 1.595 ;
      RECT  6.9 0.445 7.005 0.475 ;
      RECT  6.9 0.475 7.49 0.595 ;
      RECT  7.39 0.595 7.49 0.71 ;
      RECT  6.9 0.595 7.01 1.285 ;
      RECT  6.84 1.285 7.01 1.315 ;
      RECT  6.84 1.315 7.45 1.405 ;
      RECT  7.36 1.405 7.45 1.465 ;
      RECT  7.36 1.465 7.555 1.555 ;
      RECT  0.735 0.41 1.88 0.515 ;
      RECT  1.775 0.515 1.88 0.605 ;
      RECT  4.19 0.29 4.29 0.545 ;
      RECT  4.19 0.545 5.165 0.665 ;
      RECT  3.38 0.45 4.1 0.56 ;
      RECT  3.97 0.56 4.1 0.76 ;
      RECT  3.97 0.76 5.06 0.86 ;
      RECT  3.97 0.86 4.06 1.035 ;
      RECT  4.89 0.86 5.06 1.055 ;
      RECT  3.37 1.035 4.06 1.14 ;
      RECT  3.37 1.14 3.51 1.21 ;
      RECT  3.97 1.14 4.06 1.255 ;
      RECT  3.97 1.255 4.35 1.315 ;
      RECT  3.97 1.315 4.585 1.345 ;
      RECT  4.265 1.345 4.585 1.405 ;
      RECT  4.495 1.405 4.585 1.57 ;
      RECT  4.495 1.57 4.705 1.66 ;
      RECT  7.58 0.39 7.71 0.595 ;
      RECT  7.58 0.595 8.335 0.685 ;
      RECT  8.245 0.685 8.335 0.945 ;
      RECT  7.58 0.685 7.67 0.955 ;
      RECT  7.58 0.955 7.975 1.045 ;
      RECT  7.885 1.045 7.975 1.45 ;
      RECT  7.645 1.45 7.975 1.57 ;
      RECT  2.34 0.51 3.04 0.63 ;
      RECT  2.94 0.63 3.04 0.975 ;
      RECT  2.34 0.63 2.43 1.18 ;
      RECT  2.815 0.975 3.04 1.08 ;
      RECT  2.255 1.18 2.43 1.27 ;
      RECT  8.92 0.51 9.02 0.79 ;
      RECT  8.92 0.79 10.01 0.895 ;
      RECT  3.16 0.525 3.28 0.845 ;
      RECT  3.16 0.845 3.865 0.945 ;
      RECT  3.16 0.945 3.28 1.17 ;
      RECT  2.8 1.17 3.28 1.27 ;
      RECT  5.55 0.245 5.67 0.93 ;
      RECT  5.55 0.93 6.315 0.95 ;
      RECT  5.405 0.95 6.315 1.04 ;
      RECT  5.405 1.04 5.525 1.145 ;
      RECT  4.18 1.045 4.745 1.145 ;
      RECT  4.18 1.145 5.525 1.15 ;
      RECT  4.65 1.15 5.525 1.25 ;
      RECT  6.71 0.49 6.81 1.025 ;
      RECT  1.3 1.055 1.56 1.165 ;
      RECT  1.3 1.165 1.39 1.21 ;
      RECT  0.325 0.535 0.445 0.735 ;
      RECT  0.325 0.735 0.65 0.845 ;
      RECT  0.56 0.845 0.65 1.21 ;
      RECT  0.065 1.21 1.39 1.3 ;
      RECT  0.065 1.3 0.185 1.61 ;
      RECT  0.61 1.39 1.39 1.485 ;
      RECT  0.61 1.485 1.945 1.49 ;
      RECT  1.29 1.49 1.945 1.6 ;
      RECT  4.0 1.455 4.12 1.555 ;
      RECT  3.045 1.555 4.12 1.66 ;
      LAYER M2 ;
      RECT  0.485 0.35 4.33 0.45 ;
      RECT  2.895 0.55 6.85 0.65 ;
      RECT  7.35 0.55 9.065 0.65 ;
      LAYER V1 ;
      RECT  0.525 0.35 0.625 0.45 ;
      RECT  4.19 0.35 4.29 0.45 ;
      RECT  2.94 0.55 3.04 0.65 ;
      RECT  6.71 0.55 6.81 0.65 ;
      RECT  7.39 0.55 7.49 0.65 ;
      RECT  8.92 0.55 9.02 0.65 ;
  END
END SEN_FSDPRBQO_6
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBQO_8
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBQO_8
  CLASS CORE ;
  FOREIGN SEN_FSDPRBQO_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.6 8.05 1.16 ;
      RECT  7.95 1.16 8.21 1.33 ;
      RECT  5.825 0.575 5.93 0.985 ;
      LAYER M2 ;
      RECT  5.785 0.75 8.09 0.85 ;
      LAYER V1 ;
      RECT  7.95 0.75 8.05 0.85 ;
      RECT  5.825 0.75 5.925 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1581 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.62 ;
      RECT  0.75 0.62 0.95 0.71 ;
      RECT  0.85 0.71 0.95 0.955 ;
      RECT  0.85 0.955 2.05 1.045 ;
      RECT  1.95 1.045 2.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.715 0.51 11.445 0.69 ;
      RECT  10.91 0.69 11.09 1.095 ;
      RECT  10.91 1.095 11.4 1.11 ;
      RECT  9.715 1.11 11.4 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 0.945 8.84 1.115 ;
      RECT  4.83 0.67 4.94 1.16 ;
      RECT  3.5 0.72 3.61 1.125 ;
      RECT  0.35 0.71 0.495 0.95 ;
      RECT  0.35 0.95 0.54 1.05 ;
      LAYER M2 ;
      RECT  0.36 0.95 8.785 1.05 ;
      LAYER V1 ;
      RECT  8.645 0.95 8.745 1.05 ;
      RECT  4.84 0.95 4.94 1.05 ;
      RECT  3.51 0.95 3.61 1.05 ;
      RECT  0.4 0.95 0.5 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END RD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.69 0.71 2.79 1.195 ;
      RECT  1.805 0.75 1.985 0.775 ;
      RECT  1.06 0.775 1.985 0.865 ;
      LAYER M2 ;
      RECT  1.805 0.75 2.83 0.85 ;
      LAYER V1 ;
      RECT  2.69 0.75 2.79 0.85 ;
      RECT  1.845 0.75 1.945 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1104 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 1.015 2.375 1.115 ;
      RECT  2.15 1.115 2.25 1.39 ;
      RECT  0.665 0.8 0.76 1.135 ;
      RECT  0.665 1.135 1.85 1.2 ;
      RECT  0.15 0.71 0.25 1.2 ;
      RECT  0.15 1.2 1.85 1.225 ;
      RECT  0.15 1.225 0.76 1.29 ;
      RECT  1.75 1.225 1.85 1.39 ;
      RECT  1.75 1.39 2.25 1.48 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0474 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.075 0.51 9.25 0.68 ;
      RECT  9.13 0.68 9.25 1.165 ;
      RECT  9.13 1.165 9.265 1.335 ;
    END
    ANTENNADIFFAREA 0.106 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.405 0.195 1.75 ;
      RECT  0.0 1.75 12.0 1.85 ;
      RECT  0.615 1.605 0.785 1.75 ;
      RECT  2.65 1.61 2.82 1.75 ;
      RECT  3.375 1.615 3.545 1.75 ;
      RECT  4.895 1.45 5.015 1.75 ;
      RECT  5.365 1.45 5.485 1.75 ;
      RECT  5.92 1.45 6.04 1.75 ;
      RECT  6.485 1.37 6.605 1.75 ;
      RECT  7.005 1.405 7.125 1.75 ;
      RECT  8.58 1.61 8.755 1.75 ;
      RECT  9.39 1.605 9.56 1.75 ;
      RECT  9.96 1.39 10.105 1.75 ;
      RECT  10.48 1.39 10.625 1.75 ;
      RECT  11.0 1.39 11.145 1.75 ;
      RECT  11.535 1.205 11.655 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.0 0.05 ;
      RECT  2.79 0.05 2.96 0.185 ;
      RECT  3.355 0.05 3.475 0.24 ;
      RECT  8.815 0.05 8.935 0.24 ;
      RECT  9.345 0.05 9.515 0.24 ;
      RECT  5.94 0.05 6.11 0.305 ;
      RECT  6.46 0.05 6.63 0.315 ;
      RECT  6.98 0.05 7.15 0.315 ;
      RECT  0.315 0.05 0.435 0.36 ;
      RECT  5.445 0.05 5.56 0.365 ;
      RECT  5.0 0.05 5.12 0.38 ;
      RECT  9.96 0.05 10.11 0.41 ;
      RECT  10.48 0.05 10.63 0.41 ;
      RECT  11.0 0.05 11.15 0.41 ;
      RECT  11.535 0.05 11.655 0.63 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  7.5 0.14 8.59 0.23 ;
      RECT  8.5 0.23 8.59 0.33 ;
      RECT  7.5 0.23 7.67 0.355 ;
      RECT  8.02 0.23 8.19 0.39 ;
      RECT  8.5 0.33 9.595 0.42 ;
      RECT  9.49 0.42 9.595 0.805 ;
      RECT  9.49 0.805 10.82 0.92 ;
      RECT  9.49 0.92 9.58 1.425 ;
      RECT  7.4 1.425 9.58 1.515 ;
      RECT  7.4 1.515 8.115 1.55 ;
      RECT  1.17 0.14 2.545 0.24 ;
      RECT  0.55 0.33 2.22 0.42 ;
      RECT  0.55 0.42 0.64 0.45 ;
      RECT  0.055 0.175 0.175 0.45 ;
      RECT  0.055 0.45 0.64 0.54 ;
      RECT  7.76 0.33 7.93 0.42 ;
      RECT  7.76 0.42 7.915 0.445 ;
      RECT  6.24 0.27 6.345 0.405 ;
      RECT  6.24 0.405 7.37 0.445 ;
      RECT  7.28 0.25 7.37 0.405 ;
      RECT  6.24 0.445 7.915 0.495 ;
      RECT  7.28 0.495 7.915 0.51 ;
      RECT  7.28 0.51 7.855 0.535 ;
      RECT  7.685 0.535 7.855 1.095 ;
      RECT  6.2 1.095 7.855 1.22 ;
      RECT  2.31 0.335 4.03 0.425 ;
      RECT  2.88 0.425 4.03 0.445 ;
      RECT  2.31 0.425 2.4 0.515 ;
      RECT  2.88 0.445 2.97 1.41 ;
      RECT  1.05 0.51 1.14 0.515 ;
      RECT  1.05 0.515 2.4 0.605 ;
      RECT  1.05 0.605 1.14 0.68 ;
      RECT  2.88 1.41 3.745 1.43 ;
      RECT  2.435 1.43 3.745 1.48 ;
      RECT  2.435 1.48 4.105 1.5 ;
      RECT  2.435 1.5 2.995 1.52 ;
      RECT  3.645 1.5 4.105 1.59 ;
      RECT  2.435 1.52 2.525 1.57 ;
      RECT  1.2 1.495 1.37 1.57 ;
      RECT  1.2 1.57 2.525 1.66 ;
      RECT  3.985 1.59 4.105 1.66 ;
      RECT  5.645 0.395 6.145 0.485 ;
      RECT  6.055 0.485 6.145 0.585 ;
      RECT  5.645 0.485 5.735 0.815 ;
      RECT  6.055 0.585 7.1 0.675 ;
      RECT  7.01 0.675 7.1 0.78 ;
      RECT  7.01 0.78 7.45 0.95 ;
      RECT  5.21 0.815 5.735 0.905 ;
      RECT  5.61 0.905 5.735 1.075 ;
      RECT  5.61 1.075 5.805 1.18 ;
      RECT  8.28 0.32 8.41 0.49 ;
      RECT  8.28 0.49 8.37 0.93 ;
      RECT  8.28 0.93 8.405 1.02 ;
      RECT  8.31 1.02 8.405 1.245 ;
      RECT  8.31 1.245 9.04 1.335 ;
      RECT  8.93 0.84 9.04 1.245 ;
      RECT  4.095 0.525 4.265 0.535 ;
      RECT  3.32 0.535 4.265 0.63 ;
      RECT  4.095 0.63 4.265 0.645 ;
      RECT  3.32 0.63 3.41 0.9 ;
      RECT  3.73 0.63 3.825 0.965 ;
      RECT  3.71 0.965 3.825 1.01 ;
      RECT  3.71 1.01 4.4 1.11 ;
      RECT  3.71 1.11 3.815 1.135 ;
      RECT  4.23 1.11 4.4 1.21 ;
      RECT  4.355 0.47 5.38 0.56 ;
      RECT  5.26 0.56 5.38 0.7 ;
      RECT  4.355 0.56 4.445 0.75 ;
      RECT  5.03 0.56 5.12 1.035 ;
      RECT  4.29 0.75 4.445 0.92 ;
      RECT  5.03 1.035 5.35 1.155 ;
      RECT  2.51 0.515 2.715 0.615 ;
      RECT  2.51 0.615 2.6 0.775 ;
      RECT  2.12 0.775 2.6 0.895 ;
      RECT  2.48 0.895 2.6 1.225 ;
      RECT  11.805 0.215 11.925 0.745 ;
      RECT  11.555 0.745 11.925 0.85 ;
      RECT  11.805 0.85 11.925 1.615 ;
      RECT  8.46 0.65 8.75 0.85 ;
      RECT  6.02 0.765 6.89 0.87 ;
      RECT  6.02 0.87 6.11 1.27 ;
      RECT  4.72 1.27 6.11 1.3 ;
      RECT  3.06 0.535 3.23 1.0 ;
      RECT  3.06 1.0 3.265 1.17 ;
      RECT  3.175 1.17 3.265 1.23 ;
      RECT  3.175 1.23 4.085 1.3 ;
      RECT  3.175 1.3 6.11 1.32 ;
      RECT  3.935 1.32 6.11 1.36 ;
      RECT  3.935 1.36 4.805 1.39 ;
      RECT  4.685 1.39 4.805 1.62 ;
      RECT  0.91 1.315 1.66 1.405 ;
      RECT  0.91 1.405 1.01 1.425 ;
      RECT  0.29 1.425 1.01 1.515 ;
      LAYER M2 ;
      RECT  8.46 0.75 11.755 0.85 ;
      LAYER V1 ;
      RECT  8.51 0.75 8.61 0.85 ;
      RECT  11.595 0.75 11.695 0.85 ;
  END
END SEN_FSDPRBQO_8
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBSBQ_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBSBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDPRBSBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.775 0.555 3.875 1.125 ;
      RECT  3.775 1.125 4.105 1.22 ;
      RECT  1.58 0.865 1.885 0.97 ;
      RECT  1.785 0.97 1.885 1.09 ;
      LAYER M2 ;
      RECT  1.745 0.95 3.915 1.05 ;
      LAYER V1 ;
      RECT  3.775 0.95 3.875 1.05 ;
      RECT  1.785 0.95 1.885 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.115 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.31 5.9 0.505 ;
      RECT  5.75 0.505 5.85 1.11 ;
      RECT  5.55 1.11 5.85 1.3 ;
      RECT  5.55 1.3 5.65 1.43 ;
      RECT  5.52 1.43 5.65 1.6 ;
    END
    ANTENNADIFFAREA 0.137 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.94 0.48 5.05 0.91 ;
      RECT  2.605 0.55 3.075 0.65 ;
      LAYER M2 ;
      RECT  2.895 0.55 4.305 0.65 ;
      RECT  4.205 0.65 4.305 0.75 ;
      RECT  4.205 0.75 5.08 0.85 ;
      LAYER V1 ;
      RECT  4.94 0.75 5.04 0.85 ;
      RECT  2.935 0.55 3.035 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.14 4.45 0.23 ;
      RECT  4.35 0.23 4.45 0.31 ;
      RECT  3.35 0.23 3.45 0.535 ;
      RECT  4.35 0.31 4.65 0.49 ;
      RECT  4.55 0.49 4.65 0.51 ;
      RECT  4.55 0.51 4.67 0.69 ;
      RECT  3.2 0.535 3.45 0.625 ;
      RECT  3.2 0.625 3.29 0.77 ;
      RECT  3.09 0.77 3.29 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.37 0.5 0.65 0.61 ;
      RECT  0.55 0.61 0.65 1.01 ;
      RECT  0.55 1.01 1.45 1.1 ;
      RECT  1.345 0.91 1.45 1.01 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.375 1.14 4.495 1.22 ;
      RECT  4.375 1.22 4.78 1.31 ;
      RECT  4.66 1.31 4.78 1.75 ;
      RECT  0.38 1.44 0.53 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  1.425 1.615 1.595 1.75 ;
      RECT  2.745 1.575 2.895 1.75 ;
      RECT  3.295 1.39 3.445 1.75 ;
      RECT  5.245 1.455 5.395 1.75 ;
      RECT  5.775 1.41 5.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  4.645 0.05 4.815 0.21 ;
      RECT  1.245 0.05 1.395 0.36 ;
      RECT  0.31 0.05 0.46 0.38 ;
      RECT  3.015 0.05 3.165 0.405 ;
      RECT  5.515 0.05 5.635 0.605 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.485 0.245 2.115 0.365 ;
      RECT  1.485 0.365 1.575 0.45 ;
      RECT  0.735 0.215 1.03 0.335 ;
      RECT  0.94 0.335 1.03 0.45 ;
      RECT  0.94 0.45 1.575 0.54 ;
      RECT  4.76 0.3 5.385 0.39 ;
      RECT  5.265 0.39 5.385 0.68 ;
      RECT  4.76 0.39 4.85 0.78 ;
      RECT  5.265 0.68 5.46 0.77 ;
      RECT  5.37 0.77 5.46 0.89 ;
      RECT  4.335 0.665 4.445 0.78 ;
      RECT  4.335 0.78 4.85 0.87 ;
      RECT  5.37 0.89 5.64 1.0 ;
      RECT  5.37 1.0 5.46 1.23 ;
      RECT  4.95 1.23 5.46 1.35 ;
      RECT  3.575 0.32 3.75 0.44 ;
      RECT  3.575 0.44 3.685 1.145 ;
      RECT  2.605 1.145 3.685 1.255 ;
      RECT  3.84 0.325 4.245 0.445 ;
      RECT  4.155 0.445 4.245 0.96 ;
      RECT  4.155 0.96 4.705 1.02 ;
      RECT  4.155 1.02 5.27 1.05 ;
      RECT  5.17 0.88 5.27 1.02 ;
      RECT  4.615 1.05 5.27 1.11 ;
      RECT  4.195 1.05 4.285 1.31 ;
      RECT  3.83 1.31 4.285 1.4 ;
      RECT  3.83 1.4 3.945 1.61 ;
      RECT  1.675 0.51 2.095 0.6 ;
      RECT  1.675 0.6 1.795 0.715 ;
      RECT  1.995 0.6 2.095 1.195 ;
      RECT  1.67 1.195 2.095 1.285 ;
      RECT  1.67 1.285 2.32 1.315 ;
      RECT  1.995 1.315 2.32 1.375 ;
      RECT  2.23 1.375 2.32 1.57 ;
      RECT  2.23 1.57 2.52 1.66 ;
      RECT  2.21 0.2 2.33 0.965 ;
      RECT  2.21 0.965 3.485 1.055 ;
      RECT  3.385 0.725 3.485 0.965 ;
      RECT  2.21 1.055 2.33 1.195 ;
      RECT  3.965 0.535 4.065 0.99 ;
      RECT  0.08 0.19 0.17 1.26 ;
      RECT  0.08 1.26 0.735 1.35 ;
      RECT  0.645 1.35 0.735 1.48 ;
      RECT  0.08 1.35 0.17 1.61 ;
      RECT  0.645 1.48 1.28 1.59 ;
      RECT  0.895 1.215 1.505 1.335 ;
      RECT  1.415 1.335 1.505 1.405 ;
      RECT  1.415 1.405 1.79 1.465 ;
      RECT  1.415 1.465 2.12 1.525 ;
      RECT  1.7 1.525 2.12 1.585 ;
      RECT  2.455 1.35 2.625 1.39 ;
      RECT  2.455 1.39 3.15 1.48 ;
      RECT  3.03 1.48 3.15 1.615 ;
      RECT  4.385 1.405 4.505 1.49 ;
      RECT  4.04 1.49 4.505 1.6 ;
      LAYER M2 ;
      RECT  1.955 0.75 4.105 0.85 ;
      LAYER V1 ;
      RECT  1.995 0.75 2.095 0.85 ;
      RECT  3.965 0.75 4.065 0.85 ;
  END
END SEN_FSDPRBSBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBSBQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBSBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPRBSBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.775 0.555 3.875 1.125 ;
      RECT  3.775 1.125 4.105 1.22 ;
      RECT  1.58 0.845 1.885 0.95 ;
      RECT  1.785 0.95 1.885 1.09 ;
      LAYER M2 ;
      RECT  1.745 0.95 3.915 1.05 ;
      LAYER V1 ;
      RECT  3.775 0.95 3.875 1.05 ;
      RECT  1.785 0.95 1.885 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.115 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.31 5.875 0.505 ;
      RECT  5.75 0.505 5.85 1.11 ;
      RECT  5.75 1.11 6.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.94 0.48 5.05 0.93 ;
      RECT  2.605 0.55 3.075 0.65 ;
      LAYER M2 ;
      RECT  2.895 0.55 4.305 0.65 ;
      RECT  4.205 0.65 4.305 0.75 ;
      RECT  4.205 0.75 5.08 0.85 ;
      LAYER V1 ;
      RECT  4.94 0.75 5.04 0.85 ;
      RECT  2.935 0.55 3.035 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.14 4.45 0.23 ;
      RECT  4.35 0.23 4.45 0.31 ;
      RECT  3.35 0.23 3.45 0.535 ;
      RECT  4.35 0.31 4.65 0.49 ;
      RECT  4.55 0.49 4.65 0.51 ;
      RECT  4.55 0.51 4.67 0.69 ;
      RECT  3.2 0.535 3.45 0.625 ;
      RECT  3.2 0.625 3.29 0.77 ;
      RECT  3.09 0.77 3.29 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.405 0.5 0.65 0.61 ;
      RECT  0.55 0.61 0.65 1.01 ;
      RECT  0.55 1.01 1.45 1.1 ;
      RECT  1.345 0.9 1.45 1.01 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.375 1.14 4.495 1.22 ;
      RECT  4.375 1.22 4.78 1.31 ;
      RECT  4.66 1.31 4.78 1.75 ;
      RECT  0.38 1.44 0.53 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  1.425 1.615 1.595 1.75 ;
      RECT  2.745 1.575 2.895 1.75 ;
      RECT  3.295 1.39 3.445 1.75 ;
      RECT  5.245 1.44 5.39 1.75 ;
      RECT  5.485 1.44 5.635 1.75 ;
      RECT  6.005 1.41 6.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  4.645 0.05 4.815 0.21 ;
      RECT  0.31 0.05 0.46 0.38 ;
      RECT  1.245 0.05 1.395 0.385 ;
      RECT  3.02 0.05 3.17 0.39 ;
      RECT  5.495 0.05 5.615 0.585 ;
      RECT  6.015 0.05 6.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.485 0.245 2.09 0.365 ;
      RECT  1.485 0.365 1.575 0.475 ;
      RECT  0.735 0.215 1.03 0.335 ;
      RECT  0.94 0.335 1.03 0.475 ;
      RECT  0.94 0.475 1.575 0.565 ;
      RECT  4.76 0.3 5.385 0.39 ;
      RECT  5.265 0.39 5.385 0.68 ;
      RECT  4.76 0.39 4.85 0.78 ;
      RECT  5.265 0.68 5.635 0.77 ;
      RECT  5.535 0.77 5.635 1.23 ;
      RECT  4.335 0.64 4.445 0.78 ;
      RECT  4.335 0.78 4.85 0.87 ;
      RECT  4.95 1.23 5.635 1.35 ;
      RECT  3.575 0.32 3.75 0.44 ;
      RECT  3.575 0.44 3.685 1.145 ;
      RECT  2.605 1.145 3.685 1.255 ;
      RECT  3.84 0.325 4.245 0.445 ;
      RECT  4.155 0.445 4.245 0.96 ;
      RECT  4.155 0.96 4.705 1.04 ;
      RECT  4.155 1.04 5.27 1.05 ;
      RECT  5.17 0.88 5.27 1.04 ;
      RECT  4.615 1.05 5.27 1.13 ;
      RECT  4.195 1.05 4.285 1.31 ;
      RECT  3.83 1.31 4.285 1.4 ;
      RECT  3.83 1.4 3.945 1.61 ;
      RECT  1.675 0.51 2.095 0.6 ;
      RECT  1.675 0.6 1.795 0.715 ;
      RECT  1.995 0.6 2.095 1.195 ;
      RECT  1.67 1.195 2.095 1.285 ;
      RECT  1.67 1.285 2.32 1.315 ;
      RECT  1.995 1.315 2.32 1.375 ;
      RECT  2.23 1.375 2.32 1.57 ;
      RECT  2.23 1.57 2.52 1.66 ;
      RECT  2.21 0.2 2.33 0.965 ;
      RECT  2.21 0.965 3.485 1.055 ;
      RECT  3.385 0.755 3.485 0.965 ;
      RECT  2.21 1.055 2.33 1.195 ;
      RECT  3.965 0.535 4.065 0.99 ;
      RECT  0.08 0.19 0.17 1.26 ;
      RECT  0.08 1.26 0.735 1.35 ;
      RECT  0.645 1.35 0.735 1.48 ;
      RECT  0.08 1.35 0.17 1.61 ;
      RECT  0.645 1.48 1.28 1.59 ;
      RECT  0.895 1.215 1.505 1.335 ;
      RECT  1.415 1.335 1.505 1.405 ;
      RECT  1.415 1.405 1.79 1.465 ;
      RECT  1.415 1.465 2.12 1.525 ;
      RECT  1.7 1.525 2.12 1.585 ;
      RECT  2.43 1.35 2.625 1.39 ;
      RECT  2.43 1.39 3.15 1.48 ;
      RECT  3.03 1.48 3.15 1.615 ;
      RECT  4.385 1.405 4.505 1.49 ;
      RECT  4.04 1.49 4.505 1.6 ;
      LAYER M2 ;
      RECT  1.955 0.75 4.105 0.85 ;
      LAYER V1 ;
      RECT  1.995 0.75 2.095 0.85 ;
      RECT  3.965 0.75 4.065 0.85 ;
  END
END SEN_FSDPRBSBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBSBQ_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBSBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDPRBSBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.775 0.555 3.875 1.125 ;
      RECT  3.775 1.125 4.105 1.22 ;
      RECT  1.58 0.845 1.885 0.95 ;
      RECT  1.785 0.95 1.885 1.09 ;
      LAYER M2 ;
      RECT  1.745 0.95 3.915 1.05 ;
      LAYER V1 ;
      RECT  3.775 0.95 3.875 1.05 ;
      RECT  1.785 0.95 1.885 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.115 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.31 5.875 0.51 ;
      RECT  5.75 0.51 6.45 0.69 ;
      RECT  6.35 0.69 6.45 1.11 ;
      RECT  5.75 1.11 6.45 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.94 0.48 5.05 0.9 ;
      RECT  2.605 0.55 3.075 0.65 ;
      LAYER M2 ;
      RECT  2.895 0.55 4.305 0.65 ;
      RECT  4.205 0.65 4.305 0.75 ;
      RECT  4.205 0.75 5.08 0.85 ;
      LAYER V1 ;
      RECT  4.94 0.75 5.04 0.85 ;
      RECT  2.935 0.55 3.035 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.14 4.45 0.23 ;
      RECT  4.35 0.23 4.45 0.31 ;
      RECT  3.35 0.23 3.45 0.525 ;
      RECT  4.35 0.31 4.65 0.49 ;
      RECT  4.55 0.49 4.65 0.51 ;
      RECT  4.55 0.51 4.67 0.69 ;
      RECT  3.2 0.525 3.45 0.615 ;
      RECT  3.2 0.615 3.29 0.77 ;
      RECT  3.09 0.77 3.29 0.875 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.155 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.405 0.5 0.65 0.61 ;
      RECT  0.55 0.61 0.65 1.01 ;
      RECT  0.55 1.01 1.45 1.1 ;
      RECT  1.345 0.9 1.45 1.01 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.375 1.14 4.495 1.22 ;
      RECT  4.375 1.22 4.78 1.31 ;
      RECT  4.66 1.31 4.78 1.75 ;
      RECT  0.365 1.44 0.515 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.425 1.615 1.595 1.75 ;
      RECT  2.745 1.575 2.895 1.75 ;
      RECT  3.295 1.39 3.445 1.75 ;
      RECT  5.245 1.44 5.39 1.75 ;
      RECT  5.485 1.44 5.635 1.75 ;
      RECT  6.015 1.415 6.135 1.75 ;
      RECT  6.58 1.21 6.7 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  4.645 0.05 4.815 0.21 ;
      RECT  1.245 0.05 1.395 0.385 ;
      RECT  3.02 0.05 3.17 0.39 ;
      RECT  0.31 0.05 0.46 0.405 ;
      RECT  6.0 0.05 6.15 0.41 ;
      RECT  5.495 0.05 5.615 0.585 ;
      RECT  6.58 0.05 6.7 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.485 0.245 2.115 0.365 ;
      RECT  1.485 0.365 1.575 0.475 ;
      RECT  0.735 0.215 1.03 0.335 ;
      RECT  0.94 0.335 1.03 0.475 ;
      RECT  0.94 0.475 1.575 0.565 ;
      RECT  4.76 0.3 5.385 0.39 ;
      RECT  5.265 0.39 5.385 0.68 ;
      RECT  4.76 0.39 4.85 0.78 ;
      RECT  5.265 0.68 5.635 0.77 ;
      RECT  5.535 0.77 5.635 0.785 ;
      RECT  4.335 0.64 4.445 0.78 ;
      RECT  4.335 0.78 4.85 0.87 ;
      RECT  5.535 0.785 6.205 0.895 ;
      RECT  5.535 0.895 5.635 1.23 ;
      RECT  4.95 1.23 5.635 1.35 ;
      RECT  3.575 0.32 3.75 0.44 ;
      RECT  3.575 0.44 3.685 1.145 ;
      RECT  2.59 1.145 3.685 1.255 ;
      RECT  3.84 0.325 4.245 0.445 ;
      RECT  4.155 0.445 4.245 0.96 ;
      RECT  4.155 0.96 4.705 1.01 ;
      RECT  4.155 1.01 5.27 1.05 ;
      RECT  5.17 0.86 5.27 1.01 ;
      RECT  4.615 1.05 5.27 1.1 ;
      RECT  4.195 1.05 4.285 1.31 ;
      RECT  3.83 1.31 4.285 1.4 ;
      RECT  3.83 1.4 3.945 1.61 ;
      RECT  1.675 0.51 2.095 0.6 ;
      RECT  1.675 0.6 1.795 0.715 ;
      RECT  1.995 0.6 2.095 1.195 ;
      RECT  1.695 1.195 2.095 1.285 ;
      RECT  1.695 1.285 2.3 1.315 ;
      RECT  1.995 1.315 2.3 1.375 ;
      RECT  2.21 1.375 2.3 1.57 ;
      RECT  2.21 1.57 2.52 1.66 ;
      RECT  2.21 0.23 2.33 0.965 ;
      RECT  2.21 0.965 3.485 1.055 ;
      RECT  3.385 0.725 3.485 0.965 ;
      RECT  2.21 1.055 2.33 1.195 ;
      RECT  3.965 0.535 4.065 1.015 ;
      RECT  0.08 0.2 0.17 1.26 ;
      RECT  0.08 1.26 0.735 1.35 ;
      RECT  0.645 1.35 0.735 1.48 ;
      RECT  0.08 1.35 0.17 1.61 ;
      RECT  0.645 1.48 1.28 1.59 ;
      RECT  0.89 1.215 1.505 1.335 ;
      RECT  1.415 1.335 1.505 1.405 ;
      RECT  1.415 1.405 1.79 1.465 ;
      RECT  1.415 1.465 2.12 1.525 ;
      RECT  1.7 1.525 2.12 1.585 ;
      RECT  2.43 1.35 2.625 1.39 ;
      RECT  2.43 1.39 3.15 1.48 ;
      RECT  3.03 1.48 3.15 1.615 ;
      RECT  4.385 1.405 4.505 1.49 ;
      RECT  4.04 1.49 4.505 1.6 ;
      LAYER M2 ;
      RECT  1.955 0.75 4.105 0.85 ;
      LAYER V1 ;
      RECT  1.995 0.75 2.095 0.85 ;
      RECT  3.965 0.75 4.065 0.85 ;
  END
END SEN_FSDPRBSBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBSBQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear/set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBSBQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDPRBSBQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.59 0.74 4.69 1.19 ;
      RECT  1.765 0.77 1.91 1.105 ;
      LAYER M2 ;
      RECT  1.77 0.95 4.73 1.05 ;
      LAYER V1 ;
      RECT  4.59 0.95 4.69 1.05 ;
      RECT  1.81 0.95 1.91 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0762 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.51 0.31 6.65 0.49 ;
      RECT  6.55 0.49 6.65 1.31 ;
      RECT  6.495 1.31 6.65 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.46 0.495 5.66 0.665 ;
      RECT  5.54 0.665 5.66 0.89 ;
      RECT  3.43 0.51 3.66 0.69 ;
      RECT  3.43 0.69 3.52 0.925 ;
      LAYER M2 ;
      RECT  3.52 0.55 5.69 0.65 ;
      LAYER V1 ;
      RECT  5.55 0.55 5.65 0.65 ;
      RECT  3.56 0.55 3.66 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.14 5.52 0.23 ;
      RECT  5.43 0.23 5.52 0.315 ;
      RECT  3.75 0.23 3.84 0.8 ;
      RECT  5.43 0.315 5.84 0.405 ;
      RECT  5.75 0.405 5.84 0.51 ;
      RECT  5.75 0.51 6.05 0.69 ;
      RECT  5.95 0.69 6.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.057 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.51 0.65 0.6 ;
      RECT  0.55 0.6 0.65 1.005 ;
      RECT  0.55 1.005 1.495 1.095 ;
      RECT  1.405 1.095 1.495 1.175 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.3 7.13 0.69 ;
      RECT  7.03 0.69 7.13 1.11 ;
      RECT  6.95 1.11 7.13 1.49 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  5.4 1.16 5.84 1.25 ;
      RECT  5.72 1.25 5.84 1.75 ;
      RECT  0.385 1.44 0.525 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  1.465 1.615 1.635 1.75 ;
      RECT  2.03 1.615 2.2 1.75 ;
      RECT  3.285 1.47 3.455 1.75 ;
      RECT  3.84 1.43 4.01 1.75 ;
      RECT  6.225 1.6 6.395 1.75 ;
      RECT  6.755 1.215 6.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  5.61 0.05 5.725 0.225 ;
      RECT  1.27 0.05 1.44 0.305 ;
      RECT  1.81 0.05 1.93 0.305 ;
      RECT  0.325 0.05 0.445 0.385 ;
      RECT  3.515 0.05 3.635 0.385 ;
      RECT  6.755 0.05 6.86 0.57 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  2.02 0.18 2.62 0.27 ;
      RECT  2.02 0.27 2.11 0.395 ;
      RECT  2.5 0.27 2.62 0.43 ;
      RECT  0.745 0.24 1.15 0.36 ;
      RECT  1.06 0.36 1.15 0.395 ;
      RECT  1.06 0.395 2.11 0.485 ;
      RECT  1.35 0.485 1.44 0.825 ;
      RECT  1.35 0.825 1.675 0.915 ;
      RECT  1.585 0.915 1.675 1.305 ;
      RECT  0.925 1.305 1.675 1.395 ;
      RECT  1.585 1.395 1.675 1.42 ;
      RECT  1.585 1.42 2.68 1.525 ;
      RECT  2.76 0.22 2.925 0.4 ;
      RECT  2.825 0.4 2.925 1.015 ;
      RECT  2.75 1.015 2.925 1.135 ;
      RECT  3.93 0.35 4.11 0.45 ;
      RECT  3.985 0.45 4.11 0.8 ;
      RECT  4.655 0.335 5.34 0.45 ;
      RECT  4.41 0.34 4.555 0.51 ;
      RECT  4.41 0.51 4.5 1.25 ;
      RECT  3.015 0.2 3.14 0.395 ;
      RECT  3.015 0.395 3.105 1.25 ;
      RECT  3.015 1.25 4.5 1.31 ;
      RECT  3.015 1.31 4.795 1.34 ;
      RECT  3.015 1.34 3.69 1.355 ;
      RECT  4.41 1.34 4.795 1.405 ;
      RECT  3.57 1.355 3.69 1.61 ;
      RECT  4.625 1.405 4.795 1.43 ;
      RECT  1.53 0.575 2.1 0.68 ;
      RECT  2.0 0.68 2.1 1.235 ;
      RECT  1.765 1.235 2.925 1.325 ;
      RECT  2.835 1.325 2.925 1.525 ;
      RECT  2.835 1.525 3.08 1.625 ;
      RECT  4.78 0.59 4.925 0.76 ;
      RECT  4.78 0.76 4.885 1.11 ;
      RECT  4.78 1.11 4.95 1.2 ;
      RECT  6.745 0.78 6.94 0.96 ;
      RECT  6.745 0.96 6.845 1.11 ;
      RECT  2.2 0.36 2.305 0.97 ;
      RECT  2.2 0.97 2.66 1.06 ;
      RECT  2.56 0.89 2.66 0.97 ;
      RECT  2.2 1.06 2.425 1.125 ;
      RECT  5.31 0.75 5.41 0.98 ;
      RECT  5.31 0.98 6.23 1.07 ;
      RECT  6.14 0.185 6.23 0.98 ;
      RECT  5.98 1.07 6.1 1.595 ;
      RECT  3.195 0.725 3.285 1.015 ;
      RECT  3.195 1.015 4.29 1.13 ;
      RECT  4.2 0.32 4.29 1.015 ;
      RECT  5.065 0.585 5.165 1.16 ;
      RECT  5.065 1.16 5.305 1.25 ;
      RECT  5.195 1.25 5.305 1.46 ;
      RECT  5.195 1.46 5.63 1.55 ;
      RECT  6.32 0.29 6.42 1.16 ;
      RECT  6.215 1.16 6.42 1.255 ;
      RECT  6.215 1.255 6.315 1.49 ;
      RECT  0.08 0.2 0.17 1.26 ;
      RECT  0.08 1.26 0.835 1.35 ;
      RECT  0.745 1.35 0.835 1.565 ;
      RECT  0.08 1.35 0.17 1.61 ;
      RECT  0.745 1.565 1.31 1.66 ;
      RECT  4.91 1.345 5.1 1.515 ;
      RECT  4.91 1.515 5.01 1.54 ;
      RECT  4.34 1.495 4.535 1.54 ;
      RECT  4.34 1.54 5.01 1.63 ;
      LAYER M2 ;
      RECT  2.785 0.35 4.11 0.45 ;
      RECT  5.16 0.35 6.46 0.45 ;
      RECT  1.96 0.75 4.925 0.85 ;
      RECT  5.025 0.95 6.885 1.05 ;
      RECT  4.88 1.35 6.355 1.45 ;
      LAYER V1 ;
      RECT  2.825 0.35 2.925 0.45 ;
      RECT  3.97 0.35 4.07 0.45 ;
      RECT  5.2 0.35 5.3 0.45 ;
      RECT  6.32 0.35 6.42 0.45 ;
      RECT  2.0 0.75 2.1 0.85 ;
      RECT  4.785 0.75 4.885 0.85 ;
      RECT  5.065 0.95 5.165 1.05 ;
      RECT  6.745 0.95 6.845 1.05 ;
      RECT  4.96 1.35 5.06 1.45 ;
      RECT  6.215 1.35 6.315 1.45 ;
  END
END SEN_FSDPRBSBQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBSBQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear/set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBSBQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDPRBSBQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.11 0.95 6.29 1.265 ;
      RECT  5.19 0.735 5.63 0.845 ;
      RECT  5.53 0.845 5.63 1.09 ;
      LAYER M2 ;
      RECT  5.49 0.95 6.29 1.05 ;
      LAYER V1 ;
      RECT  6.15 0.95 6.25 1.05 ;
      RECT  5.53 0.95 5.63 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0981 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.73 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0846 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.9 0.31 8.05 0.49 ;
      RECT  7.95 0.49 8.05 1.11 ;
      RECT  7.895 1.11 8.05 1.29 ;
    END
    ANTENNADIFFAREA 0.218 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.615 0.87 6.715 1.29 ;
      RECT  3.63 1.12 3.97 1.25 ;
      LAYER M2 ;
      RECT  3.79 1.15 6.755 1.25 ;
      LAYER V1 ;
      RECT  6.615 1.15 6.715 1.25 ;
      RECT  3.83 1.15 3.93 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0846 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.015 0.495 7.115 1.04 ;
      RECT  3.895 0.51 4.105 0.85 ;
      LAYER M2 ;
      RECT  3.965 0.55 7.155 0.65 ;
      LAYER V1 ;
      RECT  7.015 0.55 7.115 0.65 ;
      RECT  4.005 0.55 4.105 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.505 1.33 0.595 ;
      RECT  1.24 0.595 1.33 0.63 ;
      RECT  0.35 0.595 0.45 1.12 ;
      RECT  1.24 0.63 1.405 0.8 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.087 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.685 1.115 0.855 ;
      RECT  0.95 0.855 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.41 0.29 8.53 0.46 ;
      RECT  8.15 0.46 8.53 0.55 ;
      RECT  8.15 0.55 8.25 1.245 ;
      RECT  8.15 1.245 8.53 1.335 ;
      RECT  8.41 1.335 8.53 1.51 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.415 0.455 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.855 1.63 1.025 1.75 ;
      RECT  3.285 1.54 3.405 1.75 ;
      RECT  3.835 1.52 3.955 1.75 ;
      RECT  4.35 1.48 4.52 1.75 ;
      RECT  5.195 1.44 5.315 1.75 ;
      RECT  6.47 1.615 6.64 1.75 ;
      RECT  7.015 1.395 7.135 1.75 ;
      RECT  7.63 1.39 7.75 1.75 ;
      RECT  8.15 1.44 8.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  0.855 0.05 1.025 0.17 ;
      RECT  6.775 0.05 6.915 0.225 ;
      RECT  8.15 0.05 8.27 0.345 ;
      RECT  3.27 0.05 3.44 0.35 ;
      RECT  7.625 0.05 7.745 0.36 ;
      RECT  0.335 0.05 0.455 0.38 ;
      RECT  3.82 0.05 3.96 0.385 ;
      RECT  5.445 0.05 5.585 0.39 ;
      RECT  4.925 0.05 5.045 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.115 0.14 1.785 0.23 ;
      RECT  1.115 0.23 1.205 0.285 ;
      RECT  1.665 0.23 1.785 0.36 ;
      RECT  0.545 0.285 1.205 0.375 ;
      RECT  5.93 0.14 6.685 0.23 ;
      RECT  6.595 0.23 6.685 0.315 ;
      RECT  5.93 0.23 6.07 0.385 ;
      RECT  6.595 0.315 7.295 0.405 ;
      RECT  5.93 0.385 6.02 1.395 ;
      RECT  7.205 0.405 7.295 0.79 ;
      RECT  7.205 0.79 7.605 0.89 ;
      RECT  5.93 1.395 6.07 1.48 ;
      RECT  5.42 1.48 6.07 1.57 ;
      RECT  4.61 0.235 4.785 0.405 ;
      RECT  4.61 0.405 4.7 0.91 ;
      RECT  4.61 0.91 4.75 1.2 ;
      RECT  6.175 0.32 6.395 0.41 ;
      RECT  6.175 0.41 6.265 0.75 ;
      RECT  6.175 0.75 6.525 0.85 ;
      RECT  6.435 0.85 6.525 1.38 ;
      RECT  6.2 1.38 6.91 1.5 ;
      RECT  1.42 0.32 1.525 0.45 ;
      RECT  1.42 0.45 2.1 0.54 ;
      RECT  1.84 0.54 2.1 0.555 ;
      RECT  1.84 0.555 1.93 1.205 ;
      RECT  1.42 1.205 2.045 1.295 ;
      RECT  1.42 1.295 1.525 1.375 ;
      RECT  1.925 1.295 2.045 1.385 ;
      RECT  1.925 1.385 2.645 1.505 ;
      RECT  7.385 0.2 7.49 0.45 ;
      RECT  7.385 0.45 7.805 0.54 ;
      RECT  7.715 0.54 7.805 1.13 ;
      RECT  6.355 0.54 6.895 0.65 ;
      RECT  6.805 0.65 6.895 1.13 ;
      RECT  6.805 1.13 7.805 1.22 ;
      RECT  7.275 1.22 7.395 1.615 ;
      RECT  5.19 0.27 5.31 0.555 ;
      RECT  4.84 0.555 5.31 0.645 ;
      RECT  4.84 0.645 4.94 1.0 ;
      RECT  4.84 1.0 5.03 1.17 ;
      RECT  2.725 0.465 3.725 0.585 ;
      RECT  4.195 0.29 4.295 0.73 ;
      RECT  4.195 0.73 4.325 0.8 ;
      RECT  4.235 0.8 4.325 0.9 ;
      RECT  3.24 0.87 3.515 0.94 ;
      RECT  3.24 0.94 4.15 0.97 ;
      RECT  3.425 0.97 4.15 1.03 ;
      RECT  4.06 1.03 4.15 1.07 ;
      RECT  4.06 1.07 4.52 1.16 ;
      RECT  4.43 0.205 4.52 1.07 ;
      RECT  2.655 0.91 2.94 1.09 ;
      RECT  8.35 0.67 8.45 1.09 ;
      RECT  1.24 0.915 1.345 1.115 ;
      RECT  1.24 1.115 1.33 1.21 ;
      RECT  0.065 0.22 0.185 1.21 ;
      RECT  0.065 1.21 1.33 1.3 ;
      RECT  0.715 0.685 0.805 1.21 ;
      RECT  0.065 1.3 0.185 1.59 ;
      RECT  2.03 0.695 2.13 1.115 ;
      RECT  2.22 0.2 2.32 1.18 ;
      RECT  2.22 1.18 2.865 1.27 ;
      RECT  2.745 1.27 2.865 1.425 ;
      RECT  5.72 0.41 5.825 1.26 ;
      RECT  4.82 1.26 5.825 1.29 ;
      RECT  4.2 1.29 5.825 1.34 ;
      RECT  2.47 0.215 3.18 0.335 ;
      RECT  2.47 0.335 2.56 0.7 ;
      RECT  2.47 0.7 3.135 0.79 ;
      RECT  3.03 0.79 3.135 1.34 ;
      RECT  3.03 1.34 5.825 1.35 ;
      RECT  3.03 1.35 4.89 1.39 ;
      RECT  3.03 1.39 4.275 1.43 ;
      RECT  3.03 1.43 3.675 1.45 ;
      RECT  3.555 1.45 3.675 1.58 ;
      RECT  0.545 1.43 1.19 1.465 ;
      RECT  0.545 1.465 1.835 1.52 ;
      RECT  1.09 1.52 1.835 1.555 ;
      LAYER M2 ;
      RECT  2.18 0.35 4.335 0.45 ;
      RECT  1.99 0.75 4.98 0.85 ;
      RECT  6.345 0.75 8.49 0.85 ;
      RECT  2.8 0.95 4.75 1.05 ;
      LAYER V1 ;
      RECT  2.22 0.35 2.32 0.45 ;
      RECT  4.195 0.35 4.295 0.45 ;
      RECT  2.03 0.75 2.13 0.85 ;
      RECT  4.84 0.75 4.94 0.85 ;
      RECT  6.385 0.75 6.485 0.85 ;
      RECT  8.35 0.75 8.45 0.85 ;
      RECT  2.84 0.95 2.94 1.05 ;
      RECT  4.61 0.95 4.71 1.05 ;
  END
END SEN_FSDPRBSBQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBSBQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear/set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBSBQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDPRBSBQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 0.31 8.65 0.71 ;
      RECT  8.245 0.71 8.65 0.815 ;
      LAYER M2 ;
      RECT  8.51 0.35 9.255 0.45 ;
      LAYER V1 ;
      RECT  8.55 0.35 8.65 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1266 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.815 ;
      RECT  0.55 0.815 1.25 0.925 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1092 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  11.235 0.51 11.86 0.69 ;
      RECT  11.75 0.69 11.86 1.11 ;
      RECT  11.155 1.03 11.54 1.11 ;
      RECT  11.155 1.11 11.86 1.12 ;
      RECT  11.45 1.12 11.86 1.29 ;
    END
    ANTENNADIFFAREA 0.464 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.095 0.645 9.195 0.75 ;
      RECT  8.76 0.75 9.195 0.85 ;
      RECT  8.76 0.85 8.85 1.02 ;
      RECT  8.355 0.95 8.445 1.02 ;
      RECT  8.355 1.02 8.85 1.12 ;
      RECT  5.955 0.675 6.445 0.85 ;
      LAYER M2 ;
      RECT  6.065 0.75 9.11 0.85 ;
      LAYER V1 ;
      RECT  8.97 0.75 9.07 0.85 ;
      RECT  6.105 0.75 6.205 0.85 ;
      RECT  6.305 0.75 6.405 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1197 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.19 0.89 10.29 1.11 ;
      RECT  10.19 1.11 10.45 1.29 ;
      RECT  4.35 0.84 4.625 1.05 ;
      LAYER M2 ;
      RECT  4.445 0.95 10.33 1.05 ;
      LAYER V1 ;
      RECT  10.19 0.95 10.29 1.05 ;
      RECT  4.485 0.95 4.585 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.078 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.275 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1035 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.65 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.01 0.34 10.1 0.51 ;
      RECT  10.01 0.51 10.65 0.69 ;
      RECT  10.55 0.31 10.65 0.51 ;
      RECT  10.01 0.69 10.1 1.11 ;
      RECT  9.855 1.11 10.1 1.29 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.4 0.445 1.75 ;
      RECT  0.0 1.75 12.2 1.85 ;
      RECT  0.845 1.39 0.965 1.75 ;
      RECT  2.585 1.48 2.705 1.75 ;
      RECT  4.495 1.63 4.665 1.75 ;
      RECT  5.08 1.325 5.185 1.75 ;
      RECT  5.295 1.48 5.465 1.75 ;
      RECT  5.815 1.48 5.985 1.75 ;
      RECT  6.335 1.48 6.505 1.75 ;
      RECT  7.64 1.48 7.81 1.75 ;
      RECT  8.185 1.44 8.305 1.75 ;
      RECT  8.705 1.41 8.81 1.75 ;
      RECT  10.085 1.615 10.255 1.75 ;
      RECT  10.92 1.43 11.04 1.75 ;
      RECT  11.44 1.38 11.56 1.75 ;
      RECT  12.015 1.21 12.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.2 0.05 ;
      RECT  5.94 0.05 6.06 0.225 ;
      RECT  6.48 0.05 6.6 0.225 ;
      RECT  8.37 0.05 8.49 0.24 ;
      RECT  1.8 0.05 1.915 0.375 ;
      RECT  4.365 0.05 4.485 0.375 ;
      RECT  2.815 0.05 2.935 0.385 ;
      RECT  0.085 0.05 0.225 0.39 ;
      RECT  10.255 0.05 10.375 0.42 ;
      RECT  11.495 0.05 11.615 0.42 ;
      RECT  8.985 0.05 9.105 0.445 ;
      RECT  10.975 0.05 11.095 0.56 ;
      RECT  12.015 0.05 12.135 0.59 ;
      RECT  2.305 0.05 2.41 0.615 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.1 0.15 3.96 0.245 ;
      RECT  3.1 0.245 3.19 1.015 ;
      RECT  3.1 1.015 3.325 1.065 ;
      RECT  2.815 1.065 3.325 1.185 ;
      RECT  9.285 0.16 9.89 0.25 ;
      RECT  9.285 0.25 9.375 1.035 ;
      RECT  9.15 1.035 9.375 1.125 ;
      RECT  9.15 1.125 9.265 1.35 ;
      RECT  9.085 1.35 9.265 1.45 ;
      RECT  4.78 0.165 5.525 0.255 ;
      RECT  4.78 0.255 4.9 0.465 ;
      RECT  5.435 0.255 5.525 0.475 ;
      RECT  4.105 0.31 4.225 0.465 ;
      RECT  4.105 0.465 4.9 0.555 ;
      RECT  7.545 0.235 8.24 0.325 ;
      RECT  7.545 0.325 7.635 0.495 ;
      RECT  5.615 0.495 7.635 0.565 ;
      RECT  5.37 0.565 7.635 0.585 ;
      RECT  5.37 0.585 5.705 0.655 ;
      RECT  7.025 0.585 7.115 1.04 ;
      RECT  5.37 0.655 5.47 0.91 ;
      RECT  6.715 1.04 7.115 1.13 ;
      RECT  6.715 1.13 6.805 1.29 ;
      RECT  5.53 1.29 6.805 1.39 ;
      RECT  6.635 1.39 6.805 1.49 ;
      RECT  6.635 1.49 7.31 1.58 ;
      RECT  0.55 0.28 1.01 0.38 ;
      RECT  0.83 0.38 1.01 0.45 ;
      RECT  1.1 0.26 1.71 0.38 ;
      RECT  1.62 0.38 1.71 0.48 ;
      RECT  1.62 0.48 2.215 0.585 ;
      RECT  5.635 0.315 7.44 0.405 ;
      RECT  7.765 0.42 7.935 0.51 ;
      RECT  7.765 0.51 7.855 0.675 ;
      RECT  7.205 0.675 7.855 0.765 ;
      RECT  7.205 0.765 7.295 1.22 ;
      RECT  6.895 1.22 7.295 1.25 ;
      RECT  6.895 1.25 7.55 1.34 ;
      RECT  6.895 1.34 6.985 1.39 ;
      RECT  7.45 1.34 7.55 1.51 ;
      RECT  2.5 0.19 2.66 0.55 ;
      RECT  8.74 0.21 8.83 0.55 ;
      RECT  8.74 0.55 8.99 0.65 ;
      RECT  3.35 0.43 3.52 0.6 ;
      RECT  3.43 0.6 3.52 1.3 ;
      RECT  0.805 0.54 1.53 0.63 ;
      RECT  1.44 0.63 1.53 0.69 ;
      RECT  1.44 0.69 2.255 0.78 ;
      RECT  1.44 0.78 1.53 1.105 ;
      RECT  2.165 0.78 2.255 1.18 ;
      RECT  1.44 1.105 1.655 1.195 ;
      RECT  2.06 1.18 2.255 1.3 ;
      RECT  2.06 1.3 3.52 1.39 ;
      RECT  9.66 0.36 9.78 0.725 ;
      RECT  10.92 0.795 11.645 0.89 ;
      RECT  10.92 0.89 11.01 1.24 ;
      RECT  10.92 1.24 11.25 1.33 ;
      RECT  11.15 1.33 11.25 1.51 ;
      RECT  4.72 0.785 4.98 0.895 ;
      RECT  4.72 0.895 4.81 1.27 ;
      RECT  3.61 0.405 3.715 1.27 ;
      RECT  3.61 1.27 4.81 1.36 ;
      RECT  3.61 1.36 3.7 1.48 ;
      RECT  3.065 1.48 3.7 1.57 ;
      RECT  9.48 0.34 9.57 0.895 ;
      RECT  9.48 0.895 9.92 0.985 ;
      RECT  9.83 0.815 9.92 0.895 ;
      RECT  9.48 0.985 9.57 1.215 ;
      RECT  9.425 1.215 9.57 1.305 ;
      RECT  9.425 1.305 9.515 1.54 ;
      RECT  8.445 1.23 8.995 1.32 ;
      RECT  8.905 1.32 8.995 1.54 ;
      RECT  8.445 1.32 8.565 1.61 ;
      RECT  8.905 1.54 9.515 1.63 ;
      RECT  2.91 0.51 3.01 0.935 ;
      RECT  6.535 0.77 6.935 0.95 ;
      RECT  6.535 0.95 6.625 1.0 ;
      RECT  5.59 1.0 6.625 1.1 ;
      RECT  5.59 1.1 5.68 1.11 ;
      RECT  5.16 0.345 5.28 1.105 ;
      RECT  4.9 1.105 5.28 1.11 ;
      RECT  4.9 1.11 5.68 1.2 ;
      RECT  4.9 1.2 4.99 1.45 ;
      RECT  4.185 1.45 4.99 1.54 ;
      RECT  8.025 0.49 8.125 1.02 ;
      RECT  7.385 1.02 8.125 1.11 ;
      RECT  7.385 1.11 8.045 1.12 ;
      RECT  7.925 1.12 8.045 1.59 ;
      RECT  3.855 0.385 3.975 1.035 ;
      RECT  3.855 1.035 4.25 1.155 ;
      RECT  4.15 0.69 4.25 1.035 ;
      RECT  1.88 0.87 2.05 1.04 ;
      RECT  1.88 1.04 1.97 1.285 ;
      RECT  0.37 0.165 0.46 1.03 ;
      RECT  0.37 1.03 1.35 1.12 ;
      RECT  0.37 1.12 0.46 1.22 ;
      RECT  1.26 1.12 1.35 1.285 ;
      RECT  0.065 1.22 0.46 1.31 ;
      RECT  1.26 1.285 1.97 1.375 ;
      RECT  0.065 1.31 0.185 1.61 ;
      RECT  0.585 1.21 1.17 1.3 ;
      RECT  0.585 1.3 0.705 1.405 ;
      RECT  1.08 1.3 1.17 1.465 ;
      RECT  1.08 1.465 1.93 1.57 ;
      RECT  10.74 0.25 10.83 1.405 ;
      RECT  9.605 1.405 10.83 1.5 ;
      RECT  9.605 1.5 9.695 1.605 ;
      LAYER M2 ;
      RECT  0.83 0.35 2.64 0.45 ;
      RECT  2.87 0.55 9.8 0.65 ;
      RECT  4.11 0.75 5.51 0.85 ;
      RECT  7.41 1.35 11.29 1.45 ;
      LAYER V1 ;
      RECT  0.87 0.35 0.97 0.45 ;
      RECT  2.5 0.35 2.6 0.45 ;
      RECT  2.91 0.55 3.01 0.65 ;
      RECT  8.025 0.55 8.125 0.65 ;
      RECT  8.78 0.55 8.88 0.65 ;
      RECT  9.66 0.55 9.76 0.65 ;
      RECT  4.15 0.75 4.25 0.85 ;
      RECT  5.37 0.75 5.47 0.85 ;
      RECT  7.45 1.35 7.55 1.45 ;
      RECT  9.125 1.35 9.225 1.45 ;
      RECT  11.15 1.35 11.25 1.45 ;
  END
END SEN_FSDPRBSBQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBSBQO_6
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear/set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBSBQO_6
  CLASS CORE ;
  FOREIGN SEN_FSDPRBSBQO_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.35 0.31 9.45 0.77 ;
      RECT  9.14 0.77 9.62 0.865 ;
      LAYER M2 ;
      RECT  9.31 0.35 10.29 0.45 ;
      LAYER V1 ;
      RECT  9.35 0.35 9.45 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1491 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.785 ;
      RECT  0.55 0.785 1.28 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  12.035 0.51 13.25 0.69 ;
      RECT  12.92 0.69 13.05 1.11 ;
      RECT  12.035 1.11 13.25 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.92 0.71 10.02 0.97 ;
      RECT  9.345 0.97 10.02 1.06 ;
      RECT  9.345 1.06 9.435 1.2 ;
      RECT  6.15 0.75 7.295 0.895 ;
      LAYER M2 ;
      RECT  6.915 0.75 10.06 0.85 ;
      LAYER V1 ;
      RECT  9.92 0.75 10.02 0.85 ;
      RECT  6.955 0.75 7.055 0.85 ;
      RECT  7.155 0.75 7.255 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1512 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.15 0.71 11.275 1.195 ;
      RECT  4.605 0.91 5.03 1.09 ;
      LAYER M2 ;
      RECT  4.89 0.95 11.315 1.05 ;
      LAYER V1 ;
      RECT  11.175 0.95 11.275 1.05 ;
      RECT  4.93 0.95 5.03 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0876 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.255 0.975 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1164 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.65 0.91 ;
      RECT  2.35 0.91 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.75 0.385 10.985 0.505 ;
      RECT  10.75 0.505 10.85 1.115 ;
      RECT  10.695 1.115 10.85 1.285 ;
    END
    ANTENNADIFFAREA 0.105 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  9.705 1.175 9.825 1.3 ;
      RECT  9.175 1.3 9.825 1.39 ;
      RECT  9.175 1.39 9.295 1.75 ;
      RECT  0.325 1.375 0.445 1.75 ;
      RECT  0.0 1.75 13.6 1.85 ;
      RECT  0.86 1.44 1.0 1.75 ;
      RECT  2.5 1.46 2.67 1.75 ;
      RECT  4.485 1.395 4.605 1.75 ;
      RECT  4.99 1.615 5.16 1.75 ;
      RECT  5.545 1.215 5.665 1.75 ;
      RECT  6.065 1.455 6.185 1.75 ;
      RECT  6.585 1.455 6.705 1.75 ;
      RECT  7.23 1.455 7.35 1.75 ;
      RECT  10.94 1.63 11.11 1.75 ;
      RECT  11.75 1.435 11.92 1.75 ;
      RECT  12.295 1.38 12.415 1.75 ;
      RECT  12.815 1.39 12.935 1.75 ;
      RECT  13.36 1.21 13.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 13.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
      RECT  11.85 1.75 11.95 1.85 ;
      RECT  12.45 1.75 12.55 1.85 ;
      RECT  13.05 1.75 13.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 13.6 0.05 ;
      RECT  6.37 0.05 6.54 0.22 ;
      RECT  6.91 0.05 7.08 0.22 ;
      RECT  9.26 0.05 9.38 0.22 ;
      RECT  1.75 0.05 1.855 0.365 ;
      RECT  12.295 0.05 12.415 0.38 ;
      RECT  12.815 0.05 12.935 0.38 ;
      RECT  4.565 0.05 4.685 0.385 ;
      RECT  0.07 0.05 0.205 0.39 ;
      RECT  2.755 0.05 2.895 0.39 ;
      RECT  5.85 0.05 5.97 0.415 ;
      RECT  11.075 0.05 11.195 0.42 ;
      RECT  9.805 0.05 9.925 0.485 ;
      RECT  11.775 0.05 11.895 0.585 ;
      RECT  2.255 0.05 2.36 0.59 ;
      RECT  13.36 0.05 13.48 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 13.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
      RECT  11.85 -0.05 11.95 0.05 ;
      RECT  12.45 -0.05 12.55 0.05 ;
      RECT  13.05 -0.05 13.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.04 0.16 4.125 0.25 ;
      RECT  3.04 0.25 3.145 1.0 ;
      RECT  3.04 1.0 3.345 1.06 ;
      RECT  2.77 1.06 3.345 1.17 ;
      RECT  2.77 1.17 2.94 1.19 ;
      RECT  10.11 0.145 10.735 0.255 ;
      RECT  10.11 0.255 10.21 1.245 ;
      RECT  9.945 1.245 10.21 1.365 ;
      RECT  8.51 0.19 9.135 0.28 ;
      RECT  9.015 0.28 9.135 0.39 ;
      RECT  8.51 0.28 8.615 0.545 ;
      RECT  5.48 0.545 8.615 0.635 ;
      RECT  5.48 0.635 7.73 0.66 ;
      RECT  5.48 0.66 5.58 0.91 ;
      RECT  7.625 0.66 7.73 1.245 ;
      RECT  5.755 1.245 7.73 1.365 ;
      RECT  7.61 1.365 7.73 1.48 ;
      RECT  7.61 1.48 8.82 1.595 ;
      RECT  4.94 0.2 5.715 0.32 ;
      RECT  4.94 0.32 5.06 0.485 ;
      RECT  4.28 0.485 5.06 0.605 ;
      RECT  0.56 0.235 1.0 0.34 ;
      RECT  0.82 0.34 1.0 0.45 ;
      RECT  1.09 0.22 1.66 0.34 ;
      RECT  1.57 0.34 1.66 0.48 ;
      RECT  1.57 0.48 2.165 0.6 ;
      RECT  2.45 0.235 2.61 0.42 ;
      RECT  2.45 0.42 2.55 0.59 ;
      RECT  6.08 0.335 8.415 0.455 ;
      RECT  3.25 0.365 3.915 0.47 ;
      RECT  3.81 0.47 3.915 1.215 ;
      RECT  3.81 1.215 5.21 1.305 ;
      RECT  5.12 0.89 5.21 1.215 ;
      RECT  3.81 1.305 4.105 1.31 ;
      RECT  3.985 1.31 4.105 1.48 ;
      RECT  3.255 1.48 4.105 1.585 ;
      RECT  9.56 0.195 9.66 0.55 ;
      RECT  9.56 0.55 9.74 0.65 ;
      RECT  3.485 0.575 3.72 0.68 ;
      RECT  3.63 0.68 3.72 1.28 ;
      RECT  1.39 0.48 1.48 0.54 ;
      RECT  0.805 0.54 1.48 0.665 ;
      RECT  1.39 0.665 1.48 0.715 ;
      RECT  1.39 0.715 2.25 0.805 ;
      RECT  1.465 0.805 1.585 1.165 ;
      RECT  2.16 0.805 2.25 1.24 ;
      RECT  1.97 1.24 2.25 1.28 ;
      RECT  1.97 1.28 3.72 1.37 ;
      RECT  3.045 1.37 3.72 1.39 ;
      RECT  3.045 1.39 3.165 1.58 ;
      RECT  8.755 0.37 8.86 0.725 ;
      RECT  8.35 0.725 8.86 0.815 ;
      RECT  8.35 0.815 8.45 1.27 ;
      RECT  7.845 1.27 8.56 1.39 ;
      RECT  10.48 0.345 10.6 0.725 ;
      RECT  2.85 0.51 2.95 0.8 ;
      RECT  2.74 0.8 2.95 0.97 ;
      RECT  10.3 0.355 10.39 0.845 ;
      RECT  10.3 0.845 10.66 1.025 ;
      RECT  10.3 1.025 10.39 1.48 ;
      RECT  9.385 1.48 10.39 1.6 ;
      RECT  11.74 0.79 12.81 0.89 ;
      RECT  11.74 0.89 11.84 1.31 ;
      RECT  8.95 0.51 9.05 0.95 ;
      RECT  8.585 0.95 9.05 1.12 ;
      RECT  8.93 1.12 9.05 1.31 ;
      RECT  4.055 0.375 4.175 1.015 ;
      RECT  4.055 1.015 4.515 1.125 ;
      RECT  4.415 0.71 4.515 1.015 ;
      RECT  5.3 0.425 5.39 1.015 ;
      RECT  5.3 1.015 7.475 1.115 ;
      RECT  7.385 0.77 7.475 1.015 ;
      RECT  5.3 1.115 5.405 1.42 ;
      RECT  4.695 1.42 5.405 1.525 ;
      RECT  1.79 0.925 2.065 1.035 ;
      RECT  1.79 1.035 1.88 1.255 ;
      RECT  0.35 0.19 0.44 1.08 ;
      RECT  0.065 1.08 1.36 1.17 ;
      RECT  1.27 1.17 1.36 1.255 ;
      RECT  0.065 1.17 0.185 1.61 ;
      RECT  1.27 1.255 1.88 1.345 ;
      RECT  0.535 1.26 1.18 1.35 ;
      RECT  1.09 1.35 1.18 1.46 ;
      RECT  1.09 1.46 1.895 1.58 ;
      RECT  11.525 0.2 11.65 1.405 ;
      RECT  10.545 1.405 11.65 1.52 ;
      RECT  10.545 1.52 10.635 1.61 ;
      LAYER M2 ;
      RECT  0.82 0.35 2.59 0.45 ;
      RECT  2.81 0.55 10.62 0.65 ;
      RECT  4.375 0.75 5.62 0.85 ;
      RECT  8.31 1.15 11.88 1.25 ;
      LAYER V1 ;
      RECT  0.86 0.35 0.96 0.45 ;
      RECT  2.45 0.35 2.55 0.45 ;
      RECT  2.85 0.55 2.95 0.65 ;
      RECT  8.95 0.55 9.05 0.65 ;
      RECT  9.6 0.55 9.7 0.65 ;
      RECT  10.48 0.55 10.58 0.65 ;
      RECT  4.415 0.75 4.515 0.85 ;
      RECT  5.48 0.75 5.58 0.85 ;
      RECT  8.35 1.15 8.45 1.25 ;
      RECT  10.11 1.15 10.21 1.25 ;
      RECT  11.74 1.15 11.84 1.25 ;
  END
END SEN_FSDPRBSBQO_6
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPRBSBQO_8
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-clear/set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),clear=!RD,preset=!SD,clear_preset_var1=0):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPRBSBQO_8
  CLASS CORE ;
  FOREIGN SEN_FSDPRBSBQO_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.535 0.31 9.635 0.76 ;
      RECT  9.535 0.76 9.69 0.775 ;
      RECT  9.3 0.775 9.69 0.865 ;
      LAYER M2 ;
      RECT  9.495 0.35 10.49 0.45 ;
      LAYER V1 ;
      RECT  9.535 0.35 9.635 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.76 ;
      RECT  0.55 0.76 1.235 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  12.255 0.51 13.965 0.69 ;
      RECT  13.48 0.69 13.65 1.11 ;
      RECT  12.15 1.11 13.975 1.29 ;
    END
    ANTENNADIFFAREA 0.88 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.79 0.75 10.2 0.85 ;
      RECT  10.095 0.85 10.195 0.94 ;
      RECT  9.79 0.85 9.89 1.0 ;
      RECT  9.335 1.0 9.89 1.11 ;
      RECT  6.185 0.745 7.11 0.855 ;
      LAYER M2 ;
      RECT  6.73 0.75 10.2 0.85 ;
      LAYER V1 ;
      RECT  10.06 0.75 10.16 0.85 ;
      RECT  6.77 0.75 6.87 0.85 ;
      RECT  6.97 0.75 7.07 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.18 ;
  END RD
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.35 0.78 11.45 1.2 ;
      RECT  4.605 0.91 4.93 1.09 ;
      LAYER M2 ;
      RECT  4.79 0.95 11.49 1.05 ;
      LAYER V1 ;
      RECT  11.35 0.95 11.45 1.05 ;
      RECT  4.83 0.95 4.93 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.26 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1188 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.65 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0474 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  11.0 0.22 11.105 0.51 ;
      RECT  11.0 0.51 11.45 0.69 ;
      RECT  11.15 0.69 11.25 1.12 ;
      RECT  10.835 1.12 11.25 1.24 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  9.175 1.2 9.825 1.29 ;
      RECT  9.705 1.29 9.825 1.37 ;
      RECT  9.175 1.29 9.295 1.75 ;
      RECT  0.325 1.4 0.445 1.75 ;
      RECT  0.0 1.75 14.4 1.85 ;
      RECT  0.845 1.415 0.965 1.75 ;
      RECT  2.5 1.48 2.67 1.75 ;
      RECT  4.485 1.39 4.605 1.75 ;
      RECT  4.99 1.61 5.16 1.75 ;
      RECT  5.545 1.2 5.665 1.75 ;
      RECT  6.065 1.44 6.185 1.75 ;
      RECT  6.585 1.44 6.705 1.75 ;
      RECT  7.105 1.44 7.225 1.75 ;
      RECT  8.655 1.29 8.775 1.75 ;
      RECT  11.13 1.6 11.3 1.75 ;
      RECT  11.935 1.185 12.055 1.75 ;
      RECT  12.47 1.4 12.59 1.75 ;
      RECT  13.02 1.39 13.14 1.75 ;
      RECT  13.57 1.39 13.69 1.75 ;
      RECT  14.13 1.21 14.25 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 14.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 14.4 0.05 ;
      RECT  9.415 0.05 9.585 0.185 ;
      RECT  5.94 0.05 6.11 0.215 ;
      RECT  6.48 0.05 6.65 0.215 ;
      RECT  7.02 0.05 7.19 0.215 ;
      RECT  1.75 0.05 1.855 0.36 ;
      RECT  4.565 0.05 4.685 0.36 ;
      RECT  2.765 0.05 2.885 0.385 ;
      RECT  11.245 0.05 11.365 0.385 ;
      RECT  0.065 0.05 0.205 0.39 ;
      RECT  12.515 0.05 12.635 0.42 ;
      RECT  13.035 0.05 13.155 0.42 ;
      RECT  13.56 0.05 13.68 0.42 ;
      RECT  9.975 0.05 10.095 0.45 ;
      RECT  2.255 0.05 2.36 0.585 ;
      RECT  11.965 0.05 12.085 0.585 ;
      RECT  14.13 0.05 14.25 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 14.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.865 0.14 5.565 0.23 ;
      RECT  5.445 0.23 5.565 0.385 ;
      RECT  4.865 0.23 4.985 0.45 ;
      RECT  4.28 0.45 4.985 0.57 ;
      RECT  10.29 0.14 10.9 0.245 ;
      RECT  10.29 0.245 10.38 1.06 ;
      RECT  10.25 1.06 10.38 1.135 ;
      RECT  10.25 1.135 10.35 1.235 ;
      RECT  10.095 1.235 10.35 1.355 ;
      RECT  3.04 0.14 4.13 0.25 ;
      RECT  3.04 0.25 3.145 1.08 ;
      RECT  2.745 1.08 3.44 1.19 ;
      RECT  7.315 0.22 8.525 0.33 ;
      RECT  5.655 0.33 8.525 0.34 ;
      RECT  5.655 0.34 7.435 0.45 ;
      RECT  0.545 0.215 0.9 0.335 ;
      RECT  0.72 0.335 0.9 0.45 ;
      RECT  1.065 0.215 1.66 0.335 ;
      RECT  1.57 0.335 1.66 0.475 ;
      RECT  1.57 0.475 2.165 0.595 ;
      RECT  11.56 0.215 11.86 0.335 ;
      RECT  11.56 0.335 11.65 1.38 ;
      RECT  10.62 1.38 11.65 1.495 ;
      RECT  10.62 1.495 10.71 1.58 ;
      RECT  8.615 0.245 9.345 0.365 ;
      RECT  8.615 0.365 8.735 0.475 ;
      RECT  7.935 0.475 8.735 0.565 ;
      RECT  5.38 0.565 8.735 0.595 ;
      RECT  5.38 0.595 8.03 0.655 ;
      RECT  5.38 0.655 5.48 0.89 ;
      RECT  7.94 0.655 8.03 0.99 ;
      RECT  7.38 0.99 8.03 1.08 ;
      RECT  7.38 1.08 7.485 1.245 ;
      RECT  5.755 1.245 7.485 1.35 ;
      RECT  7.365 1.35 7.485 1.47 ;
      RECT  7.365 1.47 8.565 1.585 ;
      RECT  2.45 0.235 2.625 0.415 ;
      RECT  2.45 0.415 2.55 0.59 ;
      RECT  3.235 0.34 3.915 0.46 ;
      RECT  3.81 0.46 3.915 1.21 ;
      RECT  3.81 1.21 5.11 1.3 ;
      RECT  5.02 0.785 5.11 1.21 ;
      RECT  3.985 1.3 4.105 1.495 ;
      RECT  3.255 1.495 4.105 1.6 ;
      RECT  9.725 0.25 9.815 0.55 ;
      RECT  9.725 0.55 9.905 0.655 ;
      RECT  3.485 0.55 3.71 0.67 ;
      RECT  3.62 0.67 3.71 1.3 ;
      RECT  1.375 0.455 1.48 0.54 ;
      RECT  0.805 0.54 1.48 0.64 ;
      RECT  1.375 0.64 1.48 0.71 ;
      RECT  1.375 0.71 2.25 0.795 ;
      RECT  1.45 0.795 2.25 0.8 ;
      RECT  1.45 0.8 1.555 1.17 ;
      RECT  2.16 0.8 2.25 1.22 ;
      RECT  2.01 1.22 2.25 1.3 ;
      RECT  2.01 1.3 3.71 1.39 ;
      RECT  3.06 1.39 3.71 1.405 ;
      RECT  3.06 1.405 3.15 1.53 ;
      RECT  10.65 0.51 10.91 0.705 ;
      RECT  8.915 0.475 9.02 0.71 ;
      RECT  8.125 0.71 9.02 0.8 ;
      RECT  8.125 0.8 8.225 1.24 ;
      RECT  7.625 1.17 7.745 1.24 ;
      RECT  7.625 1.24 8.315 1.345 ;
      RECT  10.47 0.36 10.56 0.825 ;
      RECT  10.47 0.825 11.06 0.92 ;
      RECT  10.47 0.92 10.56 1.21 ;
      RECT  10.44 1.21 10.56 1.285 ;
      RECT  10.44 1.285 10.53 1.47 ;
      RECT  9.385 1.47 10.53 1.585 ;
      RECT  2.85 0.49 2.95 0.83 ;
      RECT  2.76 0.83 2.95 0.94 ;
      RECT  11.74 0.785 13.38 0.895 ;
      RECT  11.74 0.895 11.84 1.31 ;
      RECT  7.2 0.79 7.85 0.9 ;
      RECT  7.2 0.9 7.29 1.01 ;
      RECT  5.2 0.32 5.29 1.01 ;
      RECT  5.2 1.01 7.29 1.11 ;
      RECT  5.2 1.11 5.395 1.115 ;
      RECT  5.295 1.115 5.395 1.4 ;
      RECT  4.72 1.4 5.395 1.52 ;
      RECT  9.11 0.51 9.21 0.995 ;
      RECT  8.315 0.995 9.21 1.095 ;
      RECT  8.915 1.095 9.035 1.53 ;
      RECT  4.055 0.34 4.175 1.02 ;
      RECT  4.055 1.02 4.515 1.12 ;
      RECT  4.415 0.69 4.515 1.02 ;
      RECT  1.83 0.92 2.07 1.03 ;
      RECT  1.83 1.03 1.92 1.26 ;
      RECT  0.35 0.19 0.455 0.99 ;
      RECT  0.35 0.99 1.36 1.08 ;
      RECT  0.35 1.08 0.44 1.22 ;
      RECT  1.27 1.08 1.36 1.26 ;
      RECT  0.065 1.22 0.44 1.31 ;
      RECT  1.27 1.26 1.92 1.35 ;
      RECT  0.065 1.31 0.185 1.61 ;
      RECT  0.535 1.2 1.18 1.32 ;
      RECT  1.09 1.32 1.18 1.465 ;
      RECT  1.09 1.465 1.865 1.585 ;
      LAYER M2 ;
      RECT  0.72 0.35 2.59 0.45 ;
      RECT  2.81 0.55 10.79 0.65 ;
      RECT  4.375 0.75 5.52 0.85 ;
      RECT  8.085 1.15 11.88 1.25 ;
      LAYER V1 ;
      RECT  0.76 0.35 0.86 0.45 ;
      RECT  2.45 0.35 2.55 0.45 ;
      RECT  2.85 0.55 2.95 0.65 ;
      RECT  9.11 0.55 9.21 0.65 ;
      RECT  9.765 0.55 9.865 0.65 ;
      RECT  10.65 0.55 10.75 0.65 ;
      RECT  4.415 0.75 4.515 0.85 ;
      RECT  5.38 0.75 5.48 0.85 ;
      RECT  8.125 1.15 8.225 1.25 ;
      RECT  10.25 1.15 10.35 1.25 ;
      RECT  11.74 1.15 11.84 1.25 ;
  END
END SEN_FSDPRBSBQO_8
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPSBQ_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPSBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDPSBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.94 0.71 2.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.84 0.83 0.93 ;
      RECT  0.35 0.93 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 5.95 0.69 ;
      RECT  5.86 0.69 5.95 1.11 ;
      RECT  5.75 1.11 5.95 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.92 0.87 5.06 1.23 ;
      RECT  3.385 0.905 3.84 1.055 ;
      LAYER M2 ;
      RECT  3.44 0.95 5.085 1.05 ;
      LAYER V1 ;
      RECT  4.945 0.95 5.045 1.05 ;
      RECT  3.485 0.95 3.585 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.49 ;
      RECT  0.35 0.49 1.265 0.51 ;
      RECT  0.15 0.51 1.265 0.59 ;
      RECT  0.15 0.59 0.555 0.69 ;
      RECT  1.15 0.59 1.265 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.88 0.25 1.5 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.61 0.225 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  1.315 1.605 1.485 1.75 ;
      RECT  1.95 1.6 2.12 1.75 ;
      RECT  3.26 1.505 3.43 1.75 ;
      RECT  3.665 1.5 3.835 1.75 ;
      RECT  4.795 1.52 4.965 1.75 ;
      RECT  5.565 0.99 5.66 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  1.065 0.05 1.235 0.19 ;
      RECT  1.945 0.05 2.115 0.19 ;
      RECT  3.215 0.05 3.425 0.32 ;
      RECT  5.01 0.05 5.18 0.325 ;
      RECT  0.075 0.05 0.205 0.39 ;
      RECT  5.555 0.05 5.66 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.575 0.18 0.705 0.295 ;
      RECT  0.575 0.295 2.66 0.385 ;
      RECT  2.535 0.18 2.66 0.295 ;
      RECT  2.77 0.215 2.95 0.335 ;
      RECT  2.845 0.335 2.95 0.66 ;
      RECT  2.845 0.66 3.87 0.765 ;
      RECT  2.845 0.765 2.95 1.24 ;
      RECT  2.765 1.24 2.95 1.36 ;
      RECT  4.26 0.215 4.46 0.335 ;
      RECT  4.37 0.335 4.46 0.67 ;
      RECT  4.37 0.67 5.27 0.76 ;
      RECT  5.17 0.76 5.27 0.94 ;
      RECT  4.69 0.76 4.78 1.14 ;
      RECT  4.26 1.14 4.78 1.23 ;
      RECT  4.26 1.23 4.38 1.6 ;
      RECT  4.655 0.4 4.825 0.44 ;
      RECT  4.655 0.44 5.45 0.57 ;
      RECT  5.295 0.26 5.45 0.44 ;
      RECT  5.36 0.57 5.45 0.8 ;
      RECT  5.36 0.8 5.77 0.9 ;
      RECT  5.36 0.9 5.45 1.05 ;
      RECT  5.29 1.05 5.45 1.165 ;
      RECT  5.29 1.165 5.405 1.325 ;
      RECT  3.75 0.38 4.055 0.5 ;
      RECT  3.96 0.5 4.055 1.17 ;
      RECT  3.145 0.87 3.255 1.17 ;
      RECT  3.145 1.17 4.055 1.24 ;
      RECT  3.145 1.24 4.125 1.275 ;
      RECT  3.96 1.275 4.125 1.415 ;
      RECT  2.275 0.48 2.4 0.55 ;
      RECT  2.275 0.55 2.755 0.65 ;
      RECT  2.275 0.65 2.4 0.83 ;
      RECT  2.275 0.83 2.7 0.94 ;
      RECT  2.275 0.94 2.395 1.22 ;
      RECT  1.67 0.49 1.82 0.67 ;
      RECT  1.73 0.67 1.82 1.38 ;
      RECT  1.705 1.38 1.82 1.4 ;
      RECT  1.705 1.4 2.33 1.49 ;
      RECT  2.24 1.49 2.33 1.57 ;
      RECT  1.705 1.49 1.825 1.61 ;
      RECT  2.24 1.57 3.1 1.66 ;
      RECT  4.145 0.44 4.25 0.87 ;
      RECT  4.145 0.87 4.59 1.03 ;
      RECT  1.375 0.5 1.47 0.99 ;
      RECT  1.375 0.99 1.64 1.16 ;
      RECT  1.375 1.16 1.48 1.2 ;
      RECT  0.93 0.7 1.02 1.2 ;
      RECT  0.93 1.2 1.48 1.3 ;
      RECT  0.93 1.3 1.02 1.57 ;
      RECT  0.37 1.57 1.02 1.66 ;
      RECT  0.58 1.2 0.7 1.335 ;
      RECT  0.58 1.335 0.84 1.46 ;
      RECT  2.53 1.11 2.65 1.35 ;
      RECT  2.45 1.35 2.65 1.45 ;
      RECT  4.52 1.34 5.2 1.43 ;
      RECT  4.52 1.43 4.64 1.62 ;
      RECT  5.095 1.43 5.2 1.62 ;
      LAYER M2 ;
      RECT  2.575 0.55 4.29 0.65 ;
      RECT  0.66 1.35 2.635 1.45 ;
      LAYER V1 ;
      RECT  2.615 0.55 2.715 0.65 ;
      RECT  4.15 0.55 4.25 0.65 ;
      RECT  0.7 1.35 0.8 1.45 ;
      RECT  2.49 1.35 2.59 1.45 ;
  END
END SEN_FSDPSBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPSBQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPSBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPSBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.94 0.71 2.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.84 0.83 0.93 ;
      RECT  0.35 0.93 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.895 0.51 6.25 0.69 ;
      RECT  6.15 0.69 6.25 1.015 ;
      RECT  5.895 1.015 6.25 1.115 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.92 0.87 5.06 1.23 ;
      RECT  3.385 0.905 3.84 1.055 ;
      LAYER M2 ;
      RECT  3.44 0.95 5.085 1.05 ;
      LAYER V1 ;
      RECT  4.945 0.95 5.045 1.05 ;
      RECT  3.485 0.95 3.585 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.49 ;
      RECT  0.35 0.49 1.265 0.51 ;
      RECT  0.15 0.51 1.265 0.59 ;
      RECT  0.15 0.59 0.555 0.69 ;
      RECT  1.15 0.59 1.265 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.88 0.25 1.5 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.61 0.225 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  1.315 1.605 1.485 1.75 ;
      RECT  1.95 1.6 2.12 1.75 ;
      RECT  3.26 1.505 3.43 1.75 ;
      RECT  3.665 1.5 3.835 1.75 ;
      RECT  4.795 1.52 4.965 1.75 ;
      RECT  5.63 1.21 5.75 1.75 ;
      RECT  6.2 1.21 6.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  1.065 0.05 1.235 0.19 ;
      RECT  1.945 0.05 2.115 0.19 ;
      RECT  3.215 0.05 3.425 0.32 ;
      RECT  5.05 0.05 5.26 0.345 ;
      RECT  0.075 0.05 0.205 0.39 ;
      RECT  6.195 0.05 6.325 0.39 ;
      RECT  5.65 0.05 5.77 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.575 0.18 0.705 0.295 ;
      RECT  0.575 0.295 2.66 0.385 ;
      RECT  2.535 0.17 2.66 0.295 ;
      RECT  2.77 0.215 2.95 0.335 ;
      RECT  2.845 0.335 2.95 0.66 ;
      RECT  2.845 0.66 3.87 0.765 ;
      RECT  2.845 0.765 2.95 1.24 ;
      RECT  2.765 1.24 2.95 1.36 ;
      RECT  4.26 0.215 4.46 0.335 ;
      RECT  4.37 0.335 4.46 0.67 ;
      RECT  4.37 0.67 5.325 0.76 ;
      RECT  5.225 0.76 5.325 0.96 ;
      RECT  4.69 0.76 4.78 1.14 ;
      RECT  4.26 1.14 4.78 1.23 ;
      RECT  4.26 1.23 4.38 1.6 ;
      RECT  4.655 0.4 4.825 0.44 ;
      RECT  4.655 0.44 5.505 0.57 ;
      RECT  5.415 0.57 5.505 0.795 ;
      RECT  5.415 0.795 6.06 0.895 ;
      RECT  5.415 0.895 5.505 1.175 ;
      RECT  5.29 1.175 5.505 1.29 ;
      RECT  3.75 0.38 4.055 0.5 ;
      RECT  3.96 0.5 4.055 1.17 ;
      RECT  3.145 0.87 3.255 1.17 ;
      RECT  3.145 1.17 4.055 1.24 ;
      RECT  3.145 1.24 4.125 1.275 ;
      RECT  3.96 1.275 4.125 1.415 ;
      RECT  2.275 0.48 2.4 0.55 ;
      RECT  2.275 0.55 2.755 0.65 ;
      RECT  2.275 0.65 2.4 0.83 ;
      RECT  2.275 0.83 2.7 0.94 ;
      RECT  2.275 0.94 2.395 1.22 ;
      RECT  1.67 0.49 1.82 0.67 ;
      RECT  1.73 0.67 1.82 1.38 ;
      RECT  1.705 1.38 1.82 1.4 ;
      RECT  1.705 1.4 2.33 1.49 ;
      RECT  2.24 1.49 2.33 1.57 ;
      RECT  1.705 1.49 1.825 1.61 ;
      RECT  2.24 1.57 3.1 1.66 ;
      RECT  4.145 0.44 4.25 0.87 ;
      RECT  4.145 0.87 4.59 1.03 ;
      RECT  1.375 0.5 1.47 0.99 ;
      RECT  1.375 0.99 1.64 1.16 ;
      RECT  1.375 1.16 1.48 1.2 ;
      RECT  0.93 0.7 1.02 1.2 ;
      RECT  0.93 1.2 1.48 1.3 ;
      RECT  0.93 1.3 1.02 1.57 ;
      RECT  0.37 1.57 1.02 1.66 ;
      RECT  0.58 1.2 0.7 1.335 ;
      RECT  0.58 1.335 0.84 1.46 ;
      RECT  2.53 1.11 2.65 1.35 ;
      RECT  2.45 1.35 2.65 1.45 ;
      RECT  4.52 1.34 5.2 1.43 ;
      RECT  4.52 1.43 4.64 1.62 ;
      RECT  5.095 1.43 5.2 1.62 ;
      LAYER M2 ;
      RECT  2.575 0.55 4.29 0.65 ;
      RECT  0.66 1.35 2.635 1.45 ;
      LAYER V1 ;
      RECT  2.615 0.55 2.715 0.65 ;
      RECT  4.15 0.55 4.25 0.65 ;
      RECT  0.7 1.35 0.8 1.45 ;
      RECT  2.49 1.35 2.59 1.45 ;
  END
END SEN_FSDPSBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPSBQ_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-/set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPSBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDPSBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.94 0.71 2.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0528 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.84 0.83 0.93 ;
      RECT  0.35 0.93 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.31 6.46 0.51 ;
      RECT  5.75 0.51 6.46 0.69 ;
      RECT  6.35 0.69 6.46 1.015 ;
      RECT  5.8 1.015 6.46 1.115 ;
      RECT  6.35 1.115 6.46 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.92 0.87 5.06 1.23 ;
      RECT  3.385 0.905 3.84 1.055 ;
      LAYER M2 ;
      RECT  3.44 0.95 5.085 1.05 ;
      LAYER V1 ;
      RECT  4.945 0.95 5.045 1.05 ;
      RECT  3.485 0.95 3.585 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.49 ;
      RECT  0.35 0.49 1.265 0.51 ;
      RECT  0.15 0.51 1.265 0.59 ;
      RECT  0.15 0.59 0.555 0.69 ;
      RECT  1.15 0.59 1.265 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.88 0.25 1.5 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.018 ;
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.61 0.225 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.315 1.605 1.485 1.75 ;
      RECT  1.95 1.6 2.12 1.75 ;
      RECT  3.26 1.505 3.43 1.75 ;
      RECT  3.665 1.5 3.835 1.75 ;
      RECT  4.795 1.52 4.965 1.75 ;
      RECT  5.58 1.215 5.695 1.75 ;
      RECT  6.095 1.21 6.215 1.75 ;
      RECT  6.615 1.21 6.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  1.065 0.05 1.235 0.19 ;
      RECT  1.945 0.05 2.115 0.19 ;
      RECT  3.235 0.05 3.445 0.32 ;
      RECT  5.05 0.05 5.26 0.345 ;
      RECT  5.57 0.05 5.7 0.365 ;
      RECT  0.075 0.05 0.205 0.39 ;
      RECT  6.09 0.05 6.22 0.4 ;
      RECT  6.615 0.05 6.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.575 0.18 0.705 0.295 ;
      RECT  0.575 0.295 2.66 0.385 ;
      RECT  2.535 0.17 2.66 0.295 ;
      RECT  2.77 0.215 2.95 0.335 ;
      RECT  2.845 0.335 2.95 0.66 ;
      RECT  2.845 0.66 3.87 0.765 ;
      RECT  2.845 0.765 2.95 1.24 ;
      RECT  2.765 1.24 2.95 1.36 ;
      RECT  4.26 0.215 4.46 0.335 ;
      RECT  4.37 0.335 4.46 0.67 ;
      RECT  4.37 0.67 5.325 0.76 ;
      RECT  5.225 0.76 5.325 0.95 ;
      RECT  4.69 0.76 4.78 1.14 ;
      RECT  4.26 1.14 4.78 1.23 ;
      RECT  4.26 1.23 4.38 1.6 ;
      RECT  4.655 0.4 4.825 0.44 ;
      RECT  4.655 0.44 5.505 0.57 ;
      RECT  5.415 0.57 5.505 0.795 ;
      RECT  5.415 0.795 6.25 0.895 ;
      RECT  5.415 0.895 5.505 1.05 ;
      RECT  5.27 1.05 5.505 1.165 ;
      RECT  3.75 0.38 4.055 0.5 ;
      RECT  3.96 0.5 4.055 1.17 ;
      RECT  3.145 0.87 3.255 1.17 ;
      RECT  3.145 1.17 4.055 1.24 ;
      RECT  3.145 1.24 4.125 1.275 ;
      RECT  3.96 1.275 4.125 1.415 ;
      RECT  2.275 0.48 2.4 0.55 ;
      RECT  2.275 0.55 2.755 0.65 ;
      RECT  2.275 0.65 2.4 0.83 ;
      RECT  2.275 0.83 2.7 0.94 ;
      RECT  2.275 0.94 2.395 1.22 ;
      RECT  1.67 0.49 1.82 0.67 ;
      RECT  1.73 0.67 1.82 1.38 ;
      RECT  1.705 1.38 1.82 1.4 ;
      RECT  1.705 1.4 2.33 1.49 ;
      RECT  2.24 1.49 2.33 1.57 ;
      RECT  1.705 1.49 1.825 1.61 ;
      RECT  2.24 1.57 3.1 1.66 ;
      RECT  4.145 0.44 4.25 0.87 ;
      RECT  4.145 0.87 4.59 1.03 ;
      RECT  1.375 0.5 1.47 0.99 ;
      RECT  1.375 0.99 1.64 1.16 ;
      RECT  1.375 1.16 1.48 1.2 ;
      RECT  0.93 0.7 1.02 1.2 ;
      RECT  0.93 1.2 1.48 1.3 ;
      RECT  0.93 1.3 1.02 1.57 ;
      RECT  0.37 1.57 1.02 1.66 ;
      RECT  0.58 1.2 0.7 1.335 ;
      RECT  0.58 1.335 0.84 1.46 ;
      RECT  2.53 1.11 2.65 1.35 ;
      RECT  2.45 1.35 2.65 1.45 ;
      RECT  4.52 1.34 5.2 1.43 ;
      RECT  4.52 1.43 4.64 1.62 ;
      RECT  5.095 1.43 5.2 1.62 ;
      LAYER M2 ;
      RECT  2.575 0.55 4.29 0.65 ;
      RECT  0.66 1.35 2.635 1.45 ;
      LAYER V1 ;
      RECT  2.615 0.55 2.715 0.65 ;
      RECT  4.15 0.55 4.25 0.65 ;
      RECT  0.7 1.35 0.8 1.45 ;
      RECT  2.49 1.35 2.59 1.45 ;
  END
END SEN_FSDPSBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPSBQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPSBQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDPSBQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.51 0.71 4.65 0.9 ;
      RECT  4.55 0.9 4.65 1.25 ;
      RECT  4.55 1.25 4.935 1.34 ;
      RECT  4.845 1.34 4.935 1.43 ;
      RECT  4.845 1.43 5.17 1.53 ;
      RECT  3.27 0.69 3.37 0.925 ;
      RECT  3.27 0.925 4.0 1.025 ;
      LAYER M2 ;
      RECT  3.23 0.75 4.65 0.85 ;
      LAYER V1 ;
      RECT  4.51 0.75 4.61 0.85 ;
      RECT  3.27 0.75 3.37 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0744 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.485 1.08 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0639 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.625 0.165 6.745 0.45 ;
      RECT  6.385 0.45 6.745 0.54 ;
      RECT  6.385 0.54 6.475 0.91 ;
      RECT  6.35 0.91 6.475 1.11 ;
      RECT  6.35 1.11 6.74 1.29 ;
      RECT  6.635 1.29 6.74 1.61 ;
    END
    ANTENNADIFFAREA 0.139 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.13 0.27 6.25 0.45 ;
      RECT  6.13 0.45 6.295 0.55 ;
      RECT  6.195 0.55 6.295 0.69 ;
      RECT  1.97 0.49 2.07 0.71 ;
      RECT  1.75 0.71 2.07 0.89 ;
      LAYER M2 ;
      RECT  1.93 0.55 6.335 0.65 ;
      LAYER V1 ;
      RECT  6.195 0.55 6.295 0.65 ;
      RECT  1.97 0.55 2.07 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0597 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.295 0.71 0.475 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.395 0.505 0.85 0.605 ;
      RECT  0.735 0.605 0.85 1.03 ;
      RECT  0.735 1.03 0.87 1.12 ;
      RECT  0.78 1.12 0.87 1.365 ;
      RECT  0.78 1.365 1.58 1.455 ;
      RECT  1.38 1.455 1.58 1.495 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.645 0.51 5.735 1.11 ;
      RECT  5.55 1.11 5.735 1.31 ;
      RECT  5.55 1.31 5.65 1.49 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.49 0.505 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  1.59 1.63 1.76 1.75 ;
      RECT  2.16 1.63 2.33 1.75 ;
      RECT  3.24 1.525 3.41 1.75 ;
      RECT  4.08 1.385 4.2 1.75 ;
      RECT  5.325 1.57 5.495 1.75 ;
      RECT  5.845 1.44 5.965 1.75 ;
      RECT  6.365 1.4 6.485 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  4.07 0.05 4.24 0.195 ;
      RECT  5.32 0.05 5.49 0.24 ;
      RECT  3.245 0.05 3.415 0.335 ;
      RECT  6.365 0.05 6.485 0.36 ;
      RECT  1.55 0.05 1.68 0.385 ;
      RECT  0.325 0.05 0.445 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.77 0.18 2.5 0.27 ;
      RECT  2.385 0.27 2.5 0.465 ;
      RECT  1.77 0.27 1.86 0.475 ;
      RECT  0.835 0.215 1.395 0.325 ;
      RECT  1.305 0.325 1.395 0.475 ;
      RECT  1.305 0.475 1.86 0.565 ;
      RECT  1.305 0.565 1.395 1.105 ;
      RECT  0.96 1.105 1.395 1.185 ;
      RECT  0.96 1.185 1.825 1.275 ;
      RECT  1.735 1.275 1.825 1.43 ;
      RECT  1.735 1.43 2.6 1.54 ;
      RECT  4.375 0.175 5.11 0.275 ;
      RECT  4.375 0.275 4.465 0.31 ;
      RECT  4.11 0.31 4.465 0.4 ;
      RECT  4.11 0.4 4.2 0.705 ;
      RECT  3.46 0.63 3.55 0.705 ;
      RECT  3.46 0.705 4.2 0.8 ;
      RECT  3.815 0.495 3.93 0.705 ;
      RECT  4.11 0.8 4.2 1.16 ;
      RECT  3.785 1.16 4.2 1.255 ;
      RECT  5.83 0.225 5.96 0.33 ;
      RECT  5.205 0.33 5.96 0.395 ;
      RECT  5.205 0.395 5.915 0.42 ;
      RECT  5.205 0.42 5.305 0.815 ;
      RECT  5.825 0.42 5.915 1.26 ;
      RECT  5.825 1.26 6.225 1.35 ;
      RECT  6.105 1.35 6.225 1.615 ;
      RECT  3.55 0.19 3.67 0.45 ;
      RECT  2.895 0.45 3.67 0.54 ;
      RECT  2.895 0.54 2.985 0.72 ;
      RECT  2.86 0.72 2.985 0.89 ;
      RECT  2.895 0.89 2.985 1.165 ;
      RECT  2.895 1.165 3.695 1.255 ;
      RECT  4.65 0.41 4.935 0.525 ;
      RECT  4.795 0.525 4.935 1.16 ;
      RECT  2.16 0.41 2.255 0.605 ;
      RECT  2.16 0.605 2.25 1.25 ;
      RECT  1.915 1.145 2.02 1.25 ;
      RECT  1.915 1.25 2.78 1.34 ;
      RECT  2.69 1.34 2.78 1.345 ;
      RECT  2.69 1.345 3.85 1.435 ;
      RECT  3.06 1.435 3.15 1.59 ;
      RECT  3.74 1.435 3.85 1.66 ;
      RECT  4.33 0.5 4.55 0.62 ;
      RECT  4.33 0.62 4.42 1.025 ;
      RECT  4.33 1.025 4.445 1.115 ;
      RECT  4.355 1.115 4.445 1.46 ;
      RECT  4.355 1.46 4.74 1.575 ;
      RECT  5.025 0.38 5.115 0.905 ;
      RECT  5.025 0.905 5.555 0.995 ;
      RECT  5.46 0.76 5.555 0.905 ;
      RECT  5.025 0.995 5.115 1.165 ;
      RECT  5.025 1.165 5.27 1.28 ;
      RECT  2.34 0.835 2.435 0.945 ;
      RECT  2.34 0.945 2.745 0.99 ;
      RECT  2.655 0.245 2.745 0.945 ;
      RECT  2.34 0.99 2.805 1.035 ;
      RECT  2.665 1.035 2.805 1.16 ;
      RECT  6.565 0.635 6.745 0.965 ;
      RECT  6.005 0.71 6.105 0.975 ;
      RECT  6.005 0.975 6.24 1.08 ;
      RECT  0.065 0.18 0.185 1.31 ;
      RECT  0.065 1.31 0.69 1.4 ;
      RECT  0.6 1.4 0.69 1.545 ;
      RECT  0.065 1.4 0.185 1.61 ;
      RECT  0.6 1.545 1.305 1.66 ;
      LAYER M2 ;
      RECT  4.795 0.75 6.73 0.85 ;
      LAYER V1 ;
      RECT  4.835 0.75 4.935 0.85 ;
      RECT  6.005 0.75 6.105 0.85 ;
      RECT  6.59 0.75 6.69 0.85 ;
  END
END SEN_FSDPSBQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPSBQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPSBQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDPSBQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.48 7.11 0.92 ;
      RECT  6.255 0.605 6.435 0.89 ;
      RECT  5.08 0.74 5.715 0.855 ;
      LAYER M2 ;
      RECT  5.535 0.75 7.15 0.85 ;
      LAYER V1 ;
      RECT  7.01 0.75 7.11 0.85 ;
      RECT  6.335 0.75 6.435 0.85 ;
      RECT  5.575 0.75 5.675 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0981 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.435 0.7 2.45 0.79 ;
      RECT  2.35 0.79 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0834 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.97 0.19 9.075 0.45 ;
      RECT  8.97 0.45 9.25 0.54 ;
      RECT  9.15 0.54 9.25 1.105 ;
      RECT  8.98 1.105 9.25 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.53 0.665 8.685 0.91 ;
      RECT  8.585 0.91 8.685 1.115 ;
      RECT  4.605 0.775 4.79 1.09 ;
      LAYER M2 ;
      RECT  4.565 0.95 8.725 1.05 ;
      LAYER V1 ;
      RECT  8.585 0.95 8.685 1.05 ;
      RECT  4.605 0.95 4.705 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.069 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.665 0.45 1.265 ;
      RECT  0.35 1.265 1.585 1.355 ;
      RECT  1.415 1.225 1.585 1.265 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.087 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.505 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.84 0.31 8.05 0.485 ;
      RECT  7.95 0.485 8.05 1.015 ;
      RECT  7.775 1.015 8.05 1.12 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.63 0.5 1.75 ;
      RECT  0.0 1.75 9.4 1.85 ;
      RECT  1.415 1.445 1.585 1.75 ;
      RECT  2.445 1.48 2.615 1.75 ;
      RECT  3.95 1.405 4.07 1.75 ;
      RECT  4.52 1.4 4.64 1.75 ;
      RECT  5.08 1.215 5.2 1.75 ;
      RECT  5.865 1.6 6.035 1.75 ;
      RECT  7.515 1.63 7.685 1.75 ;
      RECT  8.08 1.63 8.25 1.75 ;
      RECT  8.72 1.455 8.825 1.75 ;
      RECT  9.215 1.41 9.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      RECT  1.905 0.05 2.075 0.195 ;
      RECT  5.865 0.05 6.035 0.195 ;
      RECT  8.645 0.05 8.815 0.32 ;
      RECT  9.225 0.05 9.345 0.36 ;
      RECT  0.065 0.05 0.2 0.385 ;
      RECT  5.375 0.05 5.495 0.385 ;
      RECT  3.97 0.05 4.09 0.39 ;
      RECT  2.68 0.05 2.81 0.395 ;
      RECT  7.535 0.05 7.675 0.42 ;
      RECT  4.775 0.05 4.925 0.435 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.63 0.14 1.54 0.23 ;
      RECT  0.63 0.23 0.72 0.91 ;
      RECT  0.63 0.91 2.25 1.0 ;
      RECT  0.885 1.0 1.055 1.175 ;
      RECT  2.16 1.0 2.25 1.265 ;
      RECT  2.16 1.265 3.305 1.39 ;
      RECT  3.185 0.23 3.305 1.265 ;
      RECT  2.16 1.39 2.25 1.43 ;
      RECT  1.915 1.43 2.25 1.53 ;
      RECT  5.62 0.26 5.715 0.365 ;
      RECT  5.62 0.365 6.32 0.395 ;
      RECT  5.62 0.395 6.615 0.455 ;
      RECT  6.19 0.455 6.615 0.5 ;
      RECT  6.525 0.5 6.615 1.27 ;
      RECT  6.525 1.27 6.84 1.275 ;
      RECT  6.19 1.275 6.84 1.365 ;
      RECT  6.67 1.365 6.84 1.405 ;
      RECT  6.19 1.365 6.28 1.41 ;
      RECT  5.555 1.41 6.28 1.51 ;
      RECT  0.85 0.325 2.59 0.415 ;
      RECT  0.37 0.2 0.46 0.475 ;
      RECT  0.12 0.475 0.46 0.565 ;
      RECT  0.12 0.565 0.22 1.29 ;
      RECT  8.32 0.42 8.88 0.51 ;
      RECT  8.32 0.51 8.41 0.765 ;
      RECT  8.775 0.51 8.88 0.785 ;
      RECT  8.775 0.785 9.035 0.895 ;
      RECT  8.775 0.895 8.865 1.27 ;
      RECT  8.535 1.27 8.865 1.365 ;
      RECT  8.535 1.365 8.63 1.45 ;
      RECT  6.39 0.175 6.81 0.26 ;
      RECT  6.39 0.26 7.11 0.305 ;
      RECT  6.72 0.305 7.11 0.38 ;
      RECT  6.72 0.38 6.81 1.01 ;
      RECT  6.72 1.01 7.07 1.18 ;
      RECT  6.97 1.18 7.07 1.45 ;
      RECT  6.97 1.45 8.63 1.515 ;
      RECT  6.41 1.475 6.58 1.515 ;
      RECT  6.41 1.515 8.63 1.54 ;
      RECT  6.41 1.54 7.1 1.62 ;
      RECT  5.065 0.245 5.17 0.545 ;
      RECT  5.065 0.545 6.075 0.635 ;
      RECT  5.985 0.635 6.075 1.085 ;
      RECT  5.985 1.085 6.435 1.15 ;
      RECT  6.345 1.005 6.435 1.085 ;
      RECT  5.35 1.15 6.435 1.175 ;
      RECT  5.35 1.175 6.075 1.25 ;
      RECT  5.35 1.25 5.45 1.47 ;
      RECT  1.055 0.505 2.37 0.595 ;
      RECT  3.81 0.525 4.97 0.615 ;
      RECT  3.81 0.615 4.39 0.62 ;
      RECT  4.88 0.615 4.97 0.95 ;
      RECT  3.81 0.62 3.9 0.755 ;
      RECT  4.3 0.62 4.39 1.21 ;
      RECT  4.88 0.95 5.895 1.05 ;
      RECT  5.805 0.77 5.895 0.95 ;
      RECT  4.88 1.05 4.97 1.455 ;
      RECT  4.185 1.21 4.39 1.3 ;
      RECT  4.74 1.455 4.97 1.555 ;
      RECT  7.2 0.205 7.32 0.635 ;
      RECT  7.2 0.635 7.785 0.725 ;
      RECT  7.675 0.725 7.785 0.84 ;
      RECT  7.2 0.725 7.31 1.015 ;
      RECT  7.2 1.015 7.415 1.115 ;
      RECT  2.965 0.23 3.055 0.845 ;
      RECT  2.965 0.845 3.095 0.98 ;
      RECT  2.815 0.98 3.095 1.08 ;
      RECT  2.815 1.08 2.905 1.175 ;
      RECT  3.465 0.215 3.565 0.95 ;
      RECT  3.395 0.95 3.565 0.97 ;
      RECT  3.395 0.97 4.21 1.06 ;
      RECT  4.11 0.83 4.21 0.97 ;
      RECT  3.395 1.06 3.49 1.285 ;
      RECT  8.14 0.19 8.23 1.085 ;
      RECT  8.14 1.085 8.495 1.175 ;
      RECT  8.405 1.005 8.495 1.085 ;
      RECT  8.14 1.175 8.23 1.265 ;
      RECT  7.275 1.265 8.23 1.36 ;
      RECT  1.675 1.11 1.98 1.225 ;
      RECT  1.675 1.225 1.805 1.615 ;
      RECT  3.59 1.15 3.77 1.25 ;
      RECT  3.59 1.25 3.69 1.525 ;
      RECT  2.71 1.525 3.69 1.64 ;
      RECT  0.07 1.38 0.19 1.445 ;
      RECT  0.07 1.445 1.325 1.535 ;
      RECT  0.07 1.535 0.285 1.55 ;
      LAYER M2 ;
      RECT  0.08 1.15 1.815 1.25 ;
      RECT  3.59 1.15 5.53 1.25 ;
      LAYER V1 ;
      RECT  0.12 1.15 0.22 1.25 ;
      RECT  1.675 1.15 1.775 1.25 ;
      RECT  3.63 1.15 3.73 1.25 ;
      RECT  5.39 1.15 5.49 1.25 ;
  END
END SEN_FSDPSBQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPSBQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPSBQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDPSBQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.05 0.69 7.15 0.945 ;
      RECT  6.95 0.945 7.15 1.115 ;
      RECT  2.4 0.71 2.615 0.89 ;
      RECT  2.4 0.89 2.49 1.05 ;
      LAYER M2 ;
      RECT  2.475 0.75 7.22 0.85 ;
      LAYER V1 ;
      RECT  7.05 0.75 7.15 0.85 ;
      RECT  2.515 0.75 2.615 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1266 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.85 0.895 ;
      LAYER M2 ;
      RECT  1.15 0.75 1.935 0.85 ;
      LAYER V1 ;
      RECT  1.35 0.75 1.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.655 0.29 8.745 0.44 ;
      RECT  8.655 0.44 9.265 0.53 ;
      RECT  9.15 0.53 9.265 1.11 ;
      RECT  8.64 1.11 9.265 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.17 0.82 8.45 0.92 ;
      RECT  8.35 0.92 8.45 1.29 ;
      RECT  4.125 0.99 4.365 1.18 ;
      RECT  4.125 1.18 4.225 1.29 ;
      LAYER M2 ;
      RECT  4.085 1.15 8.49 1.25 ;
      LAYER V1 ;
      RECT  8.35 1.15 8.45 1.25 ;
      RECT  4.125 1.15 4.225 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0834 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.89 ;
      RECT  0.35 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1035 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.66 ;
      RECT  0.55 0.66 1.05 0.76 ;
      RECT  0.95 0.76 1.05 1.02 ;
      RECT  0.95 1.02 1.165 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.575 0.45 7.75 0.69 ;
      RECT  7.575 0.69 7.665 1.575 ;
      LAYER M2 ;
      RECT  7.475 0.55 8.475 0.65 ;
      LAYER V1 ;
      RECT  7.65 0.55 7.75 0.65 ;
    END
    ANTENNADIFFAREA 0.093 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.435 0.47 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.83 1.615 1.0 1.75 ;
      RECT  2.475 1.615 2.645 1.75 ;
      RECT  4.13 1.385 4.235 1.75 ;
      RECT  4.61 1.45 4.78 1.75 ;
      RECT  5.165 1.21 5.285 1.75 ;
      RECT  5.685 1.385 5.805 1.75 ;
      RECT  7.275 1.48 7.445 1.75 ;
      RECT  7.84 1.395 7.96 1.75 ;
      RECT  8.38 1.39 8.5 1.75 ;
      RECT  8.9 1.39 9.02 1.75 ;
      RECT  9.41 1.41 9.54 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  1.665 0.05 1.835 0.18 ;
      RECT  2.24 0.05 2.42 0.18 ;
      RECT  2.82 0.05 2.99 0.18 ;
      RECT  7.3 0.05 7.47 0.18 ;
      RECT  8.875 0.05 9.045 0.32 ;
      RECT  4.09 0.05 4.26 0.345 ;
      RECT  0.365 0.05 0.505 0.38 ;
      RECT  9.41 0.05 9.54 0.39 ;
      RECT  5.685 0.05 5.805 0.435 ;
      RECT  8.355 0.05 8.525 0.515 ;
      RECT  5.16 0.05 5.28 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.33 0.165 3.44 0.27 ;
      RECT  0.845 0.27 3.44 0.36 ;
      RECT  0.845 0.36 2.31 0.37 ;
      RECT  2.925 0.36 3.015 1.135 ;
      RECT  2.22 0.37 2.31 1.22 ;
      RECT  2.925 1.135 3.445 1.23 ;
      RECT  1.445 1.22 2.31 1.31 ;
      RECT  1.445 1.31 1.615 1.36 ;
      RECT  8.045 0.16 8.145 0.27 ;
      RECT  6.755 0.27 8.145 0.36 ;
      RECT  6.755 0.36 6.845 0.415 ;
      RECT  8.055 0.36 8.145 0.62 ;
      RECT  6.22 0.415 6.845 0.505 ;
      RECT  6.22 0.505 6.31 1.315 ;
      RECT  8.055 0.62 8.67 0.71 ;
      RECT  8.58 0.71 8.67 0.785 ;
      RECT  8.58 0.785 9.04 0.895 ;
      RECT  6.22 1.315 6.88 1.405 ;
      RECT  6.76 1.405 6.88 1.635 ;
      RECT  5.96 0.21 6.655 0.305 ;
      RECT  6.485 0.305 6.655 0.32 ;
      RECT  5.96 0.305 6.05 0.53 ;
      RECT  5.425 0.375 5.545 0.53 ;
      RECT  5.425 0.53 6.05 0.62 ;
      RECT  5.96 0.62 6.05 1.06 ;
      RECT  5.375 1.06 6.05 1.18 ;
      RECT  5.96 1.18 6.05 1.495 ;
      RECT  5.96 1.495 6.63 1.6 ;
      RECT  4.35 0.215 5.07 0.32 ;
      RECT  3.6 0.19 3.805 0.36 ;
      RECT  3.715 0.36 3.805 0.73 ;
      RECT  3.715 0.73 4.63 0.82 ;
      RECT  4.54 0.82 4.63 0.915 ;
      RECT  3.945 0.82 4.035 1.54 ;
      RECT  4.54 0.915 4.77 1.015 ;
      RECT  2.97 1.54 4.035 1.66 ;
      RECT  3.895 0.475 5.0 0.565 ;
      RECT  3.895 0.565 4.065 0.6 ;
      RECT  4.91 0.565 5.0 0.765 ;
      RECT  4.91 0.765 5.85 0.875 ;
      RECT  4.91 0.875 5.0 1.27 ;
      RECT  4.38 1.27 5.0 1.36 ;
      RECT  4.91 1.36 5.0 1.54 ;
      RECT  4.38 1.36 4.48 1.605 ;
      RECT  2.51 0.49 2.805 0.58 ;
      RECT  2.705 0.58 2.805 1.14 ;
      RECT  2.47 1.14 2.805 1.23 ;
      RECT  2.47 1.23 2.56 1.4 ;
      RECT  2.18 1.4 2.56 1.525 ;
      RECT  6.96 0.485 7.48 0.585 ;
      RECT  7.39 0.585 7.48 1.26 ;
      RECT  7.04 1.26 7.48 1.35 ;
      RECT  7.04 1.35 7.16 1.615 ;
      RECT  1.115 0.475 2.12 0.595 ;
      RECT  3.105 0.545 3.625 0.665 ;
      RECT  3.535 0.665 3.625 1.35 ;
      RECT  2.72 1.35 3.625 1.45 ;
      RECT  6.65 0.71 6.96 0.83 ;
      RECT  6.65 0.83 6.755 1.135 ;
      RECT  6.65 1.135 6.82 1.225 ;
      RECT  7.875 0.45 7.965 0.965 ;
      RECT  7.8 0.965 7.965 1.045 ;
      RECT  7.8 1.045 8.235 1.135 ;
      RECT  8.12 1.135 8.235 1.615 ;
      RECT  2.04 0.695 2.13 1.0 ;
      RECT  1.265 1.0 2.13 1.09 ;
      RECT  1.265 1.09 1.355 1.255 ;
      RECT  0.065 0.2 0.185 1.255 ;
      RECT  0.065 1.255 1.355 1.345 ;
      RECT  0.065 1.345 0.185 1.59 ;
      RECT  3.755 0.91 3.855 1.37 ;
      RECT  0.56 1.435 1.395 1.475 ;
      RECT  0.56 1.475 1.9 1.525 ;
      RECT  1.305 1.525 1.9 1.575 ;
      LAYER M2 ;
      RECT  2.665 0.95 6.79 1.05 ;
      LAYER V1 ;
      RECT  2.705 0.95 2.805 1.05 ;
      RECT  3.755 0.95 3.855 1.05 ;
      RECT  6.65 0.95 6.75 1.05 ;
  END
END SEN_FSDPSBQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPSBQO_6
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPSBQO_6
  CLASS CORE ;
  FOREIGN SEN_FSDPSBQO_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.35 0.75 8.535 0.85 ;
      RECT  8.35 0.85 8.53 0.945 ;
      RECT  8.23 0.945 8.53 1.115 ;
      RECT  2.695 0.75 2.985 0.93 ;
      LAYER M2 ;
      RECT  2.805 0.75 8.535 0.85 ;
      LAYER V1 ;
      RECT  8.395 0.75 8.495 0.85 ;
      RECT  2.845 0.75 2.945 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1491 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.44 0.715 1.89 0.89 ;
      LAYER M2 ;
      RECT  1.28 0.75 2.105 0.85 ;
      LAYER V1 ;
      RECT  1.75 0.75 1.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1266 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.93 0.19 10.045 0.36 ;
      RECT  9.955 0.36 10.045 0.51 ;
      RECT  9.955 0.51 11.075 0.69 ;
      RECT  10.72 0.69 10.85 1.11 ;
      RECT  9.915 1.11 11.075 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.55 0.71 9.68 0.95 ;
      RECT  9.58 0.95 9.68 1.29 ;
      RECT  4.895 0.95 5.055 1.35 ;
      LAYER M2 ;
      RECT  4.915 1.15 9.76 1.25 ;
      LAYER V1 ;
      RECT  9.58 1.15 9.68 1.25 ;
      RECT  4.955 1.15 5.055 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.345 0.51 0.445 0.785 ;
      RECT  0.235 0.785 0.445 0.955 ;
      LAYER M2 ;
      RECT  0.305 0.55 0.845 0.65 ;
      LAYER V1 ;
      RECT  0.345 0.55 0.445 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1164 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.535 0.56 0.625 0.71 ;
      RECT  0.535 0.71 1.185 0.89 ;
      RECT  0.75 0.28 0.85 0.71 ;
      RECT  1.015 0.89 1.185 0.955 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0429 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.91 0.51 9.05 1.43 ;
      RECT  8.855 1.43 9.05 1.6 ;
    END
    ANTENNADIFFAREA 0.09 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.395 0.455 1.75 ;
      RECT  0.0 1.75 11.4 1.85 ;
      RECT  0.83 1.48 1.0 1.75 ;
      RECT  2.48 1.62 2.65 1.75 ;
      RECT  3.06 1.57 3.18 1.75 ;
      RECT  4.76 1.45 4.93 1.75 ;
      RECT  5.4 1.45 5.57 1.75 ;
      RECT  5.945 1.34 6.065 1.75 ;
      RECT  6.435 1.235 6.555 1.75 ;
      RECT  6.955 1.235 7.075 1.75 ;
      RECT  8.545 1.45 8.715 1.75 ;
      RECT  9.14 1.39 9.25 1.75 ;
      RECT  9.64 1.415 9.77 1.75 ;
      RECT  10.175 1.415 10.295 1.75 ;
      RECT  10.695 1.415 10.815 1.75 ;
      RECT  11.21 1.21 11.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.4 0.05 ;
      RECT  5.135 0.05 5.305 0.17 ;
      RECT  8.585 0.05 8.755 0.17 ;
      RECT  2.51 0.05 2.68 0.225 ;
      RECT  3.05 0.05 3.22 0.225 ;
      RECT  1.97 0.05 2.14 0.235 ;
      RECT  6.955 0.05 7.075 0.36 ;
      RECT  6.43 0.05 6.555 0.385 ;
      RECT  9.655 0.05 9.775 0.385 ;
      RECT  0.335 0.05 0.475 0.4 ;
      RECT  4.565 0.05 4.71 0.41 ;
      RECT  10.175 0.05 10.295 0.41 ;
      RECT  10.695 0.05 10.815 0.41 ;
      RECT  11.215 0.05 11.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  7.23 0.15 7.915 0.26 ;
      RECT  7.23 0.26 7.325 0.485 ;
      RECT  6.175 0.17 6.295 0.485 ;
      RECT  6.175 0.485 7.325 0.59 ;
      RECT  7.235 0.59 7.325 1.025 ;
      RECT  6.125 1.025 7.325 1.145 ;
      RECT  7.235 1.145 7.325 1.495 ;
      RECT  7.235 1.495 7.91 1.595 ;
      RECT  1.155 0.24 1.845 0.325 ;
      RECT  1.155 0.325 2.435 0.34 ;
      RECT  1.725 0.34 2.435 0.445 ;
      RECT  3.91 0.215 4.33 0.335 ;
      RECT  4.24 0.335 4.33 0.77 ;
      RECT  4.24 0.77 5.425 0.86 ;
      RECT  5.335 0.86 5.425 0.95 ;
      RECT  4.535 0.86 4.625 1.57 ;
      RECT  5.335 0.95 5.63 1.04 ;
      RECT  3.52 1.57 4.625 1.66 ;
      RECT  8.035 0.265 9.47 0.355 ;
      RECT  8.035 0.355 8.125 0.395 ;
      RECT  9.38 0.355 9.47 0.505 ;
      RECT  7.425 0.395 8.125 0.51 ;
      RECT  9.38 0.505 9.865 0.595 ;
      RECT  7.425 0.51 7.52 1.315 ;
      RECT  9.77 0.595 9.865 0.78 ;
      RECT  9.77 0.78 10.615 0.89 ;
      RECT  7.425 1.315 8.125 1.405 ;
      RECT  8.035 1.405 8.125 1.635 ;
      RECT  0.055 0.2 0.17 0.395 ;
      RECT  0.055 0.395 0.145 1.045 ;
      RECT  0.055 1.045 2.195 1.135 ;
      RECT  2.105 0.715 2.195 1.045 ;
      RECT  0.055 1.135 0.17 1.61 ;
      RECT  4.825 0.275 5.855 0.395 ;
      RECT  2.565 0.315 3.805 0.405 ;
      RECT  3.265 0.405 3.805 0.415 ;
      RECT  2.565 0.405 2.655 0.535 ;
      RECT  3.685 0.415 3.805 0.54 ;
      RECT  3.265 0.415 3.355 1.21 ;
      RECT  0.955 0.295 1.055 0.43 ;
      RECT  0.955 0.43 1.61 0.535 ;
      RECT  1.48 0.535 2.655 0.625 ;
      RECT  2.285 0.625 2.375 1.24 ;
      RECT  3.265 1.21 3.995 1.3 ;
      RECT  1.935 1.24 2.375 1.27 ;
      RECT  1.39 1.27 2.375 1.33 ;
      RECT  1.39 1.33 2.085 1.39 ;
      RECT  8.33 0.455 8.43 0.54 ;
      RECT  8.33 0.54 8.82 0.635 ;
      RECT  8.67 0.635 8.82 0.89 ;
      RECT  8.67 0.89 8.76 1.27 ;
      RECT  8.305 1.27 8.76 1.36 ;
      RECT  8.305 1.36 8.395 1.635 ;
      RECT  4.47 0.51 6.05 0.63 ;
      RECT  4.47 0.63 4.56 0.68 ;
      RECT  5.945 0.63 6.05 0.77 ;
      RECT  5.945 0.77 6.885 0.79 ;
      RECT  5.74 0.79 6.885 0.88 ;
      RECT  5.74 0.88 5.83 1.27 ;
      RECT  5.18 1.27 5.83 1.36 ;
      RECT  5.66 1.36 5.83 1.41 ;
      RECT  5.18 1.36 5.27 1.535 ;
      RECT  2.755 0.52 3.175 0.64 ;
      RECT  3.075 0.64 3.175 1.16 ;
      RECT  2.53 1.16 3.175 1.275 ;
      RECT  2.53 1.275 2.62 1.43 ;
      RECT  2.17 1.43 2.62 1.53 ;
      RECT  3.455 0.51 3.57 0.655 ;
      RECT  3.455 0.655 4.14 0.745 ;
      RECT  4.05 0.745 4.14 0.97 ;
      RECT  4.05 0.97 4.175 1.1 ;
      RECT  4.085 1.1 4.175 1.39 ;
      RECT  2.74 1.39 4.175 1.48 ;
      RECT  9.14 0.51 9.25 0.68 ;
      RECT  9.145 0.68 9.25 1.075 ;
      RECT  9.145 1.075 9.49 1.165 ;
      RECT  9.4 1.165 9.49 1.62 ;
      RECT  8.12 0.66 8.225 0.725 ;
      RECT  7.895 0.725 8.225 0.855 ;
      RECT  7.895 0.855 8.01 1.135 ;
      RECT  7.895 1.135 8.07 1.225 ;
      RECT  4.265 0.95 4.445 1.05 ;
      RECT  4.285 1.05 4.445 1.38 ;
      RECT  0.545 1.275 1.3 1.39 ;
      RECT  1.2 1.39 1.3 1.48 ;
      RECT  1.2 1.48 1.87 1.6 ;
      LAYER M2 ;
      RECT  3.035 0.95 8.035 1.05 ;
      LAYER V1 ;
      RECT  3.075 0.95 3.175 1.05 ;
      RECT  4.305 0.95 4.405 1.05 ;
      RECT  7.895 0.95 7.995 1.05 ;
  END
END SEN_FSDPSBQO_6
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPSBQO_8
#      Description : "D-Flip Flop w/scan, pos-edge triggered, lo-async-set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=(!SE&D)|(SE&SI),preset=!SD):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPSBQO_8
  CLASS CORE ;
  FOREIGN SEN_FSDPSBQO_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.975 0.75 9.155 1.005 ;
      RECT  8.865 1.005 9.155 1.175 ;
      RECT  8.19 0.635 8.29 1.175 ;
      RECT  2.95 0.69 3.095 1.09 ;
      LAYER M2 ;
      RECT  2.945 0.75 9.155 0.85 ;
      LAYER V1 ;
      RECT  9.015 0.75 9.115 0.85 ;
      RECT  8.19 0.75 8.29 0.85 ;
      RECT  2.985 0.75 3.085 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.145 0.75 1.6 0.85 ;
      LAYER M2 ;
      RECT  1.42 0.75 2.09 0.85 ;
      LAYER V1 ;
      RECT  1.46 0.75 1.56 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.58 0.19 10.745 0.36 ;
      RECT  10.655 0.36 10.745 0.51 ;
      RECT  10.655 0.51 12.25 0.69 ;
      RECT  11.68 0.69 11.85 1.11 ;
      RECT  10.55 1.11 12.25 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END Q
  PIN SD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.23 0.725 10.33 1.31 ;
      RECT  4.935 0.98 5.115 1.25 ;
      LAYER M2 ;
      RECT  4.935 1.15 10.4 1.25 ;
      LAYER V1 ;
      RECT  10.23 1.15 10.33 1.25 ;
      RECT  4.975 1.15 5.075 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END SD
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.49 0.45 0.97 ;
      RECT  0.35 0.97 0.58 1.07 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1188 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.49 0.655 0.7 ;
      RECT  0.55 0.7 0.85 0.79 ;
      RECT  0.75 0.79 0.85 0.965 ;
      RECT  0.75 0.965 1.635 1.07 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0474 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.53 0.44 9.65 1.605 ;
    END
    ANTENNADIFFAREA 0.093 ;
  END SO
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.37 0.445 1.75 ;
      RECT  0.0 1.75 12.6 1.85 ;
      RECT  0.845 1.61 1.015 1.75 ;
      RECT  1.415 1.355 1.535 1.75 ;
      RECT  2.98 1.44 3.15 1.75 ;
      RECT  3.545 1.55 3.66 1.75 ;
      RECT  4.83 1.375 4.94 1.75 ;
      RECT  5.58 1.42 5.71 1.75 ;
      RECT  6.105 1.33 6.235 1.75 ;
      RECT  6.63 1.38 6.755 1.75 ;
      RECT  7.155 1.38 7.275 1.75 ;
      RECT  9.23 1.445 9.4 1.75 ;
      RECT  9.77 1.39 9.895 1.75 ;
      RECT  10.3 1.42 10.43 1.75 ;
      RECT  10.825 1.39 10.945 1.75 ;
      RECT  11.345 1.39 11.465 1.75 ;
      RECT  11.865 1.39 11.985 1.75 ;
      RECT  12.4 1.21 12.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.6 0.05 ;
      RECT  5.335 0.05 5.505 0.17 ;
      RECT  9.215 0.05 9.385 0.17 ;
      RECT  2.16 0.05 2.33 0.21 ;
      RECT  7.09 0.05 7.26 0.345 ;
      RECT  0.335 0.05 0.505 0.36 ;
      RECT  10.305 0.05 10.425 0.36 ;
      RECT  2.715 0.05 2.835 0.365 ;
      RECT  1.63 0.05 1.8 0.37 ;
      RECT  3.275 0.05 3.395 0.37 ;
      RECT  7.635 0.05 7.74 0.375 ;
      RECT  10.84 0.05 10.955 0.385 ;
      RECT  11.34 0.05 11.47 0.385 ;
      RECT  11.86 0.05 11.99 0.385 ;
      RECT  4.815 0.05 4.935 0.41 ;
      RECT  12.4 0.05 12.52 0.59 ;
      RECT  6.595 0.05 6.715 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.9 0.16 1.51 0.25 ;
      RECT  1.42 0.25 1.51 0.385 ;
      RECT  0.9 0.25 1.07 0.41 ;
      RECT  0.97 0.41 1.07 0.69 ;
      RECT  3.8 0.195 4.445 0.31 ;
      RECT  4.325 0.31 4.445 0.43 ;
      RECT  3.8 0.31 3.915 0.48 ;
      RECT  4.325 0.43 4.535 0.53 ;
      RECT  4.43 0.53 4.535 0.71 ;
      RECT  4.43 0.71 4.74 0.745 ;
      RECT  4.43 0.745 5.75 0.8 ;
      RECT  4.65 0.8 5.75 0.855 ;
      RECT  4.65 0.855 4.74 1.55 ;
      RECT  3.75 1.55 4.74 1.64 ;
      RECT  7.83 0.215 8.585 0.325 ;
      RECT  7.83 0.325 7.92 0.465 ;
      RECT  6.825 0.465 7.92 0.555 ;
      RECT  6.825 0.555 7.56 0.585 ;
      RECT  7.425 0.585 7.56 1.115 ;
      RECT  6.32 1.115 7.56 1.235 ;
      RECT  7.425 1.235 7.56 1.48 ;
      RECT  7.425 1.48 8.61 1.62 ;
      RECT  1.93 0.185 2.02 0.33 ;
      RECT  1.93 0.33 2.575 0.42 ;
      RECT  2.455 0.17 2.575 0.33 ;
      RECT  1.93 0.42 2.02 0.48 ;
      RECT  1.16 0.34 1.25 0.48 ;
      RECT  1.16 0.48 2.02 0.57 ;
      RECT  8.68 0.26 10.075 0.35 ;
      RECT  8.68 0.35 8.79 0.415 ;
      RECT  9.985 0.35 10.075 0.45 ;
      RECT  8.01 0.415 8.79 0.52 ;
      RECT  9.985 0.45 10.565 0.54 ;
      RECT  8.01 0.52 8.1 1.27 ;
      RECT  10.475 0.54 10.565 0.785 ;
      RECT  10.475 0.785 11.575 0.89 ;
      RECT  7.65 1.27 8.815 1.39 ;
      RECT  8.71 1.39 8.815 1.615 ;
      RECT  5.05 0.26 6.49 0.36 ;
      RECT  4.04 0.415 4.21 0.505 ;
      RECT  4.04 0.505 4.15 1.41 ;
      RECT  5.54 0.45 6.23 0.51 ;
      RECT  4.635 0.51 6.23 0.54 ;
      RECT  4.635 0.54 5.71 0.6 ;
      RECT  6.14 0.54 6.23 0.76 ;
      RECT  5.86 0.76 7.295 0.865 ;
      RECT  5.86 0.865 5.965 1.24 ;
      RECT  5.23 1.24 5.965 1.33 ;
      RECT  5.84 1.33 5.965 1.51 ;
      RECT  5.23 1.33 5.36 1.575 ;
      RECT  8.92 0.48 9.44 0.595 ;
      RECT  9.35 0.595 9.44 1.265 ;
      RECT  8.955 1.265 9.44 1.355 ;
      RECT  8.955 1.355 9.075 1.615 ;
      RECT  2.95 0.49 3.33 0.6 ;
      RECT  3.23 0.6 3.33 1.19 ;
      RECT  2.925 1.19 3.33 1.22 ;
      RECT  2.665 1.22 3.33 1.28 ;
      RECT  2.665 1.28 2.995 1.35 ;
      RECT  3.58 0.52 3.71 0.69 ;
      RECT  3.62 0.69 3.71 0.95 ;
      RECT  3.62 0.95 3.87 1.04 ;
      RECT  3.62 1.04 3.71 1.37 ;
      RECT  3.275 1.37 3.71 1.46 ;
      RECT  3.275 1.46 3.395 1.58 ;
      RECT  2.575 0.51 2.665 0.735 ;
      RECT  1.755 0.735 2.665 0.825 ;
      RECT  1.755 0.825 1.855 1.16 ;
      RECT  0.065 0.19 0.185 1.16 ;
      RECT  0.065 1.16 1.855 1.26 ;
      RECT  0.065 1.26 0.185 1.585 ;
      RECT  8.38 0.715 8.885 0.81 ;
      RECT  8.795 0.81 8.885 0.885 ;
      RECT  8.38 0.81 8.48 1.15 ;
      RECT  2.755 0.455 2.855 1.0 ;
      RECT  1.945 1.0 2.855 1.115 ;
      RECT  1.945 1.115 2.035 1.41 ;
      RECT  9.79 0.455 9.885 1.045 ;
      RECT  9.79 1.045 10.14 1.135 ;
      RECT  10.035 1.135 10.14 1.62 ;
      RECT  4.46 0.91 4.56 1.455 ;
      RECT  0.535 1.35 1.3 1.465 ;
      RECT  2.165 1.34 2.55 1.51 ;
      LAYER M2 ;
      RECT  0.93 0.55 4.18 0.65 ;
      RECT  3.19 0.95 8.52 1.05 ;
      RECT  1.11 1.35 2.35 1.45 ;
      LAYER V1 ;
      RECT  0.97 0.55 1.07 0.65 ;
      RECT  2.755 0.55 2.855 0.65 ;
      RECT  4.04 0.55 4.14 0.65 ;
      RECT  3.23 0.95 3.33 1.05 ;
      RECT  4.46 0.95 4.56 1.05 ;
      RECT  8.38 0.95 8.48 1.05 ;
      RECT  1.16 1.35 1.26 1.45 ;
      RECT  2.205 1.35 2.305 1.45 ;
  END
END SEN_FSDPSBQO_8
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPTQ_D_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, hi-sync-set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&(D|SS))|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPTQ_D_1
  CLASS CORE ;
  FOREIGN SEN_FSDPTQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.975 0.69 4.35 0.785 ;
      RECT  4.25 0.785 4.35 1.03 ;
      RECT  4.25 1.03 4.605 1.2 ;
      RECT  3.35 0.71 3.68 0.89 ;
      RECT  2.95 0.47 3.05 0.89 ;
      LAYER M2 ;
      RECT  2.91 0.75 4.39 0.85 ;
      LAYER V1 ;
      RECT  4.25 0.75 4.35 0.85 ;
      RECT  3.555 0.75 3.655 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1176 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.625 0.45 5.73 1.11 ;
      RECT  5.55 1.11 5.73 1.2 ;
      RECT  5.55 1.2 5.65 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.915 0.805 2.015 1.225 ;
      RECT  0.395 0.505 0.65 0.61 ;
      RECT  0.55 0.61 0.65 0.95 ;
      RECT  0.55 0.95 0.86 1.05 ;
      LAYER M2 ;
      RECT  0.68 0.95 2.055 1.05 ;
      LAYER V1 ;
      RECT  1.915 0.95 2.015 1.05 ;
      RECT  0.72 0.95 0.82 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.7 1.055 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END SS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.495 1.44 0.62 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  2.02 1.505 2.19 1.75 ;
      RECT  3.565 1.48 3.685 1.75 ;
      RECT  4.83 1.47 5.0 1.75 ;
      RECT  5.35 1.13 5.455 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  1.835 0.05 1.955 0.31 ;
      RECT  0.325 0.05 0.445 0.38 ;
      RECT  3.32 0.05 3.425 0.4 ;
      RECT  5.35 0.05 5.47 0.56 ;
      RECT  4.84 0.05 4.96 0.58 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.565 0.14 4.6 0.23 ;
      RECT  3.565 0.23 3.685 0.49 ;
      RECT  2.28 0.14 3.23 0.23 ;
      RECT  2.28 0.23 2.385 0.31 ;
      RECT  3.14 0.23 3.23 0.49 ;
      RECT  3.14 0.49 3.685 0.58 ;
      RECT  3.14 0.58 3.23 0.99 ;
      RECT  3.065 0.99 3.23 1.105 ;
      RECT  3.065 1.105 3.98 1.21 ;
      RECT  1.0 0.24 1.735 0.355 ;
      RECT  0.795 0.2 0.91 0.445 ;
      RECT  0.795 0.445 2.62 0.52 ;
      RECT  1.83 0.4 2.62 0.445 ;
      RECT  0.795 0.52 1.915 0.56 ;
      RECT  3.79 0.425 3.99 0.545 ;
      RECT  3.79 0.545 3.88 0.91 ;
      RECT  3.79 0.91 4.16 1.0 ;
      RECT  4.07 1.0 4.16 1.29 ;
      RECT  4.07 1.29 4.23 1.3 ;
      RECT  2.12 0.62 2.21 1.145 ;
      RECT  2.12 1.145 2.65 1.235 ;
      RECT  2.56 1.235 2.65 1.3 ;
      RECT  2.56 1.3 4.23 1.39 ;
      RECT  3.245 1.39 3.335 1.62 ;
      RECT  4.125 0.425 4.7 0.545 ;
      RECT  4.61 0.545 4.7 0.74 ;
      RECT  4.61 0.74 4.785 0.83 ;
      RECT  4.695 0.83 4.785 1.25 ;
      RECT  4.695 1.25 5.12 1.29 ;
      RECT  4.345 1.29 5.12 1.38 ;
      RECT  4.345 1.38 4.465 1.61 ;
      RECT  2.74 0.33 2.83 0.805 ;
      RECT  2.3 0.805 2.83 0.895 ;
      RECT  2.3 0.895 2.395 1.035 ;
      RECT  2.74 0.895 2.83 1.04 ;
      RECT  2.74 1.04 2.94 1.21 ;
      RECT  5.09 0.315 5.21 0.81 ;
      RECT  4.895 0.81 5.21 0.85 ;
      RECT  4.895 0.85 5.535 0.92 ;
      RECT  5.435 0.725 5.535 0.85 ;
      RECT  5.09 0.92 5.535 0.955 ;
      RECT  5.09 0.955 5.21 1.16 ;
      RECT  1.675 1.0 1.78 1.08 ;
      RECT  1.38 1.08 1.78 1.17 ;
      RECT  1.38 1.17 1.47 1.465 ;
      RECT  0.065 0.195 0.17 1.21 ;
      RECT  0.065 1.21 0.82 1.3 ;
      RECT  0.73 1.3 0.82 1.465 ;
      RECT  0.195 1.3 0.315 1.61 ;
      RECT  0.73 1.465 1.47 1.555 ;
      RECT  1.56 1.325 2.47 1.415 ;
      RECT  2.38 1.415 2.47 1.48 ;
      RECT  1.56 1.415 1.685 1.615 ;
      RECT  2.38 1.48 2.73 1.585 ;
  END
END SEN_FSDPTQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPTQ_D_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, hi-sync-set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&(D|SS))|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPTQ_D_2
  CLASS CORE ;
  FOREIGN SEN_FSDPTQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.975 0.69 4.35 0.785 ;
      RECT  4.25 0.785 4.35 1.03 ;
      RECT  4.25 1.03 4.605 1.2 ;
      RECT  3.35 0.71 3.68 0.89 ;
      RECT  2.95 0.47 3.05 0.89 ;
      LAYER M2 ;
      RECT  2.91 0.75 4.39 0.85 ;
      LAYER V1 ;
      RECT  4.25 0.75 4.35 0.85 ;
      RECT  3.555 0.75 3.655 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1176 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.575 0.455 6.05 0.575 ;
      RECT  5.95 0.575 6.05 1.11 ;
      RECT  5.635 1.11 6.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.915 0.805 2.015 1.225 ;
      RECT  0.395 0.505 0.65 0.61 ;
      RECT  0.55 0.61 0.65 0.95 ;
      RECT  0.55 0.95 0.86 1.05 ;
      LAYER M2 ;
      RECT  0.68 0.95 2.055 1.05 ;
      LAYER V1 ;
      RECT  1.915 0.95 2.015 1.05 ;
      RECT  0.72 0.95 0.82 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.7 1.055 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END SS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.49 1.39 0.62 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  2.02 1.505 2.19 1.75 ;
      RECT  3.565 1.48 3.685 1.75 ;
      RECT  4.83 1.47 5.0 1.75 ;
      RECT  5.36 1.19 5.48 1.75 ;
      RECT  5.905 1.41 6.035 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  1.835 0.05 1.955 0.31 ;
      RECT  5.905 0.05 6.035 0.36 ;
      RECT  3.32 0.05 3.425 0.4 ;
      RECT  0.325 0.05 0.445 0.415 ;
      RECT  5.36 0.05 5.48 0.56 ;
      RECT  4.84 0.05 4.96 0.595 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.565 0.14 4.6 0.23 ;
      RECT  3.565 0.23 3.685 0.49 ;
      RECT  2.29 0.14 3.23 0.23 ;
      RECT  2.29 0.23 2.385 0.31 ;
      RECT  3.14 0.23 3.23 0.49 ;
      RECT  3.14 0.49 3.685 0.58 ;
      RECT  3.14 0.58 3.23 0.99 ;
      RECT  3.055 0.99 3.23 1.095 ;
      RECT  3.055 1.095 3.98 1.21 ;
      RECT  1.005 0.24 1.735 0.355 ;
      RECT  0.795 0.205 0.915 0.445 ;
      RECT  0.795 0.445 2.62 0.52 ;
      RECT  1.83 0.4 2.62 0.445 ;
      RECT  0.795 0.52 1.915 0.56 ;
      RECT  3.79 0.425 3.985 0.545 ;
      RECT  3.79 0.545 3.88 0.9 ;
      RECT  3.79 0.9 4.16 0.99 ;
      RECT  4.07 0.99 4.16 1.29 ;
      RECT  4.07 1.29 4.23 1.3 ;
      RECT  2.12 0.62 2.21 1.13 ;
      RECT  2.12 1.13 2.65 1.235 ;
      RECT  2.56 1.235 2.65 1.3 ;
      RECT  2.56 1.3 4.23 1.39 ;
      RECT  3.245 1.39 3.335 1.65 ;
      RECT  4.1 0.425 4.75 0.545 ;
      RECT  4.66 0.545 4.75 0.74 ;
      RECT  4.66 0.74 4.785 0.83 ;
      RECT  4.695 0.83 4.785 1.25 ;
      RECT  4.695 1.25 5.115 1.29 ;
      RECT  4.345 1.29 5.115 1.38 ;
      RECT  4.345 1.38 4.465 1.61 ;
      RECT  5.09 0.45 5.21 0.785 ;
      RECT  5.09 0.785 5.75 0.825 ;
      RECT  4.875 0.825 5.75 0.89 ;
      RECT  4.875 0.89 5.21 0.995 ;
      RECT  5.105 0.995 5.21 1.16 ;
      RECT  2.725 0.33 2.845 0.805 ;
      RECT  2.3 0.805 2.845 0.895 ;
      RECT  2.3 0.895 2.395 1.035 ;
      RECT  2.74 0.895 2.845 1.04 ;
      RECT  2.74 1.04 2.94 1.21 ;
      RECT  1.675 1.025 1.78 1.135 ;
      RECT  1.385 1.135 1.78 1.225 ;
      RECT  1.385 1.225 1.475 1.465 ;
      RECT  0.065 0.2 0.17 1.21 ;
      RECT  0.065 1.21 0.835 1.3 ;
      RECT  0.745 1.3 0.835 1.465 ;
      RECT  0.195 1.3 0.315 1.615 ;
      RECT  0.745 1.465 1.475 1.555 ;
      RECT  1.565 1.325 2.47 1.415 ;
      RECT  2.38 1.415 2.47 1.48 ;
      RECT  1.565 1.415 1.685 1.595 ;
      RECT  2.38 1.48 2.735 1.585 ;
  END
END SEN_FSDPTQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPTQ_D_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, hi-sync-set, q-only"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&(D|SS))|(SE&SI))):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPTQ_D_4
  CLASS CORE ;
  FOREIGN SEN_FSDPTQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.975 0.69 4.35 0.785 ;
      RECT  4.25 0.785 4.35 1.03 ;
      RECT  4.25 1.03 4.605 1.2 ;
      RECT  3.35 0.71 3.68 0.89 ;
      RECT  2.95 0.47 3.05 0.89 ;
      LAYER M2 ;
      RECT  2.91 0.75 4.39 0.85 ;
      LAYER V1 ;
      RECT  4.25 0.75 4.35 0.85 ;
      RECT  3.555 0.75 3.655 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1176 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.57 0.455 6.25 0.575 ;
      RECT  6.15 0.575 6.25 1.11 ;
      RECT  5.615 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.915 0.805 2.015 1.225 ;
      RECT  0.37 0.505 0.65 0.61 ;
      RECT  0.55 0.61 0.65 0.95 ;
      RECT  0.55 0.95 0.86 1.05 ;
      LAYER M2 ;
      RECT  0.68 0.95 2.055 1.05 ;
      LAYER V1 ;
      RECT  1.915 0.95 2.015 1.05 ;
      RECT  0.72 0.95 0.82 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.685 1.055 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END SS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.49 1.39 0.62 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  2.02 1.505 2.19 1.75 ;
      RECT  3.565 1.48 3.685 1.75 ;
      RECT  4.83 1.47 5.0 1.75 ;
      RECT  5.36 1.215 5.48 1.75 ;
      RECT  5.88 1.38 6.0 1.75 ;
      RECT  6.41 1.21 6.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.835 0.05 1.955 0.31 ;
      RECT  5.88 0.05 6.0 0.36 ;
      RECT  3.32 0.05 3.425 0.4 ;
      RECT  0.325 0.05 0.445 0.41 ;
      RECT  5.36 0.05 5.48 0.56 ;
      RECT  4.84 0.05 4.96 0.58 ;
      RECT  6.41 0.05 6.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  3.565 0.14 4.595 0.23 ;
      RECT  3.565 0.23 3.685 0.49 ;
      RECT  2.29 0.14 3.23 0.23 ;
      RECT  2.29 0.23 2.385 0.31 ;
      RECT  3.14 0.23 3.23 0.49 ;
      RECT  3.14 0.49 3.685 0.58 ;
      RECT  3.14 0.58 3.23 0.99 ;
      RECT  3.065 0.99 3.23 1.105 ;
      RECT  3.065 1.105 3.98 1.21 ;
      RECT  1.005 0.24 1.735 0.355 ;
      RECT  0.8 0.205 0.91 0.445 ;
      RECT  0.8 0.445 2.62 0.52 ;
      RECT  1.83 0.4 2.62 0.445 ;
      RECT  0.8 0.52 1.915 0.56 ;
      RECT  3.79 0.425 3.985 0.545 ;
      RECT  3.79 0.545 3.88 0.91 ;
      RECT  3.79 0.91 4.16 1.0 ;
      RECT  4.07 1.0 4.16 1.29 ;
      RECT  4.07 1.29 4.23 1.3 ;
      RECT  2.12 0.62 2.21 1.125 ;
      RECT  2.12 1.125 2.65 1.235 ;
      RECT  2.56 1.235 2.65 1.3 ;
      RECT  2.56 1.3 4.23 1.39 ;
      RECT  3.245 1.39 3.335 1.65 ;
      RECT  4.11 0.425 4.75 0.545 ;
      RECT  4.66 0.545 4.75 0.74 ;
      RECT  4.66 0.74 4.785 0.83 ;
      RECT  4.695 0.83 4.785 1.25 ;
      RECT  4.695 1.25 5.115 1.29 ;
      RECT  4.345 1.29 5.115 1.38 ;
      RECT  4.345 1.38 4.465 1.61 ;
      RECT  5.09 0.45 5.21 0.785 ;
      RECT  5.09 0.785 6.045 0.825 ;
      RECT  4.875 0.825 6.045 0.89 ;
      RECT  4.875 0.89 5.21 0.995 ;
      RECT  5.09 0.995 5.21 1.16 ;
      RECT  2.725 0.335 2.83 0.805 ;
      RECT  2.3 0.805 2.83 0.895 ;
      RECT  2.3 0.895 2.395 1.035 ;
      RECT  2.74 0.895 2.83 1.04 ;
      RECT  2.74 1.04 2.925 1.21 ;
      RECT  1.675 1.025 1.78 1.135 ;
      RECT  1.385 1.135 1.78 1.225 ;
      RECT  1.385 1.225 1.475 1.465 ;
      RECT  0.065 0.2 0.17 1.21 ;
      RECT  0.065 1.21 0.835 1.3 ;
      RECT  0.745 1.3 0.835 1.465 ;
      RECT  0.195 1.3 0.315 1.615 ;
      RECT  0.745 1.465 1.475 1.555 ;
      RECT  1.565 1.325 2.47 1.415 ;
      RECT  2.38 1.415 2.47 1.48 ;
      RECT  1.565 1.415 1.685 1.605 ;
      RECT  2.38 1.48 2.735 1.585 ;
  END
END SEN_FSDPTQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPTQO_1
#      Description : "D-Flip Flop w/scan, pos-edge triggered, hi-sync-set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&(D|SS))|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPTQO_1
  CLASS CORE ;
  FOREIGN SEN_FSDPTQO_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.635 0.745 4.735 0.91 ;
      RECT  4.635 0.91 5.18 1.09 ;
      RECT  3.78 0.78 3.96 1.05 ;
      LAYER M2 ;
      RECT  3.78 0.95 4.775 1.05 ;
      LAYER V1 ;
      RECT  4.635 0.95 4.735 1.05 ;
      RECT  3.82 0.95 3.92 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0699 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0621 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.31 6.85 1.29 ;
    END
    ANTENNADIFFAREA 0.178 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.78 ;
      RECT  0.345 0.78 0.85 0.905 ;
      RECT  0.75 0.905 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.845 0.51 1.945 1.1 ;
      RECT  0.415 0.47 0.72 0.585 ;
      RECT  0.415 0.585 0.515 0.69 ;
      LAYER M2 ;
      RECT  0.375 0.55 1.985 0.65 ;
      LAYER V1 ;
      RECT  1.845 0.55 1.945 0.65 ;
      RECT  0.415 0.55 0.515 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0246 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.31 6.25 1.29 ;
    END
    ANTENNADIFFAREA 0.117 ;
  END SO
  PIN SS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.68 1.06 1.33 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0621 ;
  END SS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.485 1.44 0.615 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  1.995 1.43 2.115 1.75 ;
      RECT  3.365 1.51 3.535 1.75 ;
      RECT  4.19 1.39 4.31 1.75 ;
      RECT  5.51 1.61 5.68 1.75 ;
      RECT  5.85 1.61 6.02 1.75 ;
      RECT  6.44 1.22 6.56 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  4.19 0.05 4.31 0.225 ;
      RECT  5.375 0.05 5.495 0.255 ;
      RECT  5.875 0.05 5.995 0.255 ;
      RECT  3.37 0.05 3.49 0.33 ;
      RECT  1.885 0.05 1.99 0.365 ;
      RECT  0.325 0.05 0.445 0.38 ;
      RECT  6.475 0.05 6.595 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  4.65 0.14 5.02 0.23 ;
      RECT  4.93 0.23 5.02 0.31 ;
      RECT  4.65 0.23 4.74 0.315 ;
      RECT  3.88 0.315 4.74 0.405 ;
      RECT  3.88 0.405 4.14 0.435 ;
      RECT  4.05 0.435 4.14 0.6 ;
      RECT  3.57 0.6 4.14 0.69 ;
      RECT  3.57 0.69 3.67 0.94 ;
      RECT  4.05 0.69 4.14 1.15 ;
      RECT  3.895 1.15 4.14 1.24 ;
      RECT  2.08 0.18 2.695 0.27 ;
      RECT  2.575 0.27 2.695 0.46 ;
      RECT  2.08 0.27 2.17 1.25 ;
      RECT  0.81 0.19 0.915 0.435 ;
      RECT  0.81 0.435 1.71 0.555 ;
      RECT  1.62 0.555 1.71 1.25 ;
      RECT  1.62 1.25 2.515 1.34 ;
      RECT  1.62 1.34 1.71 1.425 ;
      RECT  2.425 1.34 2.515 1.495 ;
      RECT  1.43 1.425 1.71 1.545 ;
      RECT  2.425 1.495 2.7 1.6 ;
      RECT  1.005 0.22 1.795 0.33 ;
      RECT  3.67 0.295 3.79 0.42 ;
      RECT  3.39 0.42 3.79 0.51 ;
      RECT  3.39 0.51 3.48 0.71 ;
      RECT  2.965 0.71 3.48 0.88 ;
      RECT  3.39 0.88 3.48 1.15 ;
      RECT  3.39 1.15 3.805 1.24 ;
      RECT  5.105 0.345 6.05 0.435 ;
      RECT  5.105 0.435 5.225 0.6 ;
      RECT  5.95 0.435 6.05 1.415 ;
      RECT  5.175 1.415 6.05 1.52 ;
      RECT  2.785 0.305 2.955 0.475 ;
      RECT  2.785 0.475 2.875 0.71 ;
      RECT  2.46 0.71 2.875 0.8 ;
      RECT  2.46 0.8 2.56 0.94 ;
      RECT  2.785 0.8 2.875 1.03 ;
      RECT  2.785 1.03 2.91 1.2 ;
      RECT  5.45 0.525 5.75 0.62 ;
      RECT  5.45 0.62 5.545 1.03 ;
      RECT  5.45 1.03 5.635 1.12 ;
      RECT  4.425 0.52 4.68 0.64 ;
      RECT  4.425 0.64 4.515 1.245 ;
      RECT  4.425 1.245 4.87 1.365 ;
      RECT  4.825 0.435 4.93 0.69 ;
      RECT  4.825 0.69 5.36 0.78 ;
      RECT  5.27 0.78 5.36 1.21 ;
      RECT  4.96 1.21 5.825 1.3 ;
      RECT  5.725 0.71 5.825 1.21 ;
      RECT  4.96 1.3 5.085 1.6 ;
      RECT  2.26 0.39 2.37 1.07 ;
      RECT  2.26 1.07 2.695 1.16 ;
      RECT  2.605 1.16 2.695 1.315 ;
      RECT  2.605 1.315 3.265 1.33 ;
      RECT  2.605 1.33 3.93 1.405 ;
      RECT  3.175 1.405 3.93 1.42 ;
      RECT  3.175 1.42 3.265 1.59 ;
      RECT  3.82 1.42 3.93 1.66 ;
      RECT  6.425 0.69 6.525 1.13 ;
      RECT  1.44 1.11 1.53 1.22 ;
      RECT  1.2 1.22 1.53 1.31 ;
      RECT  1.2 1.31 1.29 1.44 ;
      RECT  0.065 0.19 0.185 1.22 ;
      RECT  0.065 1.22 0.84 1.31 ;
      RECT  0.065 1.31 0.31 1.32 ;
      RECT  0.75 1.31 0.84 1.44 ;
      RECT  0.19 1.32 0.31 1.61 ;
      RECT  0.75 1.44 1.29 1.53 ;
      LAYER M2 ;
      RECT  5.685 0.75 6.6 0.85 ;
      LAYER V1 ;
      RECT  5.725 0.75 5.825 0.85 ;
      RECT  6.425 0.75 6.525 0.85 ;
  END
END SEN_FSDPTQO_1
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPTQO_2
#      Description : "D-Flip Flop w/scan, pos-edge triggered, hi-sync-set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&(D|SS))|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPTQO_2
  CLASS CORE ;
  FOREIGN SEN_FSDPTQO_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.275 0.47 7.375 0.89 ;
      RECT  6.67 0.6 6.805 0.925 ;
      RECT  5.35 0.51 5.45 0.71 ;
      RECT  5.35 0.71 5.615 0.875 ;
      LAYER M2 ;
      RECT  5.395 0.75 7.415 0.85 ;
      LAYER V1 ;
      RECT  7.275 0.75 7.375 0.85 ;
      RECT  6.705 0.75 6.805 0.85 ;
      RECT  5.435 0.75 5.535 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0915 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.1 0.71 3.05 0.86 ;
      RECT  2.95 0.86 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.75 0.51 9.05 0.69 ;
      RECT  8.95 0.69 9.05 1.11 ;
      RECT  8.75 1.11 9.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.205 ;
      RECT  0.55 1.205 2.405 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.087 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0306 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.86 0.495 8.07 0.6 ;
      RECT  7.95 0.6 8.07 0.94 ;
      RECT  7.875 0.94 8.07 1.045 ;
    END
    ANTENNADIFFAREA 0.134 ;
  END SO
  PIN SS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.91 ;
      RECT  0.75 0.91 1.05 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END SS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.61 0.495 1.75 ;
      RECT  0.0 1.75 9.2 1.85 ;
      RECT  2.215 1.42 2.33 1.75 ;
      RECT  3.16 1.41 3.285 1.75 ;
      RECT  4.705 1.435 4.875 1.75 ;
      RECT  5.255 1.435 5.425 1.75 ;
      RECT  6.045 1.615 6.215 1.75 ;
      RECT  7.615 1.6 7.785 1.75 ;
      RECT  8.47 1.495 8.64 1.75 ;
      RECT  9.0 1.41 9.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.2 0.05 ;
      RECT  2.6 0.05 2.77 0.195 ;
      RECT  7.615 0.05 7.785 0.195 ;
      RECT  4.715 0.05 4.885 0.325 ;
      RECT  5.255 0.05 5.425 0.33 ;
      RECT  6.3 0.05 6.47 0.33 ;
      RECT  5.8 0.05 5.92 0.37 ;
      RECT  0.07 0.05 0.21 0.39 ;
      RECT  9.0 0.05 9.14 0.39 ;
      RECT  3.47 0.05 3.59 0.41 ;
      RECT  8.495 0.05 8.615 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.77 0.14 2.51 0.23 ;
      RECT  2.42 0.23 2.51 0.295 ;
      RECT  0.77 0.23 0.89 0.405 ;
      RECT  2.42 0.295 3.38 0.415 ;
      RECT  7.96 0.14 8.19 0.24 ;
      RECT  7.96 0.24 8.05 0.285 ;
      RECT  7.275 0.285 8.05 0.375 ;
      RECT  7.275 0.375 7.635 0.38 ;
      RECT  7.545 0.38 7.635 0.98 ;
      RECT  7.345 0.98 7.635 1.095 ;
      RECT  1.03 0.32 2.24 0.44 ;
      RECT  1.03 0.44 1.15 0.71 ;
      RECT  1.03 0.71 1.76 0.8 ;
      RECT  1.67 0.8 1.76 1.025 ;
      RECT  1.67 1.025 2.86 1.04 ;
      RECT  1.965 0.95 2.86 1.025 ;
      RECT  1.67 1.04 2.055 1.115 ;
      RECT  2.77 1.04 2.86 1.21 ;
      RECT  2.77 1.21 4.1 1.3 ;
      RECT  3.98 0.29 4.1 1.21 ;
      RECT  2.77 1.3 2.86 1.47 ;
      RECT  2.685 1.47 2.86 1.585 ;
      RECT  5.54 0.23 5.66 0.46 ;
      RECT  5.54 0.46 5.99 0.55 ;
      RECT  5.9 0.55 5.99 0.68 ;
      RECT  5.9 0.68 5.995 0.77 ;
      RECT  5.905 0.77 5.995 1.015 ;
      RECT  5.905 1.015 6.73 1.125 ;
      RECT  5.905 1.125 5.995 1.24 ;
      RECT  4.41 1.145 4.5 1.24 ;
      RECT  4.41 1.24 5.995 1.345 ;
      RECT  4.41 1.345 4.5 1.57 ;
      RECT  3.375 1.57 4.5 1.66 ;
      RECT  0.34 0.19 0.46 0.485 ;
      RECT  0.15 0.485 0.46 0.575 ;
      RECT  0.15 0.575 0.25 1.29 ;
      RECT  6.08 0.42 7.005 0.51 ;
      RECT  6.08 0.51 6.185 0.615 ;
      RECT  6.915 0.51 7.005 1.285 ;
      RECT  6.34 1.285 7.005 1.375 ;
      RECT  6.835 1.375 7.005 1.39 ;
      RECT  6.34 1.375 6.46 1.435 ;
      RECT  5.75 1.435 6.46 1.525 ;
      RECT  4.59 0.42 5.25 0.53 ;
      RECT  4.59 0.53 4.68 0.65 ;
      RECT  5.16 0.53 5.25 1.04 ;
      RECT  4.96 1.04 5.785 1.13 ;
      RECT  5.675 0.95 5.785 1.04 ;
      RECT  1.275 0.53 3.055 0.62 ;
      RECT  4.205 0.23 4.345 0.77 ;
      RECT  4.205 0.77 5.07 0.88 ;
      RECT  4.205 0.88 4.295 1.39 ;
      RECT  3.6 1.39 4.295 1.48 ;
      RECT  8.445 0.785 8.835 0.895 ;
      RECT  8.445 0.895 8.535 1.315 ;
      RECT  8.275 1.315 8.535 1.405 ;
      RECT  8.275 1.405 8.365 1.42 ;
      RECT  6.9 0.22 7.185 0.33 ;
      RECT  7.095 0.33 7.185 1.42 ;
      RECT  7.095 1.42 8.365 1.48 ;
      RECT  6.575 1.465 6.745 1.48 ;
      RECT  6.575 1.48 8.365 1.51 ;
      RECT  6.575 1.51 7.185 1.57 ;
      RECT  3.73 0.245 3.85 0.95 ;
      RECT  3.73 0.95 3.86 1.0 ;
      RECT  3.45 1.0 3.86 1.12 ;
      RECT  8.21 0.39 8.33 1.135 ;
      RECT  7.735 1.135 8.33 1.2 ;
      RECT  7.42 1.2 8.33 1.225 ;
      RECT  7.42 1.225 7.825 1.295 ;
      RECT  2.495 1.15 2.675 1.38 ;
      RECT  2.495 1.38 2.595 1.6 ;
      RECT  0.595 1.39 1.33 1.43 ;
      RECT  0.08 1.43 1.33 1.48 ;
      RECT  0.08 1.48 0.67 1.52 ;
      RECT  0.08 1.52 0.2 1.625 ;
      RECT  1.42 1.39 2.125 1.495 ;
      RECT  1.42 1.495 1.53 1.57 ;
      RECT  0.84 1.57 1.53 1.66 ;
      LAYER M2 ;
      RECT  0.11 1.15 2.675 1.25 ;
      LAYER V1 ;
      RECT  0.15 1.15 0.25 1.25 ;
      RECT  2.535 1.15 2.635 1.25 ;
  END
END SEN_FSDPTQO_2
#-----------------------------------------------------------------------
#      Cell        : SEN_FSDPTQO_4
#      Description : "D-Flip Flop w/scan, pos-edge triggered, hi-sync-set, q-only, so pin"
#      Equation    : iq,iqn=ff(clocked_on=CK,next_state=((!SE&(D|SS))|(SE&SI))):Q=iq:SO=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_FSDPTQO_4
  CLASS CORE ;
  FOREIGN SEN_FSDPTQO_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN CK
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.655 0.45 7.745 0.715 ;
      RECT  7.655 0.715 7.895 0.85 ;
      RECT  6.84 0.71 7.14 0.89 ;
      RECT  5.55 0.71 5.88 0.89 ;
      LAYER M2 ;
      RECT  5.7 0.75 7.895 0.85 ;
      LAYER V1 ;
      RECT  7.755 0.75 7.855 0.85 ;
      RECT  6.84 0.75 6.94 0.85 ;
      RECT  7.04 0.75 7.14 0.85 ;
      RECT  5.74 0.75 5.84 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1182 ;
  END CK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.965 0.72 ;
      RECT  1.35 0.72 3.05 0.81 ;
      RECT  1.35 0.81 1.965 0.89 ;
      RECT  2.95 0.81 3.05 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END D
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.15 0.51 9.85 0.69 ;
      RECT  9.75 0.69 9.85 1.11 ;
      RECT  9.15 1.11 9.85 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN SE
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.195 ;
      RECT  0.35 1.195 2.375 1.285 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1035 ;
  END SE
  PIN SI
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.65 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END SI
  PIN SO
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.35 0.31 8.5 0.49 ;
      RECT  8.35 0.49 8.45 0.93 ;
      RECT  8.35 0.93 8.52 1.02 ;
    END
    ANTENNADIFFAREA 0.119 ;
  END SO
  PIN SS
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.83 ;
      RECT  0.75 0.83 0.895 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END SS
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.61 0.48 1.75 ;
      RECT  0.0 1.75 10.2 1.85 ;
      RECT  2.17 1.415 2.285 1.75 ;
      RECT  3.21 1.39 3.33 1.75 ;
      RECT  4.81 1.43 4.98 1.75 ;
      RECT  5.33 1.43 5.5 1.75 ;
      RECT  5.875 1.42 5.995 1.75 ;
      RECT  6.395 1.59 6.565 1.75 ;
      RECT  8.075 1.615 8.245 1.75 ;
      RECT  8.865 1.48 9.035 1.75 ;
      RECT  9.41 1.38 9.53 1.75 ;
      RECT  9.95 1.21 10.07 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      RECT  2.63 0.05 2.8 0.17 ;
      RECT  6.42 0.05 6.59 0.305 ;
      RECT  5.355 0.05 5.475 0.36 ;
      RECT  5.865 0.05 6.0 0.36 ;
      RECT  8.09 0.05 8.21 0.36 ;
      RECT  4.835 0.05 4.955 0.37 ;
      RECT  3.545 0.05 3.665 0.385 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  9.41 0.05 9.53 0.42 ;
      RECT  8.89 0.05 9.01 0.585 ;
      RECT  9.95 0.05 10.07 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.71 0.14 2.54 0.23 ;
      RECT  2.45 0.23 2.54 0.29 ;
      RECT  0.71 0.23 0.8 0.42 ;
      RECT  2.45 0.29 3.455 0.4 ;
      RECT  5.62 0.29 5.73 0.45 ;
      RECT  5.62 0.45 6.08 0.54 ;
      RECT  5.99 0.54 6.08 0.655 ;
      RECT  5.99 0.655 6.54 0.745 ;
      RECT  6.45 0.745 6.54 1.06 ;
      RECT  6.45 1.06 7.13 1.17 ;
      RECT  6.45 1.17 6.54 1.23 ;
      RECT  4.515 1.11 4.605 1.23 ;
      RECT  4.515 1.23 6.54 1.32 ;
      RECT  4.515 1.32 4.605 1.56 ;
      RECT  3.48 1.56 4.605 1.66 ;
      RECT  7.835 0.19 7.925 0.45 ;
      RECT  7.835 0.45 8.075 0.54 ;
      RECT  7.985 0.54 8.075 0.625 ;
      RECT  7.985 0.625 8.26 0.795 ;
      RECT  7.985 0.795 8.075 0.96 ;
      RECT  7.77 0.96 8.075 1.07 ;
      RECT  4.0 0.3 4.19 0.49 ;
      RECT  4.1 0.49 4.19 1.115 ;
      RECT  3.97 1.115 4.19 1.22 ;
      RECT  0.345 0.19 0.465 0.5 ;
      RECT  0.15 0.5 0.465 0.59 ;
      RECT  0.15 0.59 0.25 1.29 ;
      RECT  6.17 0.395 7.365 0.5 ;
      RECT  6.17 0.5 6.27 0.565 ;
      RECT  7.26 0.5 7.365 1.29 ;
      RECT  6.75 1.29 7.365 1.38 ;
      RECT  6.75 1.38 6.84 1.41 ;
      RECT  7.255 1.38 7.365 1.455 ;
      RECT  6.135 1.41 6.84 1.5 ;
      RECT  6.135 1.5 6.255 1.625 ;
      RECT  1.165 0.53 2.12 0.54 ;
      RECT  1.165 0.54 3.11 0.62 ;
      RECT  2.03 0.62 3.11 0.63 ;
      RECT  4.335 0.19 4.45 0.765 ;
      RECT  4.335 0.765 5.165 0.865 ;
      RECT  4.335 0.865 4.425 1.335 ;
      RECT  3.735 1.335 4.425 1.455 ;
      RECT  3.805 0.19 3.91 0.83 ;
      RECT  3.805 0.83 4.01 0.91 ;
      RECT  3.55 0.91 4.01 1.0 ;
      RECT  3.55 1.0 3.64 1.24 ;
      RECT  3.43 1.24 3.64 1.36 ;
      RECT  8.815 0.785 9.65 0.895 ;
      RECT  8.815 0.895 8.905 1.3 ;
      RECT  8.685 1.3 8.905 1.39 ;
      RECT  8.685 1.39 8.775 1.435 ;
      RECT  6.95 0.175 7.665 0.265 ;
      RECT  6.95 0.265 7.12 0.305 ;
      RECT  7.475 0.265 7.665 0.36 ;
      RECT  7.475 0.36 7.565 0.94 ;
      RECT  7.475 0.94 7.655 1.11 ;
      RECT  7.565 1.11 7.655 1.435 ;
      RECT  7.565 1.435 8.775 1.525 ;
      RECT  7.565 1.525 7.655 1.545 ;
      RECT  6.97 1.47 7.14 1.545 ;
      RECT  6.97 1.545 7.655 1.65 ;
      RECT  6.065 0.865 6.325 0.975 ;
      RECT  6.065 0.975 6.155 1.05 ;
      RECT  4.695 0.47 5.345 0.585 ;
      RECT  4.695 0.585 4.795 0.64 ;
      RECT  5.255 0.585 5.345 1.04 ;
      RECT  5.045 1.04 5.345 1.05 ;
      RECT  5.045 1.05 6.155 1.14 ;
      RECT  2.35 0.9 2.84 0.99 ;
      RECT  2.35 0.99 2.44 1.0 ;
      RECT  2.75 0.99 2.84 1.465 ;
      RECT  0.93 0.335 2.36 0.425 ;
      RECT  0.985 0.425 2.36 0.44 ;
      RECT  2.175 0.44 2.36 0.45 ;
      RECT  0.985 0.44 1.075 1.0 ;
      RECT  0.985 1.0 2.44 1.105 ;
      RECT  2.655 1.465 2.84 1.585 ;
      RECT  8.62 0.19 8.725 1.12 ;
      RECT  8.165 1.12 8.725 1.21 ;
      RECT  8.165 1.21 8.255 1.22 ;
      RECT  7.87 1.22 8.255 1.325 ;
      RECT  2.53 1.08 2.635 1.21 ;
      RECT  2.465 1.21 2.635 1.3 ;
      RECT  2.465 1.3 2.555 1.635 ;
      RECT  0.065 1.39 1.305 1.48 ;
      RECT  0.065 1.48 0.185 1.615 ;
      RECT  1.395 1.375 2.08 1.495 ;
      RECT  1.395 1.495 1.515 1.57 ;
      RECT  0.825 1.57 1.515 1.66 ;
      LAYER M2 ;
      RECT  2.18 0.35 4.14 0.45 ;
      RECT  0.11 1.15 2.675 1.25 ;
      LAYER V1 ;
      RECT  2.22 0.35 2.32 0.45 ;
      RECT  4.0 0.35 4.1 0.45 ;
      RECT  0.15 1.15 0.25 1.25 ;
      RECT  2.535 1.15 2.635 1.25 ;
  END
END SEN_FSDPTQO_4
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_0P5
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_0P5
  CLASS CORE ;
  FOREIGN SEN_INV_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.215 1.75 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      RECT  0.065 0.05 0.215 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.295 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.094 ;
  END X
END SEN_INV_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_1
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_1
  CLASS CORE ;
  FOREIGN SEN_INV_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      RECT  0.08 0.05 0.2 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
END SEN_INV_1
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_2
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_2
  CLASS CORE ;
  FOREIGN SEN_INV_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.6 1.21 0.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.08 0.05 0.2 0.39 ;
      RECT  0.6 0.05 0.72 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
END SEN_INV_2
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_3
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_3
  CLASS CORE ;
  FOREIGN SEN_INV_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.74 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.14 1.24 0.255 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.67 1.4 0.79 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.67 0.05 0.79 0.36 ;
      RECT  0.14 0.05 0.255 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.38 0.45 1.05 0.57 ;
      RECT  0.95 0.57 1.05 1.11 ;
      RECT  0.35 1.11 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
END SEN_INV_3
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_4
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_4
  CLASS CORE ;
  FOREIGN SEN_INV_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.75 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.14 1.21 0.245 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.66 1.41 0.78 1.75 ;
      RECT  1.195 1.21 1.315 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.65 0.05 0.79 0.37 ;
      RECT  0.14 0.05 0.25 0.59 ;
      RECT  1.195 0.05 1.315 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.375 0.46 1.05 0.58 ;
      RECT  0.93 0.58 1.05 1.11 ;
      RECT  0.35 1.11 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
END SEN_INV_4
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_6
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_6
  CLASS CORE ;
  FOREIGN SEN_INV_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.26 0.895 ;
      RECT  0.15 0.895 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.57 1.415 0.705 1.75 ;
      RECT  1.105 1.41 1.225 1.75 ;
      RECT  1.625 1.41 1.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.57 0.05 0.715 0.385 ;
      RECT  1.09 0.05 1.235 0.385 ;
      RECT  1.625 0.05 1.745 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.3 0.5 1.48 0.62 ;
      RECT  1.35 0.62 1.48 1.11 ;
      RECT  0.34 1.11 1.48 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
END SEN_INV_6
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_8
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_8
  CLASS CORE ;
  FOREIGN SEN_INV_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.705 1.59 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.095 1.21 0.215 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.645 1.44 0.765 1.75 ;
      RECT  1.165 1.44 1.285 1.75 ;
      RECT  1.685 1.44 1.805 1.75 ;
      RECT  2.215 1.21 2.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.635 0.05 0.775 0.37 ;
      RECT  1.155 0.05 1.29 0.37 ;
      RECT  1.675 0.05 1.81 0.37 ;
      RECT  0.095 0.05 0.215 0.59 ;
      RECT  2.215 0.05 2.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.36 0.465 2.09 0.595 ;
      RECT  1.68 0.595 1.85 1.11 ;
      RECT  0.35 1.11 2.065 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
END SEN_INV_8
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_0P5
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_0P5
  CLASS CORE ;
  FOREIGN SEN_INV_AS_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.085 0.25 0.205 0.51 ;
      RECT  0.085 0.51 0.45 0.69 ;
      RECT  0.35 0.69 0.45 1.09 ;
    END
    ANTENNADIFFAREA 0.077 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.415 0.455 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.335 0.05 0.455 0.405 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.21 0.735 0.385 ;
      RECT  0.55 0.385 0.65 1.31 ;
      RECT  0.55 1.31 0.735 1.49 ;
    END
    ANTENNADIFFAREA 0.076 ;
  END X
END SEN_INV_AS_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_1
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_1
  CLASS CORE ;
  FOREIGN SEN_INV_AS_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.095 0.205 0.25 1.095 ;
    END
    ANTENNADIFFAREA 0.096 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0549 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.28 1.21 0.4 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.61 0.05 0.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.28 0.475 0.51 ;
      RECT  0.35 0.51 0.67 0.69 ;
      RECT  0.54 0.69 0.67 1.5 ;
    END
    ANTENNADIFFAREA 0.146 ;
  END X
END SEN_INV_AS_1
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_10
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_10
  CLASS CORE ;
  FOREIGN SEN_INV_AS_10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.285 0.25 0.71 ;
      RECT  0.15 0.71 1.465 0.89 ;
    END
    ANTENNADIFFAREA 0.084 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5616 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.59 1.415 0.71 1.75 ;
      RECT  1.11 1.415 1.23 1.75 ;
      RECT  1.63 1.415 1.75 1.75 ;
      RECT  2.15 1.4 2.27 1.75 ;
      RECT  2.69 1.21 2.81 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  1.11 0.05 1.23 0.35 ;
      RECT  1.63 0.05 1.75 0.35 ;
      RECT  2.15 0.05 2.27 0.385 ;
      RECT  0.56 0.05 0.68 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.8 0.44 1.85 0.51 ;
      RECT  0.8 0.51 2.65 0.56 ;
      RECT  1.63 0.56 2.65 0.69 ;
      RECT  1.63 0.69 1.85 1.11 ;
      RECT  0.325 1.11 2.53 1.29 ;
    END
    ANTENNADIFFAREA 0.965 ;
  END X
END SEN_INV_AS_10
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_12
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_12
  CLASS CORE ;
  FOREIGN SEN_INV_AS_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.17 0.25 0.71 ;
      RECT  0.15 0.71 2.155 0.89 ;
      RECT  0.15 0.89 0.25 1.29 ;
    END
    ANTENNADIFFAREA 0.095 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6576 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.13 1.41 0.26 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.63 1.46 0.8 1.75 ;
      RECT  1.15 1.46 1.32 1.75 ;
      RECT  1.67 1.46 1.84 1.75 ;
      RECT  2.19 1.455 2.36 1.75 ;
      RECT  2.71 1.455 2.88 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.63 0.05 0.8 0.33 ;
      RECT  1.15 0.05 1.32 0.33 ;
      RECT  1.67 0.05 1.84 0.33 ;
      RECT  2.19 0.05 2.36 0.33 ;
      RECT  2.71 0.05 2.88 0.33 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.42 3.115 0.605 ;
      RECT  2.35 0.605 3.115 0.69 ;
      RECT  2.35 0.69 2.65 1.11 ;
      RECT  0.35 1.11 3.115 1.335 ;
    END
    ANTENNADIFFAREA 1.187 ;
  END X
END SEN_INV_AS_12
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_16
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_16
  CLASS CORE ;
  FOREIGN SEN_INV_AS_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.205 0.25 0.71 ;
      RECT  0.15 0.71 2.145 0.89 ;
    END
    ANTENNADIFFAREA 0.105 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8796 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.345 1.445 0.515 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.865 1.445 1.035 1.75 ;
      RECT  1.385 1.445 1.555 1.75 ;
      RECT  1.905 1.445 2.075 1.75 ;
      RECT  2.425 1.445 2.595 1.75 ;
      RECT  2.945 1.445 3.115 1.75 ;
      RECT  3.465 1.445 3.635 1.75 ;
      RECT  4.005 1.41 4.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.865 0.05 1.035 0.31 ;
      RECT  1.385 0.05 1.555 0.31 ;
      RECT  1.905 0.05 2.075 0.31 ;
      RECT  2.425 0.05 2.595 0.31 ;
      RECT  2.945 0.05 3.115 0.31 ;
      RECT  3.465 0.05 3.635 0.31 ;
      RECT  0.365 0.05 0.495 0.385 ;
      RECT  4.005 0.05 4.135 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.62 0.405 3.915 0.6 ;
      RECT  2.35 0.6 3.915 0.695 ;
      RECT  2.35 0.695 2.65 1.085 ;
      RECT  0.11 1.085 3.905 1.325 ;
    END
    ANTENNADIFFAREA 1.512 ;
  END X
END SEN_INV_AS_16
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_1P5
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_1P5
  CLASS CORE ;
  FOREIGN SEN_INV_AS_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.255 0.185 0.51 ;
      RECT  0.065 0.51 0.455 0.69 ;
      RECT  0.345 0.69 0.455 0.94 ;
    END
    ANTENNADIFFAREA 0.058 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.24 1.21 0.36 1.75 ;
      RECT  0.0 1.75 1.0 1.85 ;
      RECT  0.815 1.21 0.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      RECT  0.805 0.05 0.94 0.39 ;
      RECT  0.295 0.05 0.415 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.21 0.66 1.49 ;
    END
    ANTENNADIFFAREA 0.138 ;
  END X
END SEN_INV_AS_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_2
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_2
  CLASS CORE ;
  FOREIGN SEN_INV_AS_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.495 0.25 1.1 ;
    END
    ANTENNADIFFAREA 0.063 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1098 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.275 1.41 0.405 1.75 ;
      RECT  0.0 1.75 1.0 1.85 ;
      RECT  0.795 1.41 0.925 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      RECT  0.25 0.05 0.375 0.39 ;
      RECT  0.795 0.05 0.925 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 1.5 ;
    END
    ANTENNADIFFAREA 0.214 ;
  END X
END SEN_INV_AS_2
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_3
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_3
  CLASS CORE ;
  FOREIGN SEN_INV_AS_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.125 0.215 0.25 1.1 ;
    END
    ANTENNADIFFAREA 0.108 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1644 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.155 1.41 0.285 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.68 1.21 0.8 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.94 0.05 1.065 0.39 ;
      RECT  0.41 0.05 0.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.69 0.31 0.85 0.91 ;
      RECT  0.42 0.91 1.05 1.09 ;
      RECT  0.42 1.09 0.54 1.22 ;
      RECT  0.95 1.09 1.05 1.295 ;
    END
    ANTENNADIFFAREA 0.313 ;
  END X
END SEN_INV_AS_3
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_4
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_4
  CLASS CORE ;
  FOREIGN SEN_INV_AS_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.135 0.205 0.25 0.3 ;
      RECT  0.135 0.3 0.26 0.71 ;
      RECT  0.135 0.71 0.685 0.89 ;
      RECT  0.135 0.89 0.25 1.09 ;
    END
    ANTENNADIFFAREA 0.108 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.105 1.41 0.235 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.635 1.41 0.765 1.75 ;
      RECT  1.165 1.41 1.295 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.895 0.05 1.025 0.39 ;
      RECT  0.38 0.05 0.5 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.3 1.28 0.48 ;
      RECT  0.615 0.48 1.28 0.59 ;
      RECT  1.15 0.59 1.28 1.11 ;
      RECT  0.345 1.11 1.28 1.29 ;
    END
    ANTENNADIFFAREA 0.391 ;
  END X
END SEN_INV_AS_4
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_5
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_5
  CLASS CORE ;
  FOREIGN SEN_INV_AS_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.09 0.235 0.25 0.71 ;
      RECT  0.09 0.71 1.05 0.79 ;
      RECT  0.15 0.79 1.05 0.89 ;
      RECT  0.15 0.89 0.25 1.14 ;
    END
    ANTENNADIFFAREA 0.084 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2796 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.09 1.23 0.21 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.63 1.38 0.75 1.75 ;
      RECT  1.15 1.38 1.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.63 0.05 0.75 0.35 ;
      RECT  1.15 0.05 1.27 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.41 0.325 1.53 0.44 ;
      RECT  0.34 0.44 1.53 0.56 ;
      RECT  1.14 0.56 1.25 1.11 ;
      RECT  0.35 1.11 1.53 1.29 ;
    END
    ANTENNADIFFAREA 0.55 ;
  END X
END SEN_INV_AS_5
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_6
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_6
  CLASS CORE ;
  FOREIGN SEN_INV_AS_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.14 0.21 0.25 0.71 ;
      RECT  0.14 0.71 0.89 0.89 ;
      RECT  0.14 0.89 0.25 1.1 ;
    END
    ANTENNADIFFAREA 0.12 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3288 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.18 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.57 1.41 0.695 1.75 ;
      RECT  1.09 1.41 1.22 1.75 ;
      RECT  1.61 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.03 0.05 1.16 0.39 ;
      RECT  1.565 0.05 1.695 0.39 ;
      RECT  0.495 0.05 0.615 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.485 1.47 0.595 ;
      RECT  1.35 0.595 1.47 1.11 ;
      RECT  0.55 1.11 1.47 1.205 ;
      RECT  0.32 1.205 1.47 1.295 ;
      RECT  0.32 1.295 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.548 ;
  END X
END SEN_INV_AS_6
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_AS_8
#      Description : "Symmetric rise/fall time inverter, antenna diode on input"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_AS_8
  CLASS CORE ;
  FOREIGN SEN_INV_AS_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.205 0.25 0.71 ;
      RECT  0.15 0.71 1.555 0.89 ;
      RECT  0.15 0.89 0.25 1.125 ;
    END
    ANTENNADIFFAREA 0.12 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4392 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.105 1.41 0.235 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.635 1.41 0.765 1.75 ;
      RECT  1.155 1.41 1.285 1.75 ;
      RECT  1.675 1.41 1.805 1.75 ;
      RECT  2.195 1.41 2.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.155 0.05 1.285 0.345 ;
      RECT  1.675 0.05 1.805 0.345 ;
      RECT  2.195 0.05 2.325 0.39 ;
      RECT  0.6 0.05 0.72 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.865 0.45 2.05 0.62 ;
      RECT  1.75 0.62 2.05 1.11 ;
      RECT  0.35 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.732 ;
  END X
END SEN_INV_AS_8
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_0P5
#      Description : "Symmetric rise/fall time inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_0P5
  CLASS CORE ;
  FOREIGN SEN_INV_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      RECT  0.065 0.05 0.205 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.195 0.45 1.53 ;
    END
    ANTENNADIFFAREA 0.085 ;
  END X
END SEN_INV_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_1P5
#      Description : "Symmetric rise/fall time inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_1P5
  CLASS CORE ;
  FOREIGN SEN_INV_S_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.6 1.21 0.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.065 0.05 0.205 0.39 ;
      RECT  0.59 0.05 0.73 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.2 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.142 ;
  END X
END SEN_INV_S_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_32
#      Description : "Symmetric rise/fall time inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_32
  CLASS CORE ;
  FOREIGN SEN_INV_S_32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.695 4.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.7937 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.57 1.455 0.74 1.75 ;
      RECT  1.09 1.455 1.26 1.75 ;
      RECT  1.61 1.455 1.78 1.75 ;
      RECT  2.13 1.455 2.3 1.75 ;
      RECT  2.65 1.455 2.82 1.75 ;
      RECT  3.17 1.455 3.34 1.75 ;
      RECT  3.69 1.455 3.86 1.75 ;
      RECT  4.21 1.455 4.38 1.75 ;
      RECT  4.73 1.455 4.9 1.75 ;
      RECT  5.25 1.455 5.42 1.75 ;
      RECT  5.77 1.455 5.94 1.75 ;
      RECT  6.29 1.455 6.46 1.75 ;
      RECT  6.81 1.455 6.98 1.75 ;
      RECT  7.33 1.455 7.5 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  0.57 0.05 0.74 0.305 ;
      RECT  1.09 0.05 1.26 0.305 ;
      RECT  1.61 0.05 1.78 0.305 ;
      RECT  2.13 0.05 2.3 0.305 ;
      RECT  2.65 0.05 2.82 0.305 ;
      RECT  3.17 0.05 3.34 0.305 ;
      RECT  3.69 0.05 3.86 0.305 ;
      RECT  4.21 0.05 4.38 0.305 ;
      RECT  4.73 0.05 4.9 0.305 ;
      RECT  5.25 0.05 5.42 0.305 ;
      RECT  5.77 0.05 5.94 0.305 ;
      RECT  6.29 0.05 6.46 0.305 ;
      RECT  6.81 0.05 6.98 0.305 ;
      RECT  7.33 0.05 7.5 0.305 ;
      RECT  0.075 0.05 0.195 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.6 0.325 7.735 0.405 ;
      RECT  0.285 0.405 7.735 0.525 ;
      RECT  1.9 0.525 7.735 0.57 ;
      RECT  1.9 0.57 6.25 0.595 ;
      RECT  4.75 0.595 6.25 0.755 ;
      RECT  5.65 0.755 6.25 1.005 ;
      RECT  4.75 1.005 6.25 1.11 ;
      RECT  1.95 1.11 7.73 1.21 ;
      RECT  0.285 1.21 7.73 1.33 ;
    END
    ANTENNADIFFAREA 3.048 ;
  END X
END SEN_INV_S_32
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_1
#      Description : "Symmetric rise/fall delay inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_1
  CLASS CORE ;
  FOREIGN SEN_INV_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0549 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      RECT  0.075 0.05 0.205 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.31 0.46 1.29 ;
    END
    ANTENNADIFFAREA 0.174 ;
  END X
END SEN_INV_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_12
#      Description : "Symmetric rise/fall delay inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_12
  CLASS CORE ;
  FOREIGN SEN_INV_S_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.685 2.65 0.89 ;
      RECT  0.55 0.685 1.45 0.89 ;
      LAYER M2 ;
      RECT  1.31 0.75 2.09 0.85 ;
      LAYER V1 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6576 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      RECT  1.115 1.41 1.245 1.75 ;
      RECT  1.635 1.41 1.765 1.75 ;
      RECT  2.155 1.41 2.285 1.75 ;
      RECT  2.675 1.41 2.805 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  1.635 0.05 1.765 0.365 ;
      RECT  0.595 0.05 0.725 0.39 ;
      RECT  1.115 0.05 1.245 0.39 ;
      RECT  2.155 0.05 2.285 0.39 ;
      RECT  2.675 0.05 2.805 0.39 ;
      RECT  0.08 0.05 0.2 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.5 0.455 ;
      RECT  1.35 0.455 2.05 0.485 ;
      RECT  1.9 0.31 2.05 0.455 ;
      RECT  0.34 0.31 0.46 0.485 ;
      RECT  0.34 0.485 3.06 0.575 ;
      RECT  0.86 0.33 0.98 0.485 ;
      RECT  2.42 0.33 2.54 0.485 ;
      RECT  2.945 0.31 3.06 0.485 ;
      RECT  1.55 0.575 1.85 1.11 ;
      RECT  0.34 1.11 3.06 1.29 ;
    END
    ANTENNADIFFAREA 1.17 ;
  END X
END SEN_INV_S_12
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_16
#      Description : "Symmetric rise/fall delay inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_16
  CLASS CORE ;
  FOREIGN SEN_INV_S_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.685 3.25 0.89 ;
      RECT  0.55 0.685 1.65 0.89 ;
      LAYER M2 ;
      RECT  1.51 0.75 2.29 0.85 ;
      LAYER V1 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8796 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.09 1.21 0.21 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.615 1.41 0.745 1.75 ;
      RECT  1.135 1.41 1.265 1.75 ;
      RECT  1.655 1.41 1.785 1.75 ;
      RECT  2.175 1.41 2.305 1.75 ;
      RECT  2.695 1.41 2.825 1.75 ;
      RECT  3.215 1.41 3.345 1.75 ;
      RECT  3.76 1.21 3.88 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.615 0.05 0.745 0.345 ;
      RECT  1.135 0.05 1.265 0.345 ;
      RECT  1.655 0.05 1.785 0.345 ;
      RECT  2.175 0.05 2.305 0.345 ;
      RECT  2.695 0.05 2.825 0.345 ;
      RECT  3.215 0.05 3.345 0.345 ;
      RECT  0.08 0.05 0.2 0.59 ;
      RECT  3.76 0.05 3.88 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.48 0.435 ;
      RECT  0.35 0.435 3.65 0.575 ;
      RECT  3.55 0.31 3.65 0.435 ;
      RECT  1.74 0.575 2.06 1.11 ;
      RECT  0.35 1.11 3.65 1.29 ;
    END
    ANTENNADIFFAREA 1.47 ;
  END X
END SEN_INV_S_16
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_2
#      Description : "Symmetric rise/fall delay inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_2
  CLASS CORE ;
  FOREIGN SEN_INV_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1098 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.6 1.21 0.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.205 0.39 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.31 0.46 1.29 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
END SEN_INV_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_3
#      Description : "Symmetric rise/fall time inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_3
  CLASS CORE ;
  FOREIGN SEN_INV_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1644 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.12 1.21 0.24 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.665 1.415 0.795 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.84 0.05 0.96 0.385 ;
      RECT  0.24 0.05 0.36 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.3 0.65 0.485 ;
      RECT  0.55 0.485 1.06 0.605 ;
      RECT  0.94 0.605 1.06 1.205 ;
      RECT  0.38 1.205 1.06 1.325 ;
    END
    ANTENNADIFFAREA 0.314 ;
  END X
END SEN_INV_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_4
#      Description : "Symmetric rise/fall delay inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_4
  CLASS CORE ;
  FOREIGN SEN_INV_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2196 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.1 1.21 0.22 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.635 1.415 0.765 1.75 ;
      RECT  1.18 1.21 1.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.635 0.05 0.765 0.385 ;
      RECT  1.17 0.05 1.29 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.355 0.475 1.05 0.595 ;
      RECT  0.95 0.595 1.05 1.205 ;
      RECT  0.35 1.205 1.05 1.325 ;
    END
    ANTENNADIFFAREA 0.391 ;
  END X
END SEN_INV_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_6
#      Description : "Symmetric rise/fall time inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_6
  CLASS CORE ;
  FOREIGN SEN_INV_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.04 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3288 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  0.3 0.05 0.42 0.59 ;
      RECT  1.44 0.05 1.56 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.56 0.5 1.26 0.62 ;
      RECT  1.13 0.62 1.26 1.11 ;
      RECT  0.34 1.11 1.65 1.29 ;
    END
    ANTENNADIFFAREA 0.548 ;
  END X
END SEN_INV_S_6
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_S_8
#      Description : "Symmetric rise/fall delay inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_S_8
  CLASS CORE ;
  FOREIGN SEN_INV_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.685 1.67 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4392 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.09 1.21 0.21 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  0.63 1.41 0.76 1.75 ;
      RECT  1.165 1.41 1.295 1.75 ;
      RECT  1.685 1.41 1.815 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  1.165 0.05 1.295 0.355 ;
      RECT  1.685 0.05 1.815 0.355 ;
      RECT  0.63 0.05 0.76 0.385 ;
      RECT  0.08 0.05 0.2 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.91 0.31 1.05 0.445 ;
      RECT  0.91 0.445 2.06 0.485 ;
      RECT  1.95 0.31 2.06 0.445 ;
      RECT  0.35 0.31 0.48 0.485 ;
      RECT  0.35 0.485 2.06 0.575 ;
      RECT  1.89 0.575 2.06 1.11 ;
      RECT  0.35 1.11 2.06 1.29 ;
    END
    ANTENNADIFFAREA 0.817 ;
  END X
END SEN_INV_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_0P65
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_0P65
  CLASS CORE ;
  FOREIGN SEN_INV_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0423 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      RECT  0.065 0.05 0.205 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.28 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.116 ;
  END X
END SEN_INV_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_0P8
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_0P8
  CLASS CORE ;
  FOREIGN SEN_INV_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      RECT  0.065 0.05 0.205 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 1.35 ;
    END
    ANTENNADIFFAREA 0.143 ;
  END X
END SEN_INV_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_10
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_10
  CLASS CORE ;
  FOREIGN SEN_INV_10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.7 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.595 1.42 0.715 1.75 ;
      RECT  1.115 1.42 1.235 1.75 ;
      RECT  1.635 1.42 1.755 1.75 ;
      RECT  2.155 1.42 2.275 1.75 ;
      RECT  2.71 1.21 2.83 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  0.57 0.05 0.74 0.335 ;
      RECT  1.09 0.05 1.26 0.335 ;
      RECT  1.61 0.05 1.78 0.335 ;
      RECT  2.13 0.05 2.3 0.335 ;
      RECT  0.075 0.05 0.195 0.59 ;
      RECT  2.71 0.05 2.83 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.285 0.435 2.585 0.555 ;
      RECT  0.285 0.555 2.05 0.565 ;
      RECT  1.8 0.565 2.05 1.11 ;
      RECT  1.35 1.11 2.05 1.21 ;
      RECT  0.285 1.21 2.585 1.33 ;
    END
    ANTENNADIFFAREA 1.08 ;
  END X
END SEN_INV_10
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_12
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_12
  CLASS CORE ;
  FOREIGN SEN_INV_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 2.3 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.595 1.44 0.715 1.75 ;
      RECT  1.115 1.44 1.235 1.75 ;
      RECT  1.635 1.44 1.755 1.75 ;
      RECT  2.155 1.44 2.275 1.75 ;
      RECT  2.675 1.44 2.795 1.75 ;
      RECT  3.2 1.21 3.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.57 0.05 0.74 0.325 ;
      RECT  1.09 0.05 1.26 0.325 ;
      RECT  1.61 0.05 1.78 0.325 ;
      RECT  2.13 0.05 2.3 0.325 ;
      RECT  2.65 0.05 2.82 0.325 ;
      RECT  0.075 0.05 0.195 0.59 ;
      RECT  3.2 0.05 3.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.285 0.415 3.105 0.535 ;
      RECT  1.35 0.535 2.65 0.585 ;
      RECT  2.4 0.585 2.65 1.11 ;
      RECT  1.35 1.11 2.65 1.23 ;
      RECT  0.285 1.23 3.105 1.35 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
END SEN_INV_12
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_16
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_16
  CLASS CORE ;
  FOREIGN SEN_INV_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 2.745 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.195 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.58 1.44 0.7 1.75 ;
      RECT  1.1 1.44 1.22 1.75 ;
      RECT  1.62 1.44 1.74 1.75 ;
      RECT  2.14 1.44 2.26 1.75 ;
      RECT  2.66 1.44 2.78 1.75 ;
      RECT  3.18 1.44 3.3 1.75 ;
      RECT  3.7 1.44 3.82 1.75 ;
      RECT  4.22 1.41 4.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.555 0.05 0.725 0.325 ;
      RECT  1.075 0.05 1.245 0.325 ;
      RECT  1.595 0.05 1.765 0.325 ;
      RECT  2.115 0.05 2.285 0.325 ;
      RECT  2.635 0.05 2.805 0.325 ;
      RECT  3.155 0.05 3.325 0.325 ;
      RECT  3.675 0.05 3.845 0.325 ;
      RECT  0.06 0.05 0.18 0.39 ;
      RECT  4.22 0.05 4.34 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.295 0.415 4.12 0.535 ;
      RECT  1.35 0.535 4.12 0.585 ;
      RECT  2.885 0.585 4.12 0.69 ;
      RECT  3.55 0.69 3.87 1.05 ;
      RECT  2.885 1.05 3.87 1.11 ;
      RECT  1.35 1.11 4.12 1.23 ;
      RECT  0.295 1.23 4.12 1.35 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
END SEN_INV_16
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_1P25
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_1P25
  CLASS CORE ;
  FOREIGN SEN_INV_1P25 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.7 ;
      RECT  0.15 0.7 0.455 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.585 1.41 0.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.065 0.05 0.205 0.39 ;
      RECT  0.585 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.345 0.27 0.45 0.49 ;
      RECT  0.345 0.49 0.65 0.59 ;
      RECT  0.55 0.59 0.65 1.21 ;
      RECT  0.345 1.21 0.65 1.31 ;
      RECT  0.345 1.31 0.45 1.5 ;
    END
    ANTENNADIFFAREA 0.136 ;
  END X
END SEN_INV_1P25
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_1P5
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_1P5
  CLASS CORE ;
  FOREIGN SEN_INV_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.455 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.6 1.21 0.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.59 0.05 0.73 0.39 ;
      RECT  0.08 0.05 0.2 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.49 ;
      RECT  0.35 0.49 0.65 0.59 ;
      RECT  0.55 0.59 0.65 1.02 ;
      RECT  0.35 1.02 0.65 1.12 ;
      RECT  0.35 1.12 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
END SEN_INV_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_20
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_20
  CLASS CORE ;
  FOREIGN SEN_INV_20 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 2.88 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.296 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.57 1.455 0.74 1.75 ;
      RECT  1.09 1.455 1.26 1.75 ;
      RECT  1.61 1.455 1.78 1.75 ;
      RECT  2.13 1.455 2.3 1.75 ;
      RECT  2.65 1.455 2.82 1.75 ;
      RECT  3.17 1.455 3.34 1.75 ;
      RECT  3.69 1.455 3.86 1.75 ;
      RECT  4.21 1.455 4.38 1.75 ;
      RECT  4.73 1.455 4.9 1.75 ;
      RECT  5.31 1.21 5.43 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.57 0.05 0.74 0.305 ;
      RECT  1.09 0.05 1.26 0.305 ;
      RECT  1.61 0.05 1.78 0.305 ;
      RECT  2.13 0.05 2.3 0.305 ;
      RECT  2.65 0.05 2.82 0.305 ;
      RECT  3.17 0.05 3.34 0.305 ;
      RECT  3.69 0.05 3.86 0.305 ;
      RECT  4.21 0.05 4.38 0.305 ;
      RECT  4.73 0.05 4.9 0.305 ;
      RECT  0.075 0.05 0.195 0.59 ;
      RECT  5.31 0.05 5.43 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.31 0.405 5.16 0.525 ;
      RECT  1.9 0.525 5.16 0.57 ;
      RECT  1.9 0.57 3.45 0.605 ;
      RECT  3.06 0.605 3.45 1.11 ;
      RECT  1.95 1.11 5.16 1.21 ;
      RECT  0.31 1.21 5.16 1.33 ;
    END
    ANTENNADIFFAREA 2.16 ;
  END X
END SEN_INV_20
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_24
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_24
  CLASS CORE ;
  FOREIGN SEN_INV_24 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 3.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5552 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.57 1.425 0.74 1.75 ;
      RECT  1.09 1.425 1.26 1.75 ;
      RECT  1.61 1.425 1.78 1.75 ;
      RECT  2.13 1.425 2.3 1.75 ;
      RECT  2.65 1.425 2.82 1.75 ;
      RECT  3.17 1.425 3.34 1.75 ;
      RECT  3.69 1.425 3.86 1.75 ;
      RECT  4.21 1.425 4.38 1.75 ;
      RECT  4.73 1.425 4.9 1.75 ;
      RECT  5.25 1.425 5.42 1.75 ;
      RECT  5.77 1.425 5.94 1.75 ;
      RECT  6.34 1.21 6.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.57 0.05 0.74 0.305 ;
      RECT  1.09 0.05 1.26 0.305 ;
      RECT  1.61 0.05 1.78 0.305 ;
      RECT  2.13 0.05 2.3 0.305 ;
      RECT  2.65 0.05 2.82 0.305 ;
      RECT  3.17 0.05 3.34 0.305 ;
      RECT  3.69 0.05 3.86 0.305 ;
      RECT  4.21 0.05 4.38 0.305 ;
      RECT  4.73 0.05 4.9 0.305 ;
      RECT  5.25 0.05 5.42 0.305 ;
      RECT  5.77 0.05 5.94 0.305 ;
      RECT  0.075 0.05 0.195 0.59 ;
      RECT  6.34 0.05 6.46 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.285 0.405 6.2 0.525 ;
      RECT  1.9 0.525 6.2 0.57 ;
      RECT  1.9 0.57 5.85 0.605 ;
      RECT  3.95 0.605 5.85 0.725 ;
      RECT  5.35 0.725 5.85 1.01 ;
      RECT  3.945 1.01 5.85 1.11 ;
      RECT  1.95 1.11 6.2 1.21 ;
      RECT  0.285 1.21 6.2 1.33 ;
    END
    ANTENNADIFFAREA 2.592 ;
  END X
END SEN_INV_24
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_2P5
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_2P5
  CLASS CORE ;
  FOREIGN SEN_INV_2P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.85 0.9 ;
      RECT  0.35 0.9 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.1 1.21 0.22 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.65 1.41 0.79 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.65 0.05 0.79 0.355 ;
      RECT  0.1 0.05 0.22 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.33 0.445 1.05 0.545 ;
      RECT  0.95 0.545 1.05 1.21 ;
      RECT  0.33 1.21 1.05 1.31 ;
    END
    ANTENNADIFFAREA 0.337 ;
  END X
END SEN_INV_2P5
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_32
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_32
  CLASS CORE ;
  FOREIGN SEN_INV_32 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 4.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.0736 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.57 1.455 0.74 1.75 ;
      RECT  1.09 1.455 1.26 1.75 ;
      RECT  1.61 1.455 1.78 1.75 ;
      RECT  2.13 1.455 2.3 1.75 ;
      RECT  2.65 1.455 2.82 1.75 ;
      RECT  3.17 1.455 3.34 1.75 ;
      RECT  3.69 1.455 3.86 1.75 ;
      RECT  4.21 1.455 4.38 1.75 ;
      RECT  4.73 1.455 4.9 1.75 ;
      RECT  5.25 1.455 5.42 1.75 ;
      RECT  5.77 1.455 5.94 1.75 ;
      RECT  6.29 1.455 6.46 1.75 ;
      RECT  6.81 1.455 6.98 1.75 ;
      RECT  7.33 1.455 7.5 1.75 ;
      RECT  7.85 1.455 8.02 1.75 ;
      RECT  8.41 1.21 8.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  0.57 0.05 0.74 0.305 ;
      RECT  1.09 0.05 1.26 0.305 ;
      RECT  1.61 0.05 1.78 0.305 ;
      RECT  2.13 0.05 2.3 0.305 ;
      RECT  2.65 0.05 2.82 0.305 ;
      RECT  3.17 0.05 3.34 0.305 ;
      RECT  3.69 0.05 3.86 0.305 ;
      RECT  4.21 0.05 4.38 0.305 ;
      RECT  4.73 0.05 4.9 0.305 ;
      RECT  5.25 0.05 5.42 0.305 ;
      RECT  5.77 0.05 5.94 0.305 ;
      RECT  6.29 0.05 6.46 0.305 ;
      RECT  6.81 0.05 6.98 0.305 ;
      RECT  7.33 0.05 7.5 0.305 ;
      RECT  7.85 0.05 8.02 0.305 ;
      RECT  0.075 0.05 0.195 0.59 ;
      RECT  8.41 0.05 8.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.31 0.405 8.28 0.525 ;
      RECT  1.9 0.525 8.28 0.585 ;
      RECT  1.9 0.585 7.255 0.6 ;
      RECT  4.95 0.6 7.255 0.735 ;
      RECT  6.605 0.735 7.255 1.005 ;
      RECT  4.945 1.005 7.255 1.07 ;
      RECT  1.95 1.07 7.255 1.095 ;
      RECT  1.95 1.095 8.28 1.21 ;
      RECT  0.31 1.21 8.28 1.33 ;
    END
    ANTENNADIFFAREA 3.456 ;
  END X
END SEN_INV_32
#-----------------------------------------------------------------------
#      Cell        : SEN_INV_5
#      Description : "Inverter"
#      Equation    : X=!A
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_INV_5
  CLASS CORE ;
  FOREIGN SEN_INV_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.59 1.395 0.72 1.75 ;
      RECT  1.11 1.395 1.24 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.59 0.05 0.72 0.385 ;
      RECT  1.11 0.05 1.24 0.385 ;
      RECT  0.075 0.05 0.195 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.3 1.49 0.49 ;
      RECT  0.285 0.49 1.49 0.59 ;
      RECT  1.15 0.59 1.25 1.205 ;
      RECT  0.285 1.205 1.49 1.305 ;
      RECT  1.35 1.305 1.49 1.5 ;
    END
    ANTENNADIFFAREA 0.61 ;
  END X
END SEN_INV_5
#-----------------------------------------------------------------------
#      Cell        : SEN_LDNQ_D_1
#      Description : "D-latch, neg-gate, q-only"
#      Equation    : iq,iqn=latch(enable=!G,data_in=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDNQ_D_1
  CLASS CORE ;
  FOREIGN SEN_LDNQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.3 0.65 0.72 ;
      RECT  0.46 0.72 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0438 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.925 0.4 1.02 0.48 ;
      RECT  0.75 0.48 1.02 0.57 ;
      RECT  0.75 0.57 0.85 1.005 ;
      RECT  0.23 0.92 0.33 1.005 ;
      RECT  0.23 1.005 0.85 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.485 1.945 0.665 ;
      RECT  1.75 0.665 1.85 0.99 ;
      RECT  1.75 0.99 1.945 1.16 ;
    END
    ANTENNADIFFAREA 0.158 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.445 0.45 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.245 1.315 1.375 1.75 ;
      RECT  1.565 1.23 1.685 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.29 0.05 1.41 0.36 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  1.56 0.05 1.69 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.76 0.205 1.2 0.31 ;
      RECT  1.11 0.31 1.2 0.71 ;
      RECT  0.94 0.71 1.46 0.8 ;
      RECT  1.36 0.8 1.46 0.925 ;
      RECT  0.94 0.8 1.03 1.36 ;
      RECT  0.76 1.36 1.03 1.47 ;
      RECT  0.045 0.19 0.185 0.36 ;
      RECT  0.045 0.36 0.135 1.25 ;
      RECT  0.045 1.25 0.66 1.35 ;
      RECT  0.56 1.35 0.66 1.56 ;
      RECT  0.045 1.35 0.185 1.62 ;
      RECT  0.56 1.56 1.09 1.66 ;
      RECT  1.295 0.45 1.415 0.53 ;
      RECT  1.295 0.53 1.64 0.62 ;
      RECT  1.55 0.62 1.64 1.045 ;
      RECT  1.13 0.89 1.23 1.045 ;
      RECT  1.13 1.045 1.64 1.135 ;
      RECT  1.295 1.135 1.415 1.225 ;
  END
END SEN_LDNQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_LDNQ_D_2
#      Description : "D-latch, neg-gate, q-only"
#      Equation    : iq,iqn=latch(enable=!G,data_in=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDNQ_D_2
  CLASS CORE ;
  FOREIGN SEN_LDNQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.3 0.65 0.665 ;
      RECT  0.46 0.665 0.65 0.76 ;
      RECT  0.46 0.76 0.56 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.925 0.4 1.02 0.48 ;
      RECT  0.75 0.48 1.02 0.57 ;
      RECT  0.75 0.57 0.85 0.875 ;
      RECT  0.685 0.875 0.85 1.005 ;
      RECT  0.23 0.825 0.33 1.005 ;
      RECT  0.23 1.005 0.85 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0615 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.3 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.244 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.445 0.45 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.245 1.315 1.375 1.75 ;
      RECT  1.615 1.23 1.735 1.75 ;
      RECT  2.21 1.21 2.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.29 0.05 1.41 0.36 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  1.605 0.05 1.735 0.39 ;
      RECT  2.21 0.05 2.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.74 0.205 1.2 0.31 ;
      RECT  1.11 0.31 1.2 0.71 ;
      RECT  0.94 0.71 1.46 0.78 ;
      RECT  0.94 0.78 1.655 0.8 ;
      RECT  1.36 0.8 1.655 0.89 ;
      RECT  0.94 0.8 1.03 1.36 ;
      RECT  0.76 1.36 1.03 1.47 ;
      RECT  0.045 0.19 0.185 0.36 ;
      RECT  0.045 0.36 0.135 1.25 ;
      RECT  0.045 1.25 0.66 1.35 ;
      RECT  0.56 1.35 0.66 1.56 ;
      RECT  0.045 1.35 0.185 1.63 ;
      RECT  0.56 1.56 1.09 1.66 ;
      RECT  1.295 0.45 1.415 0.53 ;
      RECT  1.295 0.53 1.835 0.62 ;
      RECT  1.745 0.62 1.835 1.045 ;
      RECT  1.13 0.89 1.23 1.045 ;
      RECT  1.13 1.045 1.835 1.135 ;
      RECT  1.295 1.135 1.415 1.225 ;
  END
END SEN_LDNQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_LDNQ_D_4
#      Description : "D-latch, neg-gate, q-only"
#      Equation    : iq,iqn=latch(enable=!G,data_in=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDNQ_D_4
  CLASS CORE ;
  FOREIGN SEN_LDNQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.3 0.65 0.6 ;
      RECT  0.45 0.6 0.65 0.695 ;
      RECT  0.45 0.695 0.55 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.145 0.4 1.24 0.48 ;
      RECT  0.75 0.48 1.24 0.57 ;
      RECT  0.75 0.57 0.85 0.78 ;
      RECT  0.685 0.78 0.85 1.005 ;
      RECT  0.225 0.75 0.325 1.005 ;
      RECT  0.225 1.005 0.85 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0699 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.0 0.45 2.675 0.55 ;
      RECT  2.55 0.55 2.675 1.225 ;
      RECT  2.01 1.225 2.675 1.33 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.445 0.45 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  1.455 1.315 1.585 1.75 ;
      RECT  1.775 1.225 1.895 1.75 ;
      RECT  2.29 1.43 2.415 1.75 ;
      RECT  2.815 1.21 2.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  1.51 0.05 1.62 0.36 ;
      RECT  2.27 0.05 2.44 0.36 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  1.77 0.05 1.9 0.39 ;
      RECT  2.815 0.05 2.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.96 0.205 1.42 0.31 ;
      RECT  1.33 0.31 1.42 0.71 ;
      RECT  1.15 0.71 1.67 0.8 ;
      RECT  1.57 0.8 1.67 0.82 ;
      RECT  1.15 0.8 1.24 1.36 ;
      RECT  1.57 0.82 2.22 0.92 ;
      RECT  0.79 1.36 1.24 1.47 ;
      RECT  0.045 0.215 0.185 0.385 ;
      RECT  0.045 0.385 0.135 1.25 ;
      RECT  0.045 1.25 0.66 1.35 ;
      RECT  0.56 1.35 0.66 1.56 ;
      RECT  0.045 1.35 0.185 1.61 ;
      RECT  0.56 1.56 1.235 1.66 ;
      RECT  1.51 0.45 1.625 0.53 ;
      RECT  1.51 0.53 1.87 0.62 ;
      RECT  1.78 0.62 1.87 0.64 ;
      RECT  1.78 0.64 2.41 0.73 ;
      RECT  2.32 0.73 2.41 1.045 ;
      RECT  1.34 0.89 1.44 1.045 ;
      RECT  1.34 1.045 2.41 1.135 ;
      RECT  1.505 1.135 1.625 1.225 ;
  END
END SEN_LDNQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_LDNRBQ_D_1
#      Description : "D-latch, neg-gate, lo-async-clear, q-only"
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDNRBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_LDNRBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 1.05 0.69 ;
      RECT  0.75 0.69 0.85 0.79 ;
      RECT  0.635 0.79 0.85 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0438 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.255 0.825 0.45 1.02 ;
      RECT  0.255 1.02 1.25 1.13 ;
      RECT  1.14 0.51 1.25 1.02 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.31 2.525 0.49 ;
      RECT  2.35 0.49 2.45 1.31 ;
      RECT  2.35 1.31 2.525 1.49 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.14 1.65 0.23 ;
      RECT  0.55 0.23 0.65 0.585 ;
      RECT  1.55 0.23 1.65 0.9 ;
      RECT  0.365 0.585 0.65 0.69 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0372 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.415 0.44 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.31 1.45 1.44 1.75 ;
      RECT  2.14 1.41 2.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.74 0.05 1.865 0.39 ;
      RECT  2.14 0.05 2.26 0.39 ;
      RECT  0.315 0.05 0.445 0.425 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.77 0.545 2.26 0.665 ;
      RECT  2.17 0.665 2.26 1.2 ;
      RECT  1.875 1.2 2.26 1.29 ;
      RECT  1.875 1.29 1.995 1.53 ;
      RECT  1.665 1.53 1.995 1.64 ;
      RECT  1.98 0.755 2.08 1.02 ;
      RECT  1.645 1.02 2.08 1.11 ;
      RECT  1.645 1.11 1.765 1.25 ;
      RECT  0.95 0.32 1.445 0.42 ;
      RECT  1.355 0.42 1.445 1.22 ;
      RECT  0.755 1.22 1.445 1.25 ;
      RECT  0.755 1.25 1.765 1.35 ;
      RECT  0.055 0.17 0.165 1.23 ;
      RECT  0.055 1.23 0.645 1.32 ;
      RECT  0.555 1.32 0.645 1.45 ;
      RECT  0.055 1.32 0.175 1.62 ;
      RECT  0.555 1.45 1.085 1.56 ;
  END
END SEN_LDNRBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_LDNRBQ_D_2
#      Description : "D-latch, neg-gate, lo-async-clear, q-only"
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDNRBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_LDNRBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 1.25 0.69 ;
      RECT  0.75 0.69 0.85 0.795 ;
      RECT  1.15 0.69 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.265 0.91 1.05 1.0 ;
      RECT  0.265 1.0 1.45 1.09 ;
      RECT  1.34 0.51 1.45 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0615 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.31 2.66 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.14 1.85 0.23 ;
      RECT  0.55 0.23 0.65 0.68 ;
      RECT  1.75 0.23 1.85 0.69 ;
      RECT  0.395 0.68 0.65 0.78 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0417 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.41 0.49 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  1.47 1.46 1.6 1.75 ;
      RECT  2.295 1.21 2.415 1.75 ;
      RECT  2.815 1.21 2.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  1.94 0.05 2.065 0.39 ;
      RECT  2.29 0.05 2.42 0.39 ;
      RECT  0.335 0.05 0.455 0.58 ;
      RECT  2.815 0.05 2.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.975 0.545 2.46 0.665 ;
      RECT  2.37 0.665 2.46 1.015 ;
      RECT  2.025 1.015 2.46 1.105 ;
      RECT  2.025 1.105 2.145 1.53 ;
      RECT  1.77 1.53 2.145 1.64 ;
      RECT  1.81 0.785 2.28 0.895 ;
      RECT  1.81 0.895 1.9 1.25 ;
      RECT  1.1 0.32 1.645 0.42 ;
      RECT  1.555 0.42 1.645 1.25 ;
      RECT  1.555 1.25 1.9 1.255 ;
      RECT  0.92 1.255 1.9 1.37 ;
      RECT  0.065 0.17 0.175 1.19 ;
      RECT  0.065 1.19 0.78 1.28 ;
      RECT  0.69 1.28 0.78 1.475 ;
      RECT  0.065 1.28 0.185 1.61 ;
      RECT  0.69 1.475 1.275 1.585 ;
  END
END SEN_LDNRBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_LDNRBQ_D_4
#      Description : "D-latch, neg-gate, lo-async-clear, q-only"
#      Equation    : iq,iqn=latch(enable=!G,data_in=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDNRBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_LDNRBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 1.25 0.69 ;
      RECT  0.75 0.69 0.85 0.815 ;
      RECT  1.15 0.69 1.25 0.89 ;
      RECT  0.645 0.815 0.85 0.915 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.78 1.05 1.025 ;
      RECT  0.265 1.025 1.05 1.035 ;
      RECT  0.265 1.035 1.48 1.125 ;
      RECT  1.34 0.51 1.48 1.035 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0699 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.31 3.26 0.45 ;
      RECT  2.61 0.45 3.26 0.565 ;
      RECT  3.15 0.565 3.26 1.205 ;
      RECT  2.61 1.205 3.26 1.325 ;
      RECT  3.15 1.325 3.26 1.49 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.14 1.85 0.23 ;
      RECT  0.55 0.23 0.65 0.635 ;
      RECT  1.75 0.23 1.85 0.635 ;
      RECT  0.35 0.635 0.65 0.725 ;
      RECT  1.75 0.635 1.98 0.745 ;
      RECT  0.35 0.725 0.515 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.405 1.415 0.535 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  1.575 1.46 1.705 1.75 ;
      RECT  2.375 1.21 2.495 1.75 ;
      RECT  2.89 1.415 3.02 1.75 ;
      RECT  3.415 1.21 3.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  2.89 0.05 3.02 0.36 ;
      RECT  1.975 0.05 2.105 0.39 ;
      RECT  2.37 0.05 2.5 0.39 ;
      RECT  0.335 0.05 0.455 0.545 ;
      RECT  3.415 0.05 3.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.21 0.32 1.66 0.42 ;
      RECT  1.57 0.42 1.66 0.835 ;
      RECT  1.57 0.835 2.88 0.935 ;
      RECT  1.57 0.935 1.66 1.25 ;
      RECT  0.98 1.25 2.055 1.37 ;
      RECT  2.08 0.5 2.2 0.655 ;
      RECT  2.08 0.655 3.06 0.745 ;
      RECT  2.97 0.745 3.06 1.025 ;
      RECT  2.08 1.025 3.06 1.115 ;
      RECT  2.08 1.115 2.25 1.135 ;
      RECT  2.15 1.135 2.25 1.53 ;
      RECT  1.95 1.53 2.25 1.64 ;
      RECT  0.065 0.19 0.175 1.225 ;
      RECT  0.065 1.225 0.78 1.315 ;
      RECT  0.69 1.315 0.78 1.48 ;
      RECT  0.065 1.315 0.185 1.59 ;
      RECT  0.69 1.48 1.32 1.59 ;
  END
END SEN_LDNRBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_LDPQ_D_1
#      Description : "D-latch, pos-gate, q-only"
#      Equation    : iq,iqn=latch(enable=G,data_in=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDPQ_D_1
  CLASS CORE ;
  FOREIGN SEN_LDPQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.51 ;
      RECT  0.35 0.51 0.65 0.7 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0438 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.235 0.83 0.325 0.91 ;
      RECT  0.235 0.91 0.85 1.0 ;
      RECT  0.75 0.51 0.85 0.91 ;
      RECT  0.35 1.0 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.485 1.945 0.665 ;
      RECT  1.75 0.665 1.85 0.99 ;
      RECT  1.75 0.99 1.945 1.16 ;
    END
    ANTENNADIFFAREA 0.158 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.29 1.495 0.46 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.46 1.495 1.63 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.455 0.05 1.625 0.23 ;
      RECT  0.31 0.05 0.44 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.74 0.205 1.345 0.31 ;
      RECT  1.255 0.31 1.345 0.34 ;
      RECT  1.255 0.34 1.65 0.43 ;
      RECT  1.55 0.43 1.65 1.31 ;
      RECT  0.75 1.31 1.65 1.405 ;
      RECT  1.305 0.52 1.405 0.795 ;
      RECT  1.15 0.795 1.405 0.885 ;
      RECT  1.305 0.885 1.405 0.99 ;
      RECT  1.305 0.99 1.445 1.16 ;
      RECT  0.945 0.425 1.035 1.13 ;
      RECT  0.56 1.13 1.035 1.22 ;
      RECT  0.56 1.22 0.66 1.305 ;
      RECT  0.055 0.17 0.175 0.36 ;
      RECT  0.055 0.36 0.145 1.305 ;
      RECT  0.055 1.305 0.66 1.405 ;
      RECT  0.56 1.405 0.66 1.57 ;
      RECT  0.055 1.405 0.185 1.62 ;
      RECT  0.56 1.57 1.09 1.66 ;
  END
END SEN_LDPQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_LDPQ_D_2
#      Description : "D-latch, pos-gate, q-only"
#      Equation    : iq,iqn=latch(enable=G,data_in=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDPQ_D_2
  CLASS CORE ;
  FOREIGN SEN_LDPQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.3 0.65 0.665 ;
      RECT  0.46 0.665 0.65 0.76 ;
      RECT  0.46 0.76 0.56 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.48 0.85 0.875 ;
      RECT  0.685 0.875 0.85 1.0 ;
      RECT  0.23 0.805 0.33 1.0 ;
      RECT  0.23 1.0 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0549 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.47 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.325 1.43 1.45 1.75 ;
      RECT  1.645 1.43 1.775 1.75 ;
      RECT  2.21 1.21 2.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.325 0.05 1.495 0.25 ;
      RECT  1.64 0.05 1.81 0.305 ;
      RECT  0.32 0.05 0.445 0.39 ;
      RECT  2.21 0.05 2.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.76 0.205 1.235 0.31 ;
      RECT  1.145 0.31 1.235 0.395 ;
      RECT  1.145 0.395 1.845 0.485 ;
      RECT  1.755 0.485 1.845 1.25 ;
      RECT  1.145 1.25 1.845 1.34 ;
      RECT  1.145 1.34 1.235 1.36 ;
      RECT  0.76 1.36 1.235 1.45 ;
      RECT  0.045 0.17 0.185 0.36 ;
      RECT  0.045 0.36 0.135 1.18 ;
      RECT  0.045 1.18 1.055 1.27 ;
      RECT  0.955 0.4 1.055 1.18 ;
      RECT  0.045 1.27 0.66 1.28 ;
      RECT  0.56 1.28 0.66 1.56 ;
      RECT  0.045 1.28 0.185 1.61 ;
      RECT  0.56 1.56 1.09 1.66 ;
      RECT  1.155 0.575 1.55 0.675 ;
      RECT  1.155 0.675 1.255 1.02 ;
      RECT  1.155 1.02 1.55 1.13 ;
  END
END SEN_LDPQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_LDPQ_D_4
#      Description : "D-latch, pos-gate, q-only"
#      Equation    : iq,iqn=latch(enable=G,data_in=D):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDPQ_D_4
  CLASS CORE ;
  FOREIGN SEN_LDPQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.3 0.65 0.74 ;
      RECT  0.45 0.74 0.65 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.005 ;
      RECT  0.225 0.73 0.325 1.005 ;
      RECT  0.225 1.005 0.85 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0627 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.0 0.43 2.66 0.53 ;
      RECT  2.55 0.53 2.66 1.225 ;
      RECT  2.01 1.225 2.66 1.33 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  1.775 1.21 1.895 1.75 ;
      RECT  2.29 1.43 2.42 1.75 ;
      RECT  2.815 1.21 2.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  2.27 0.05 2.44 0.34 ;
      RECT  0.32 0.05 0.445 0.39 ;
      RECT  1.51 0.05 1.62 0.39 ;
      RECT  1.77 0.05 1.9 0.39 ;
      RECT  2.815 0.05 2.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  0.96 0.205 1.42 0.31 ;
      RECT  1.33 0.31 1.42 0.8 ;
      RECT  1.33 0.8 2.21 0.9 ;
      RECT  1.33 0.9 1.42 1.365 ;
      RECT  0.76 1.365 1.42 1.47 ;
      RECT  0.045 0.19 0.185 0.385 ;
      RECT  0.045 0.385 0.135 1.185 ;
      RECT  0.045 1.185 1.24 1.275 ;
      RECT  1.145 0.4 1.24 1.185 ;
      RECT  0.045 1.275 0.66 1.285 ;
      RECT  0.57 1.285 0.66 1.56 ;
      RECT  0.045 1.285 0.185 1.61 ;
      RECT  0.57 1.56 1.12 1.66 ;
      RECT  1.51 0.52 1.625 0.62 ;
      RECT  1.51 0.62 2.41 0.71 ;
      RECT  2.32 0.71 2.41 0.99 ;
      RECT  1.51 0.99 2.41 1.08 ;
      RECT  1.51 1.08 1.625 1.57 ;
      RECT  1.22 1.57 1.625 1.66 ;
  END
END SEN_LDPQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_LDPRBQ_D_1
#      Description : "D-latch, pos-gate, lo-async-clear, q-only"
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDPRBQ_D_1
  CLASS CORE ;
  FOREIGN SEN_LDPRBQ_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 1.05 0.69 ;
      RECT  0.75 0.69 0.85 0.93 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0438 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.255 0.96 0.45 1.23 ;
      RECT  0.255 1.23 0.65 1.32 ;
      RECT  0.55 1.32 0.65 1.45 ;
      RECT  0.55 1.45 1.12 1.56 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.31 2.525 0.49 ;
      RECT  2.35 0.49 2.45 1.31 ;
      RECT  2.35 1.31 2.525 1.49 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.14 1.65 0.23 ;
      RECT  0.55 0.23 0.65 0.585 ;
      RECT  1.55 0.23 1.65 1.12 ;
      RECT  0.395 0.585 0.65 0.69 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0372 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.415 0.44 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.315 1.45 1.445 1.75 ;
      RECT  2.145 1.215 2.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.74 0.05 1.87 0.39 ;
      RECT  2.14 0.05 2.26 0.39 ;
      RECT  0.315 0.05 0.445 0.425 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.76 0.545 2.26 0.665 ;
      RECT  2.17 0.665 2.26 1.025 ;
      RECT  1.93 1.025 2.26 1.115 ;
      RECT  1.93 1.115 2.02 1.475 ;
      RECT  1.62 1.475 2.02 1.585 ;
      RECT  0.055 0.17 0.165 0.78 ;
      RECT  0.055 0.78 0.645 0.87 ;
      RECT  0.555 0.87 0.645 1.02 ;
      RECT  0.055 0.87 0.165 1.62 ;
      RECT  0.555 1.02 1.28 1.13 ;
      RECT  1.18 0.51 1.28 1.02 ;
      RECT  1.74 0.785 2.08 0.895 ;
      RECT  1.74 0.895 1.83 1.22 ;
      RECT  0.93 0.32 1.46 0.42 ;
      RECT  1.37 0.42 1.46 1.22 ;
      RECT  0.785 1.22 1.83 1.34 ;
  END
END SEN_LDPRBQ_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_LDPRBQ_D_2
#      Description : "D-latch, pos-gate, lo-async-clear, q-only"
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDPRBQ_D_2
  CLASS CORE ;
  FOREIGN SEN_LDPRBQ_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 1.25 0.69 ;
      RECT  0.75 0.69 0.85 0.795 ;
      RECT  1.15 0.69 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.054 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.265 1.11 0.65 1.29 ;
      RECT  0.55 1.29 0.65 1.475 ;
      RECT  0.55 1.475 1.275 1.585 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0549 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.31 2.66 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.14 1.85 0.23 ;
      RECT  0.55 0.23 0.65 0.68 ;
      RECT  1.75 0.23 1.85 0.69 ;
      RECT  0.365 0.68 0.65 0.78 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0417 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.415 0.46 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  1.47 1.46 1.6 1.75 ;
      RECT  2.295 1.21 2.415 1.75 ;
      RECT  2.815 1.21 2.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  2.29 0.05 2.42 0.385 ;
      RECT  1.94 0.05 2.07 0.39 ;
      RECT  0.335 0.05 0.455 0.59 ;
      RECT  2.815 0.05 2.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.975 0.545 2.46 0.665 ;
      RECT  2.37 0.665 2.46 1.015 ;
      RECT  2.025 1.015 2.46 1.105 ;
      RECT  2.025 1.105 2.145 1.53 ;
      RECT  1.77 1.53 2.145 1.64 ;
      RECT  0.065 0.17 0.185 0.895 ;
      RECT  0.065 0.895 1.0 0.985 ;
      RECT  0.9 0.985 1.0 1.0 ;
      RECT  0.065 0.985 0.175 1.61 ;
      RECT  0.9 1.0 1.45 1.09 ;
      RECT  1.34 0.51 1.45 1.0 ;
      RECT  1.81 0.785 2.28 0.895 ;
      RECT  1.81 0.895 1.9 1.25 ;
      RECT  1.1 0.32 1.645 0.42 ;
      RECT  1.555 0.42 1.645 1.25 ;
      RECT  1.555 1.25 1.9 1.255 ;
      RECT  0.91 1.255 1.9 1.37 ;
  END
END SEN_LDPRBQ_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_LDPRBQ_D_4
#      Description : "D-latch, pos-gate, lo-async-clear, q-only"
#      Equation    : iq,iqn=latch(enable=G,data_in=D,clear=!RD):Q=iq
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_LDPRBQ_D_4
  CLASS CORE ;
  FOREIGN SEN_LDPRBQ_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 1.25 0.69 ;
      RECT  0.75 0.69 0.85 0.73 ;
      RECT  1.15 0.69 1.25 0.89 ;
      RECT  0.715 0.73 0.85 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D
  PIN G
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.265 1.11 0.45 1.2 ;
      RECT  0.265 1.2 0.85 1.29 ;
      RECT  0.75 1.29 0.85 1.48 ;
      RECT  0.75 1.48 1.37 1.59 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0627 ;
  END G
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.31 3.26 0.45 ;
      RECT  2.58 0.45 3.26 0.565 ;
      RECT  3.15 0.565 3.26 1.205 ;
      RECT  2.61 1.205 3.26 1.325 ;
      RECT  3.15 1.325 3.26 1.49 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END Q
  PIN RD
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.14 1.85 0.23 ;
      RECT  0.55 0.23 0.65 0.51 ;
      RECT  1.75 0.23 1.85 0.635 ;
      RECT  0.35 0.51 0.65 0.6 ;
      RECT  0.35 0.6 0.565 0.84 ;
      RECT  1.75 0.635 1.955 0.745 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END RD
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.48 1.415 0.61 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  1.585 1.46 1.715 1.75 ;
      RECT  2.375 1.215 2.495 1.75 ;
      RECT  2.89 1.415 3.02 1.75 ;
      RECT  3.415 1.21 3.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  2.89 0.05 3.02 0.36 ;
      RECT  0.325 0.05 0.455 0.385 ;
      RECT  1.99 0.05 2.12 0.39 ;
      RECT  2.37 0.05 2.5 0.39 ;
      RECT  3.415 0.05 3.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  OBS
      LAYER M1 ;
      RECT  1.21 0.32 1.66 0.42 ;
      RECT  1.57 0.42 1.66 0.835 ;
      RECT  1.57 0.835 2.88 0.935 ;
      RECT  1.57 0.935 1.66 1.25 ;
      RECT  1.01 1.25 2.06 1.37 ;
      RECT  2.08 0.52 2.2 0.655 ;
      RECT  2.08 0.655 3.06 0.745 ;
      RECT  2.97 0.745 3.06 1.025 ;
      RECT  2.08 1.025 3.06 1.115 ;
      RECT  2.08 1.115 2.25 1.135 ;
      RECT  2.15 1.135 2.25 1.53 ;
      RECT  1.955 1.53 2.25 1.64 ;
      RECT  0.055 0.19 0.175 0.93 ;
      RECT  0.055 0.93 0.63 1.0 ;
      RECT  0.055 1.0 1.48 1.02 ;
      RECT  0.94 0.78 1.05 1.0 ;
      RECT  1.38 0.7 1.48 1.0 ;
      RECT  0.54 1.02 1.48 1.09 ;
      RECT  0.055 1.02 0.175 1.44 ;
      RECT  0.055 1.44 0.3 1.56 ;
  END
END SEN_LDPRBQ_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJ3_0P5
#      Description : "3-input majority"
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJ3_0P5
  CLASS CORE ;
  FOREIGN SEN_MAJ3_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.7 0.65 0.91 ;
      RECT  0.55 0.91 0.85 0.98 ;
      RECT  0.55 0.98 1.365 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.71 ;
      RECT  0.945 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0225 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.595 0.48 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.355 1.39 1.475 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.31 0.05 0.48 0.21 ;
      RECT  1.355 0.05 1.46 0.415 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.21 1.735 0.38 ;
      RECT  1.55 0.38 1.65 0.81 ;
      RECT  1.55 0.81 1.745 0.9 ;
      RECT  1.655 0.9 1.745 1.44 ;
      RECT  1.615 1.44 1.745 1.635 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.57 0.15 1.215 0.24 ;
      RECT  0.57 0.24 0.66 0.305 ;
      RECT  1.095 0.24 1.215 0.455 ;
      RECT  0.065 0.2 0.185 0.305 ;
      RECT  0.065 0.305 0.66 0.395 ;
      RECT  0.81 0.34 0.98 0.43 ;
      RECT  0.81 0.43 0.9 0.52 ;
      RECT  0.355 0.52 0.9 0.61 ;
      RECT  0.355 0.61 0.445 1.18 ;
      RECT  0.355 1.18 1.565 1.27 ;
      RECT  1.475 1.01 1.565 1.18 ;
      RECT  0.81 1.27 0.98 1.48 ;
      RECT  0.065 1.37 0.72 1.46 ;
      RECT  0.63 1.46 0.72 1.57 ;
      RECT  0.065 1.46 0.185 1.585 ;
      RECT  0.63 1.57 1.215 1.66 ;
      RECT  1.095 1.375 1.215 1.57 ;
  END
END SEN_MAJ3_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJ3_1
#      Description : "3-input majority"
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJ3_1
  CLASS CORE ;
  FOREIGN SEN_MAJ3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.71 0.845 1.245 ;
      RECT  0.745 1.245 1.46 1.335 ;
      RECT  1.34 0.75 1.46 1.245 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.115 0.71 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.34 1.615 0.51 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.44 1.425 1.57 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.36 0.05 0.49 0.39 ;
      RECT  1.445 0.05 1.575 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.74 0.31 1.86 0.49 ;
      RECT  1.76 0.49 1.86 1.11 ;
      RECT  1.74 1.11 1.86 1.49 ;
    END
    ANTENNADIFFAREA 0.238 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.615 0.24 1.35 0.36 ;
      RECT  0.615 0.36 0.715 0.48 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 0.715 0.59 ;
      RECT  0.935 0.49 1.45 0.56 ;
      RECT  0.935 0.56 1.67 0.585 ;
      RECT  1.36 0.585 1.67 0.655 ;
      RECT  0.935 0.585 1.025 1.155 ;
      RECT  1.57 0.655 1.67 0.955 ;
      RECT  0.065 1.425 1.35 1.525 ;
      RECT  0.065 1.525 0.185 1.62 ;
  END
END SEN_MAJ3_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJ3_1P5
#      Description : "3-input majority"
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJ3_1P5
  CLASS CORE ;
  FOREIGN SEN_MAJ3_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.06 ;
      RECT  0.75 1.06 1.295 1.15 ;
      RECT  1.195 0.685 1.295 1.06 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1134 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.665 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1134 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.64 1.105 0.935 ;
      LAYER M2 ;
      RECT  0.91 0.75 1.485 0.85 ;
      LAYER V1 ;
      RECT  0.95 0.75 1.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0567 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.42 0.435 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.295 1.45 1.415 1.75 ;
      RECT  1.805 1.415 1.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.295 0.05 1.415 0.345 ;
      RECT  0.315 0.05 0.435 0.385 ;
      RECT  1.805 0.05 1.935 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.57 0.31 1.675 0.475 ;
      RECT  1.57 0.475 1.85 0.565 ;
      RECT  1.75 0.565 1.85 1.11 ;
      RECT  1.57 1.11 1.85 1.3 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.57 0.2 1.205 0.32 ;
      RECT  0.57 0.32 0.66 0.475 ;
      RECT  0.055 0.165 0.175 0.475 ;
      RECT  0.055 0.475 0.66 0.565 ;
      RECT  0.75 0.435 1.48 0.55 ;
      RECT  1.39 0.55 1.48 0.795 ;
      RECT  1.39 0.795 1.66 0.905 ;
      RECT  1.39 0.905 1.48 1.24 ;
      RECT  0.71 1.24 1.48 1.36 ;
      RECT  0.055 1.24 0.615 1.33 ;
      RECT  0.525 1.33 0.615 1.465 ;
      RECT  0.055 1.33 0.175 1.63 ;
      RECT  0.525 1.465 1.205 1.585 ;
  END
END SEN_MAJ3_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJ3_2
#      Description : "3-input majority"
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJ3_2
  CLASS CORE ;
  FOREIGN SEN_MAJ3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.85 0.89 ;
      RECT  2.75 0.89 2.85 1.0 ;
      RECT  2.75 1.0 3.65 1.09 ;
      RECT  3.55 0.71 3.65 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.71 ;
      RECT  0.75 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.45 0.71 ;
      RECT  2.95 0.71 3.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.585 1.21 0.705 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.64 1.61 1.81 1.75 ;
      RECT  3.49 1.61 3.66 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  1.66 0.05 1.79 0.23 ;
      RECT  2.16 0.05 2.29 0.23 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.12 0.05 1.23 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.325 0.31 0.45 0.69 ;
      RECT  0.325 0.69 0.415 1.31 ;
      RECT  0.325 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.65 0.14 3.935 0.23 ;
      RECT  3.815 0.23 3.935 1.185 ;
      RECT  0.515 0.755 0.625 1.01 ;
      RECT  0.515 1.01 2.555 1.12 ;
      RECT  2.435 1.12 2.555 1.185 ;
      RECT  2.435 1.185 3.935 1.3 ;
      RECT  0.82 0.24 1.03 0.36 ;
      RECT  0.94 0.36 1.03 0.51 ;
      RECT  0.94 0.51 3.15 0.62 ;
      RECT  1.34 0.32 3.7 0.42 ;
      RECT  0.82 1.21 2.32 1.315 ;
      RECT  1.34 1.405 3.935 1.52 ;
      RECT  3.815 1.52 3.935 1.62 ;
  END
END SEN_MAJ3_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJ3_4
#      Description : "3-input majority"
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJ3_4
  CLASS CORE ;
  FOREIGN SEN_MAJ3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.795 4.105 0.895 ;
      RECT  2.95 0.895 3.45 1.09 ;
      RECT  3.35 1.09 3.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.435 0.71 5.25 0.895 ;
      RECT  1.55 0.71 2.65 0.895 ;
      LAYER M2 ;
      RECT  2.31 0.75 4.775 0.85 ;
      LAYER V1 ;
      RECT  4.435 0.75 4.535 0.85 ;
      RECT  4.635 0.75 4.735 0.85 ;
      RECT  2.35 0.75 2.45 0.85 ;
      RECT  2.55 0.75 2.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.504 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.79 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.36 1.425 1.49 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  1.88 1.425 2.01 1.75 ;
      RECT  2.4 1.425 2.53 1.75 ;
      RECT  2.92 1.425 3.05 1.75 ;
      RECT  4.73 1.41 4.86 1.75 ;
      RECT  5.25 1.41 5.38 1.75 ;
      RECT  5.765 1.21 5.885 1.75 ;
      RECT  6.28 1.41 6.41 1.75 ;
      RECT  6.81 1.21 6.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  2.38 0.05 2.55 0.315 ;
      RECT  2.9 0.05 3.07 0.315 ;
      RECT  1.36 0.05 1.49 0.39 ;
      RECT  1.88 0.05 2.01 0.39 ;
      RECT  4.73 0.05 4.855 0.39 ;
      RECT  5.25 0.05 5.38 0.39 ;
      RECT  6.28 0.05 6.41 0.39 ;
      RECT  5.765 0.05 5.885 0.59 ;
      RECT  6.81 0.05 6.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.025 0.51 6.66 0.69 ;
      RECT  6.55 0.69 6.66 1.11 ;
      RECT  6.025 1.11 6.66 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.215 1.225 0.335 ;
      RECT  0.065 0.335 0.185 0.39 ;
      RECT  1.105 0.335 1.225 0.485 ;
      RECT  1.105 0.485 3.33 0.505 ;
      RECT  2.145 0.405 3.33 0.485 ;
      RECT  1.105 0.505 2.265 0.605 ;
      RECT  3.41 0.24 4.595 0.36 ;
      RECT  4.475 0.36 4.595 0.485 ;
      RECT  4.475 0.485 5.675 0.605 ;
      RECT  5.55 0.79 6.44 0.895 ;
      RECT  5.55 0.895 5.65 1.01 ;
      RECT  3.49 0.505 4.335 0.595 ;
      RECT  2.755 0.595 4.335 0.625 ;
      RECT  2.755 0.625 3.6 0.685 ;
      RECT  4.215 0.625 4.335 1.01 ;
      RECT  2.755 0.685 2.845 1.01 ;
      RECT  0.27 0.485 0.99 0.605 ;
      RECT  0.9 0.605 0.99 1.01 ;
      RECT  0.34 1.01 2.845 1.13 ;
      RECT  4.215 1.01 5.65 1.1 ;
      RECT  4.215 1.1 4.335 1.135 ;
      RECT  0.34 1.13 0.445 1.24 ;
      RECT  3.64 1.135 4.335 1.255 ;
      RECT  4.475 1.19 5.675 1.305 ;
      RECT  4.475 1.305 4.595 1.44 ;
      RECT  3.41 1.44 4.595 1.56 ;
      RECT  1.105 1.22 3.26 1.335 ;
      RECT  3.17 1.335 3.26 1.37 ;
      RECT  1.105 1.335 1.225 1.4 ;
      RECT  3.17 1.37 3.305 1.54 ;
      RECT  0.065 1.4 1.225 1.52 ;
      RECT  0.065 1.52 0.185 1.61 ;
  END
END SEN_MAJ3_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJ3_6
#      Description : "3-input majority"
#      Equation    : X=(A1&A2)|(A1&A3)|(A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJ3_6
  CLASS CORE ;
  FOREIGN SEN_MAJ3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 4.13 0.89 ;
      RECT  3.35 0.89 3.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.453 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.51 5.45 0.71 ;
      RECT  4.75 0.71 5.45 0.89 ;
      RECT  2.95 0.51 3.05 0.71 ;
      RECT  1.35 0.71 3.05 0.89 ;
      LAYER M2 ;
      RECT  2.905 0.55 5.49 0.65 ;
      LAYER V1 ;
      RECT  5.35 0.55 5.45 0.65 ;
      RECT  2.95 0.55 3.05 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.453 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2265 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.365 1.45 1.485 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  1.885 1.45 2.005 1.75 ;
      RECT  2.415 1.45 2.535 1.75 ;
      RECT  2.935 1.45 3.055 1.75 ;
      RECT  4.755 1.45 4.875 1.75 ;
      RECT  5.275 1.45 5.395 1.75 ;
      RECT  5.785 1.215 5.905 1.75 ;
      RECT  6.305 1.395 6.425 1.75 ;
      RECT  6.825 1.395 6.945 1.75 ;
      RECT  7.36 1.21 7.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  1.345 0.05 1.465 0.345 ;
      RECT  1.885 0.05 2.01 0.345 ;
      RECT  2.405 0.05 2.53 0.345 ;
      RECT  4.755 0.05 4.875 0.345 ;
      RECT  6.305 0.05 6.425 0.345 ;
      RECT  6.825 0.05 6.945 0.35 ;
      RECT  5.295 0.05 5.415 0.385 ;
      RECT  2.945 0.05 3.065 0.39 ;
      RECT  5.765 0.05 5.885 0.585 ;
      RECT  7.36 0.05 7.48 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.045 0.51 7.25 0.69 ;
      RECT  6.92 0.69 7.05 1.11 ;
      RECT  6.35 1.11 7.19 1.19 ;
      RECT  5.995 1.19 7.19 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.2 1.225 0.32 ;
      RECT  0.065 0.32 0.185 0.43 ;
      RECT  1.105 0.32 1.225 0.445 ;
      RECT  1.105 0.445 2.835 0.56 ;
      RECT  3.925 0.24 4.615 0.35 ;
      RECT  4.495 0.35 4.615 0.445 ;
      RECT  4.495 0.445 5.185 0.56 ;
      RECT  6.02 0.785 6.8 0.895 ;
      RECT  6.02 0.895 6.11 0.98 ;
      RECT  3.17 0.44 4.38 0.55 ;
      RECT  4.275 0.55 4.38 0.98 ;
      RECT  3.17 0.55 3.26 1.06 ;
      RECT  4.275 0.98 6.11 1.07 ;
      RECT  0.275 0.43 0.99 0.55 ;
      RECT  0.9 0.55 0.99 1.06 ;
      RECT  0.9 1.06 3.26 1.15 ;
      RECT  4.275 1.07 4.38 1.14 ;
      RECT  3.665 1.14 4.38 1.26 ;
      RECT  0.9 1.15 0.99 1.24 ;
      RECT  0.275 1.24 0.99 1.36 ;
      RECT  1.105 1.24 3.26 1.36 ;
      RECT  3.17 1.36 3.26 1.39 ;
      RECT  1.105 1.36 1.225 1.45 ;
      RECT  3.17 1.39 3.325 1.56 ;
      RECT  0.065 1.335 0.185 1.45 ;
      RECT  0.065 1.45 1.225 1.56 ;
      RECT  4.495 1.24 5.695 1.36 ;
      RECT  4.495 1.36 4.615 1.44 ;
      RECT  3.43 1.44 4.615 1.56 ;
  END
END SEN_MAJ3_6
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_1
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_1
  CLASS CORE ;
  FOREIGN SEN_MAJI3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.0 ;
      RECT  0.15 1.0 1.05 1.09 ;
      RECT  0.95 0.71 1.05 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.895 ;
      LAYER M2 ;
      RECT  0.41 0.75 0.93 0.85 ;
      LAYER V1 ;
      RECT  0.45 0.75 0.55 0.85 ;
      RECT  0.65 0.75 0.75 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.59 1.41 0.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.45 1.25 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.86 0.17 1.52 0.29 ;
      RECT  1.405 0.29 1.52 0.39 ;
      RECT  0.86 0.29 0.95 0.51 ;
      RECT  0.34 0.38 0.455 0.51 ;
      RECT  0.34 0.51 0.95 0.6 ;
      RECT  0.305 1.21 0.94 1.32 ;
      RECT  0.85 1.32 0.94 1.51 ;
      RECT  0.85 1.51 1.52 1.63 ;
      RECT  1.4 1.41 1.52 1.51 ;
  END
END SEN_MAJI3_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_2
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_2
  CLASS CORE ;
  FOREIGN SEN_MAJI3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.84 1.72 0.9 ;
      RECT  1.55 0.9 2.18 0.98 ;
      RECT  2.005 0.835 2.18 0.9 ;
      RECT  1.55 0.98 2.05 1.1 ;
      RECT  1.95 1.1 2.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.625 0.7 2.93 0.91 ;
      RECT  0.75 0.7 1.05 0.9 ;
      LAYER M2 ;
      RECT  0.895 0.75 2.8 0.85 ;
      LAYER V1 ;
      RECT  2.655 0.75 2.755 0.85 ;
      RECT  0.935 0.75 1.035 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.845 1.41 0.975 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.365 1.41 1.495 1.75 ;
      RECT  2.655 1.485 2.825 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  2.655 0.05 2.825 0.315 ;
      RECT  0.845 0.05 0.975 0.36 ;
      RECT  1.365 0.05 1.495 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.825 0.51 2.265 0.6 ;
      RECT  1.825 0.6 2.45 0.66 ;
      RECT  1.15 0.66 2.45 0.7 ;
      RECT  1.15 0.7 1.915 0.75 ;
      RECT  2.35 0.7 2.45 1.1 ;
      RECT  1.15 0.75 1.25 1.01 ;
      RECT  0.34 0.45 0.45 1.01 ;
      RECT  0.34 1.01 1.25 1.1 ;
      RECT  0.34 1.1 0.45 1.29 ;
      RECT  2.145 1.1 2.45 1.2 ;
      RECT  2.145 1.2 2.255 1.32 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.17 0.715 0.305 ;
      RECT  0.07 0.305 0.19 0.39 ;
      RECT  0.585 0.305 0.715 0.45 ;
      RECT  0.585 0.45 1.735 0.57 ;
      RECT  1.63 0.35 1.735 0.45 ;
      RECT  1.83 0.29 2.52 0.405 ;
      RECT  1.83 0.405 3.13 0.41 ;
      RECT  2.4 0.41 3.13 0.51 ;
      RECT  0.585 1.195 1.8 1.315 ;
      RECT  0.585 1.315 0.715 1.41 ;
      RECT  0.07 1.41 0.715 1.5 ;
      RECT  0.07 1.5 0.19 1.63 ;
      RECT  2.4 1.29 3.13 1.395 ;
      RECT  2.4 1.395 2.52 1.44 ;
      RECT  1.83 1.44 2.52 1.56 ;
  END
END SEN_MAJI3_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_4
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_4
  CLASS CORE ;
  FOREIGN SEN_MAJI3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.835 4.085 0.94 ;
      RECT  2.75 0.94 3.65 1.09 ;
      RECT  3.55 1.09 3.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 5.25 0.895 ;
      RECT  1.35 0.71 2.45 0.895 ;
      LAYER M2 ;
      RECT  2.11 0.75 4.89 0.85 ;
      LAYER V1 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  2.35 0.75 2.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.855 0.895 ;
      RECT  0.15 0.895 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.365 1.41 1.495 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  1.885 1.41 2.015 1.75 ;
      RECT  2.415 1.41 2.545 1.75 ;
      RECT  2.955 1.41 3.085 1.75 ;
      RECT  4.79 1.24 4.91 1.75 ;
      RECT  5.32 1.24 5.44 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  1.345 0.05 1.515 0.345 ;
      RECT  1.865 0.05 2.035 0.345 ;
      RECT  2.385 0.05 2.555 0.345 ;
      RECT  2.905 0.05 3.075 0.345 ;
      RECT  4.755 0.05 4.885 0.39 ;
      RECT  5.305 0.05 5.435 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 4.45 0.635 ;
      RECT  2.55 0.635 4.45 0.725 ;
      RECT  2.55 0.725 2.65 1.005 ;
      RECT  4.35 0.725 4.45 1.11 ;
      RECT  0.28 0.46 1.05 0.58 ;
      RECT  0.95 0.58 1.05 1.005 ;
      RECT  0.95 1.005 2.65 1.095 ;
      RECT  0.95 1.095 1.05 1.11 ;
      RECT  0.34 1.11 1.05 1.29 ;
      RECT  3.74 1.11 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.2 1.255 0.32 ;
      RECT  0.07 0.32 0.19 0.39 ;
      RECT  1.15 0.32 1.255 0.435 ;
      RECT  1.15 0.435 3.355 0.545 ;
      RECT  3.405 0.24 4.65 0.36 ;
      RECT  4.55 0.36 4.65 0.48 ;
      RECT  4.55 0.48 5.715 0.59 ;
      RECT  5.595 0.37 5.715 0.48 ;
      RECT  4.54 1.03 5.715 1.15 ;
      RECT  5.595 1.15 5.715 1.25 ;
      RECT  4.54 1.15 4.65 1.44 ;
      RECT  3.43 1.44 4.65 1.56 ;
      RECT  1.15 1.2 3.4 1.32 ;
      RECT  1.15 1.32 1.255 1.48 ;
      RECT  0.07 1.41 0.19 1.48 ;
      RECT  0.07 1.48 1.255 1.6 ;
  END
END SEN_MAJI3_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_3
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_3
  CLASS CORE ;
  FOREIGN SEN_MAJI3_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 2.45 0.9 ;
      RECT  1.35 0.9 1.48 1.09 ;
      LAYER M2 ;
      RECT  1.085 0.95 1.775 1.05 ;
      LAYER V1 ;
      RECT  1.35 0.95 1.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.84 0.71 3.315 0.89 ;
      RECT  0.35 0.71 0.85 0.89 ;
      LAYER M2 ;
      RECT  0.475 0.75 3.49 0.85 ;
      LAYER V1 ;
      RECT  2.955 0.75 3.055 0.85 ;
      RECT  3.2 0.75 3.3 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.25 0.93 ;
      RECT  4.15 0.93 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  2.135 1.44 2.255 1.75 ;
      RECT  2.655 1.44 2.775 1.75 ;
      RECT  3.175 1.44 3.295 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.585 0.05 0.705 0.36 ;
      RECT  2.135 0.05 2.255 0.385 ;
      RECT  2.655 0.05 2.775 0.385 ;
      RECT  3.175 0.05 3.295 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.23 0.315 4.33 0.485 ;
      RECT  3.645 0.485 4.33 0.59 ;
      RECT  3.75 0.59 3.85 1.05 ;
      RECT  1.625 1.05 3.85 1.14 ;
      RECT  1.625 1.14 1.745 1.19 ;
      RECT  3.75 1.14 3.85 1.205 ;
      RECT  1.625 0.32 1.745 0.425 ;
      RECT  1.08 0.425 1.745 0.545 ;
      RECT  1.15 0.545 1.25 1.11 ;
      RECT  1.1 1.11 1.25 1.19 ;
      RECT  1.1 1.19 1.745 1.29 ;
      RECT  3.75 1.205 4.325 1.295 ;
      RECT  4.225 1.295 4.325 1.425 ;
    END
    ANTENNADIFFAREA 0.778 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.85 0.215 1.51 0.335 ;
      RECT  0.85 0.335 0.955 0.45 ;
      RECT  0.275 0.45 0.955 0.555 ;
      RECT  3.435 0.215 4.125 0.335 ;
      RECT  3.435 0.335 3.555 0.475 ;
      RECT  1.875 0.29 1.995 0.475 ;
      RECT  1.875 0.475 3.555 0.595 ;
      RECT  0.275 1.23 0.965 1.35 ;
      RECT  0.845 1.35 0.965 1.405 ;
      RECT  0.845 1.405 1.535 1.525 ;
      RECT  1.875 1.23 3.555 1.35 ;
      RECT  3.435 1.35 3.555 1.405 ;
      RECT  1.875 1.35 1.995 1.45 ;
      RECT  3.435 1.405 4.125 1.525 ;
  END
END SEN_MAJI3_3
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_5
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_5
  CLASS CORE ;
  FOREIGN SEN_MAJI3_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.915 0.785 3.895 0.895 ;
      RECT  1.915 0.895 2.05 1.145 ;
      LAYER M2 ;
      RECT  1.91 0.95 2.575 1.05 ;
      LAYER V1 ;
      RECT  1.95 0.95 2.05 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.405 0.74 5.175 0.9 ;
      RECT  0.515 0.745 1.37 0.89 ;
      LAYER M2 ;
      RECT  0.71 0.75 5.15 0.85 ;
      LAYER V1 ;
      RECT  4.455 0.75 4.555 0.85 ;
      RECT  4.7 0.75 4.8 0.85 ;
      RECT  4.945 0.75 5.045 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
      RECT  0.995 0.75 1.095 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.015 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  3.175 1.44 3.295 1.75 ;
      RECT  3.695 1.44 3.815 1.75 ;
      RECT  4.215 1.44 4.335 1.75 ;
      RECT  4.735 1.44 4.855 1.75 ;
      RECT  5.255 1.44 5.375 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  3.695 0.05 3.815 0.36 ;
      RECT  4.215 0.05 4.335 0.36 ;
      RECT  4.735 0.05 4.855 0.36 ;
      RECT  5.255 0.05 5.375 0.36 ;
      RECT  0.585 0.05 0.705 0.385 ;
      RECT  1.105 0.05 1.225 0.385 ;
      RECT  3.175 0.05 3.295 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.815 0.29 6.935 0.475 ;
      RECT  5.75 0.475 6.935 0.595 ;
      RECT  5.75 0.595 5.88 1.035 ;
      RECT  2.65 1.035 5.88 1.11 ;
      RECT  2.65 1.11 6.45 1.145 ;
      RECT  5.75 1.145 6.45 1.205 ;
      RECT  2.65 1.145 2.785 1.26 ;
      RECT  5.75 1.205 6.935 1.295 ;
      RECT  1.625 0.51 2.785 0.69 ;
      RECT  1.625 0.69 1.745 1.26 ;
      RECT  1.625 1.26 2.785 1.39 ;
      RECT  6.815 1.295 6.935 1.425 ;
    END
    ANTENNADIFFAREA 1.21 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.365 0.2 2.575 0.32 ;
      RECT  1.365 0.32 1.485 0.51 ;
      RECT  0.275 0.51 1.485 0.63 ;
      RECT  5.52 0.215 6.725 0.335 ;
      RECT  5.52 0.335 5.635 0.475 ;
      RECT  2.915 0.29 3.035 0.475 ;
      RECT  2.915 0.475 5.635 0.595 ;
      RECT  0.275 1.24 1.485 1.35 ;
      RECT  1.365 1.35 1.485 1.48 ;
      RECT  1.365 1.48 2.575 1.6 ;
      RECT  2.915 1.235 5.635 1.35 ;
      RECT  5.515 1.35 5.635 1.43 ;
      RECT  2.915 1.35 3.035 1.46 ;
      RECT  5.515 1.43 6.725 1.55 ;
  END
END SEN_MAJI3_5
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_6
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_6
  CLASS CORE ;
  FOREIGN SEN_MAJI3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.2 0.48 3.305 0.74 ;
      RECT  2.515 0.74 4.69 0.89 ;
      LAYER M2 ;
      RECT  2.855 0.55 3.55 0.65 ;
      LAYER V1 ;
      RECT  3.2 0.55 3.3 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.71 6.485 0.89 ;
      RECT  0.515 0.73 1.485 0.905 ;
      LAYER M2 ;
      RECT  0.52 0.75 6.38 0.85 ;
      LAYER V1 ;
      RECT  5.44 0.75 5.54 0.85 ;
      RECT  5.84 0.75 5.94 0.85 ;
      RECT  6.24 0.75 6.34 0.85 ;
      RECT  0.815 0.75 0.915 0.85 ;
      RECT  1.2 0.75 1.3 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.21 0.71 8.25 0.89 ;
      RECT  8.15 0.89 8.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.445 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  0.845 1.44 0.965 1.75 ;
      RECT  1.365 1.44 1.485 1.75 ;
      RECT  3.67 1.495 3.84 1.75 ;
      RECT  4.19 1.495 4.36 1.75 ;
      RECT  4.71 1.495 4.88 1.75 ;
      RECT  5.23 1.495 5.4 1.75 ;
      RECT  5.75 1.495 5.92 1.75 ;
      RECT  6.27 1.495 6.44 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  3.695 0.05 3.815 0.36 ;
      RECT  4.215 0.05 4.335 0.36 ;
      RECT  4.735 0.05 4.855 0.36 ;
      RECT  5.255 0.05 5.375 0.36 ;
      RECT  5.775 0.05 5.895 0.36 ;
      RECT  6.295 0.05 6.415 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.79 0.45 8.025 0.57 ;
      RECT  6.79 0.57 7.08 0.59 ;
      RECT  6.95 0.59 7.08 1.055 ;
      RECT  3.23 1.055 7.08 1.11 ;
      RECT  1.855 0.45 3.075 0.58 ;
      RECT  2.15 0.58 2.28 1.11 ;
      RECT  1.88 1.11 8.05 1.185 ;
      RECT  1.88 1.185 3.36 1.29 ;
      RECT  6.78 1.185 8.05 1.29 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.615 0.21 3.355 0.34 ;
      RECT  1.615 0.34 1.745 0.45 ;
      RECT  0.065 0.29 0.185 0.45 ;
      RECT  0.065 0.45 1.745 0.58 ;
      RECT  6.545 0.21 8.285 0.34 ;
      RECT  6.545 0.34 6.675 0.465 ;
      RECT  3.41 0.465 6.675 0.595 ;
      RECT  0.065 1.215 1.745 1.345 ;
      RECT  0.065 1.345 0.185 1.435 ;
      RECT  1.625 1.345 1.745 1.455 ;
      RECT  1.625 1.455 3.355 1.585 ;
      RECT  3.45 1.275 6.69 1.405 ;
      RECT  6.53 1.405 6.69 1.44 ;
      RECT  3.45 1.405 3.54 1.5 ;
      RECT  6.53 1.44 8.285 1.585 ;
  END
END SEN_MAJI3_6
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_8
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_8
  CLASS CORE ;
  FOREIGN SEN_MAJI3_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.285 0.465 4.385 0.765 ;
      RECT  3.295 0.765 6.705 0.875 ;
      LAYER M2 ;
      RECT  3.895 0.55 4.555 0.65 ;
      LAYER V1 ;
      RECT  4.285 0.55 4.385 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.915 0.745 8.76 0.875 ;
      RECT  0.55 0.71 1.89 0.89 ;
      LAYER M2 ;
      RECT  1.215 0.75 7.985 0.85 ;
      LAYER V1 ;
      RECT  7.045 0.75 7.145 0.85 ;
      RECT  7.445 0.75 7.545 0.85 ;
      RECT  7.845 0.75 7.945 0.85 ;
      RECT  1.26 0.75 1.36 0.85 ;
      RECT  1.505 0.75 1.605 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.235 0.71 10.85 0.89 ;
      RECT  10.75 0.89 10.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.445 1.75 ;
      RECT  0.0 1.75 11.0 1.85 ;
      RECT  0.845 1.44 0.965 1.75 ;
      RECT  1.365 1.44 1.485 1.75 ;
      RECT  1.885 1.44 2.005 1.75 ;
      RECT  4.725 1.48 4.895 1.75 ;
      RECT  5.245 1.48 5.415 1.75 ;
      RECT  5.765 1.48 5.935 1.75 ;
      RECT  6.285 1.48 6.455 1.75 ;
      RECT  6.805 1.48 6.975 1.75 ;
      RECT  7.325 1.48 7.495 1.75 ;
      RECT  7.845 1.48 8.015 1.75 ;
      RECT  8.365 1.48 8.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      RECT  0.3 0.05 0.47 0.345 ;
      RECT  0.82 0.05 0.99 0.345 ;
      RECT  1.34 0.05 1.51 0.345 ;
      RECT  1.885 0.05 2.005 0.345 ;
      RECT  4.725 0.05 4.895 0.355 ;
      RECT  5.245 0.05 5.415 0.355 ;
      RECT  5.765 0.05 5.935 0.355 ;
      RECT  6.285 0.05 6.455 0.355 ;
      RECT  6.805 0.05 6.975 0.355 ;
      RECT  7.325 0.05 7.495 0.355 ;
      RECT  7.845 0.05 8.015 0.355 ;
      RECT  8.365 0.05 8.51 0.355 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.885 0.45 10.615 0.59 ;
      RECT  8.885 0.59 9.12 0.595 ;
      RECT  8.95 0.595 9.12 0.975 ;
      RECT  4.23 0.975 9.12 1.11 ;
      RECT  2.405 0.51 4.11 0.64 ;
      RECT  2.405 0.64 3.12 0.69 ;
      RECT  2.95 0.69 3.12 1.11 ;
      RECT  2.405 1.11 10.65 1.13 ;
      RECT  2.405 1.13 4.4 1.29 ;
      RECT  8.95 1.13 10.65 1.29 ;
    END
    ANTENNADIFFAREA 1.736 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.095 0.185 4.385 0.355 ;
      RECT  2.095 0.355 2.265 0.435 ;
      RECT  0.065 0.435 2.265 0.605 ;
      RECT  8.6 0.19 10.85 0.36 ;
      RECT  8.6 0.36 8.77 0.445 ;
      RECT  4.505 0.445 8.77 0.615 ;
      RECT  0.065 1.18 2.265 1.35 ;
      RECT  2.095 1.35 2.265 1.44 ;
      RECT  2.095 1.44 4.37 1.61 ;
      RECT  4.49 1.22 8.795 1.39 ;
      RECT  8.625 1.39 8.795 1.435 ;
      RECT  8.625 1.435 10.875 1.605 ;
  END
END SEN_MAJI3_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_T_1
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_T_1
  CLASS CORE ;
  FOREIGN SEN_MAJI3_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.005 ;
      RECT  0.35 1.005 1.65 1.095 ;
      RECT  1.545 0.71 1.65 1.005 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.33 0.89 ;
      LAYER M2 ;
      RECT  0.85 0.75 1.415 0.85 ;
      LAYER V1 ;
      RECT  1.01 0.75 1.11 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  0.615 1.44 0.735 1.75 ;
      RECT  1.18 1.44 1.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.615 0.05 0.735 0.36 ;
      RECT  1.18 0.05 1.3 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.635 0.425 1.85 0.545 ;
      RECT  1.75 0.545 1.85 1.19 ;
      RECT  1.635 1.19 1.85 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.405 0.215 2.115 0.335 ;
      RECT  1.405 0.335 1.495 0.45 ;
      RECT  0.275 0.45 1.495 0.57 ;
      RECT  0.275 1.23 1.495 1.35 ;
      RECT  1.405 1.35 1.495 1.455 ;
      RECT  1.405 1.455 2.115 1.575 ;
  END
END SEN_MAJI3_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_T_2
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_T_2
  CLASS CORE ;
  FOREIGN SEN_MAJI3_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.045 0.5 1.145 0.71 ;
      RECT  1.045 0.71 2.05 0.89 ;
      LAYER M2 ;
      RECT  0.825 0.55 1.41 0.65 ;
      LAYER V1 ;
      RECT  1.045 0.55 1.145 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  0.35 0.71 0.695 0.89 ;
      LAYER M2 ;
      RECT  0.39 0.75 2.76 0.85 ;
      LAYER V1 ;
      RECT  2.6 0.75 2.7 0.85 ;
      RECT  0.43 0.75 0.53 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.51 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.42 0.445 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  1.615 1.44 1.735 1.75 ;
      RECT  2.135 1.44 2.255 1.75 ;
      RECT  2.655 1.44 2.775 1.75 ;
      RECT  3.175 1.44 3.295 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.325 0.05 0.445 0.365 ;
      RECT  1.615 0.05 1.735 0.385 ;
      RECT  2.135 0.05 2.255 0.385 ;
      RECT  2.655 0.05 2.775 0.385 ;
      RECT  3.175 0.05 3.295 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.67 0.44 3.85 0.56 ;
      RECT  3.75 0.56 3.85 1.055 ;
      RECT  0.82 0.495 0.95 1.055 ;
      RECT  0.82 1.055 3.85 1.155 ;
      RECT  3.75 1.155 3.85 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.435 0.215 4.125 0.335 ;
      RECT  3.435 0.335 3.555 0.475 ;
      RECT  1.3 0.475 3.555 0.595 ;
      RECT  0.585 0.22 1.25 0.34 ;
      RECT  0.585 0.34 0.705 0.455 ;
      RECT  0.065 0.26 0.185 0.455 ;
      RECT  0.065 0.455 0.705 0.545 ;
      RECT  0.065 1.24 0.705 1.33 ;
      RECT  0.585 1.33 0.705 1.415 ;
      RECT  0.065 1.33 0.185 1.435 ;
      RECT  0.585 1.415 1.275 1.535 ;
      RECT  1.365 1.245 3.545 1.35 ;
      RECT  3.44 1.35 3.545 1.405 ;
      RECT  1.365 1.35 1.465 1.46 ;
      RECT  3.44 1.405 4.125 1.525 ;
  END
END SEN_MAJI3_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_T_3
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_T_3
  CLASS CORE ;
  FOREIGN SEN_MAJI3_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.05 0.775 ;
      RECT  3.95 0.775 4.56 0.895 ;
      RECT  3.95 0.895 4.05 1.005 ;
      RECT  0.55 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.005 ;
      RECT  1.35 1.005 4.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5832 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 0.71 ;
      RECT  1.95 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5832 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.71 5.65 0.775 ;
      RECT  4.985 0.775 5.65 0.895 ;
      RECT  5.55 0.895 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  1.625 1.44 1.745 1.75 ;
      RECT  2.145 1.44 2.265 1.75 ;
      RECT  2.665 1.44 2.785 1.75 ;
      RECT  3.185 1.215 3.305 1.75 ;
      RECT  3.705 1.44 3.825 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  0.585 0.05 0.705 0.36 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  1.625 0.05 1.745 0.36 ;
      RECT  2.145 0.05 2.265 0.36 ;
      RECT  2.665 0.05 2.785 0.36 ;
      RECT  3.705 0.05 3.825 0.36 ;
      RECT  3.185 0.05 3.305 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.175 0.54 5.435 0.655 ;
      RECT  4.75 0.655 5.435 0.66 ;
      RECT  4.75 0.66 4.85 1.11 ;
      RECT  4.22 1.11 5.45 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.965 0.215 4.63 0.335 ;
      RECT  3.965 0.335 4.085 0.475 ;
      RECT  3.395 0.475 4.085 0.595 ;
      RECT  4.72 0.24 5.695 0.36 ;
      RECT  4.72 0.36 4.9 0.45 ;
      RECT  2.925 0.19 3.05 0.465 ;
      RECT  0.275 0.465 3.05 0.585 ;
      RECT  0.275 1.23 3.045 1.35 ;
      RECT  2.925 1.35 3.045 1.49 ;
      RECT  3.395 1.23 4.085 1.35 ;
      RECT  3.965 1.35 4.085 1.42 ;
      RECT  3.965 1.42 4.655 1.54 ;
      RECT  5.55 1.31 5.67 1.415 ;
      RECT  4.955 1.415 5.67 1.535 ;
      LAYER M2 ;
      RECT  2.91 0.35 4.9 0.45 ;
      RECT  2.9 1.35 5.69 1.45 ;
      LAYER V1 ;
      RECT  2.95 0.35 3.05 0.45 ;
      RECT  4.76 0.35 4.86 0.45 ;
      RECT  2.94 1.35 3.04 1.45 ;
      RECT  5.55 1.35 5.65 1.45 ;
  END
END SEN_MAJI3_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_T_4
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_T_4
  CLASS CORE ;
  FOREIGN SEN_MAJI3_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.785 ;
      RECT  1.75 0.785 4.165 0.895 ;
      RECT  1.75 0.895 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.715 0.745 6.305 0.895 ;
      RECT  0.35 0.71 1.05 0.89 ;
      LAYER M2 ;
      RECT  0.6 0.75 5.695 0.85 ;
      LAYER V1 ;
      RECT  4.845 0.75 4.945 0.85 ;
      RECT  5.2 0.75 5.3 0.85 ;
      RECT  5.555 0.75 5.655 0.85 ;
      RECT  0.64 0.75 0.74 0.85 ;
      RECT  0.84 0.75 0.94 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.65 0.895 ;
      RECT  7.55 0.895 7.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.445 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.845 1.44 0.965 1.75 ;
      RECT  2.655 1.44 2.775 1.75 ;
      RECT  3.175 1.44 3.295 1.75 ;
      RECT  3.695 1.44 3.815 1.75 ;
      RECT  4.215 1.44 4.335 1.75 ;
      RECT  4.735 1.44 4.855 1.75 ;
      RECT  5.255 1.44 5.375 1.75 ;
      RECT  5.775 1.44 5.895 1.75 ;
      RECT  6.295 1.44 6.415 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  2.655 0.05 2.775 0.425 ;
      RECT  3.175 0.05 3.295 0.425 ;
      RECT  3.695 0.05 3.815 0.425 ;
      RECT  4.215 0.05 4.335 0.425 ;
      RECT  4.735 0.05 4.855 0.425 ;
      RECT  5.255 0.05 5.375 0.425 ;
      RECT  5.775 0.05 5.895 0.425 ;
      RECT  6.295 0.05 6.415 0.425 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.79 0.47 7.505 0.59 ;
      RECT  6.95 0.59 7.05 1.05 ;
      RECT  2.15 1.05 7.05 1.105 ;
      RECT  2.15 1.105 7.45 1.14 ;
      RECT  2.15 1.14 2.25 1.205 ;
      RECT  6.815 1.14 7.45 1.29 ;
      RECT  1.34 0.47 2.055 0.59 ;
      RECT  1.55 0.59 1.65 1.11 ;
      RECT  1.345 1.11 1.65 1.205 ;
      RECT  1.345 1.205 2.25 1.315 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.555 0.215 7.715 0.335 ;
      RECT  7.595 0.335 7.715 0.445 ;
      RECT  6.555 0.335 6.675 0.515 ;
      RECT  2.395 0.425 2.515 0.515 ;
      RECT  2.395 0.515 6.675 0.635 ;
      RECT  1.105 0.22 2.315 0.34 ;
      RECT  1.105 0.34 1.225 0.475 ;
      RECT  0.065 0.29 0.185 0.475 ;
      RECT  0.065 0.475 1.225 0.595 ;
      RECT  0.065 1.225 1.225 1.35 ;
      RECT  1.105 1.35 1.225 1.43 ;
      RECT  0.065 1.35 0.185 1.435 ;
      RECT  1.105 1.43 2.305 1.55 ;
      RECT  2.395 1.23 6.675 1.35 ;
      RECT  6.555 1.35 6.675 1.43 ;
      RECT  2.395 1.35 2.515 1.46 ;
      RECT  6.555 1.43 7.715 1.55 ;
      RECT  7.595 1.325 7.715 1.43 ;
  END
END SEN_MAJI3_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_T_6
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_T_6
  CLASS CORE ;
  FOREIGN SEN_MAJI3_T_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 0.785 ;
      RECT  2.52 0.785 6.43 0.895 ;
      RECT  2.52 0.895 2.865 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1664 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.665 0.71 9.13 0.89 ;
      RECT  0.55 0.71 1.49 0.89 ;
      LAYER M2 ;
      RECT  1.11 0.75 7.83 0.85 ;
      LAYER V1 ;
      RECT  6.73 0.75 6.83 0.85 ;
      RECT  6.93 0.75 7.03 0.85 ;
      RECT  7.31 0.75 7.41 0.85 ;
      RECT  7.69 0.75 7.79 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1664 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.245 0.71 11.05 0.89 ;
      RECT  10.95 0.89 11.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.445 1.75 ;
      RECT  0.0 1.75 11.4 1.85 ;
      RECT  0.845 1.44 0.965 1.75 ;
      RECT  1.365 1.44 1.485 1.75 ;
      RECT  3.675 1.44 3.795 1.75 ;
      RECT  4.195 1.44 4.315 1.75 ;
      RECT  4.715 1.44 4.835 1.75 ;
      RECT  5.235 1.44 5.355 1.75 ;
      RECT  5.755 1.44 5.875 1.75 ;
      RECT  6.275 1.44 6.395 1.75 ;
      RECT  6.795 1.44 6.915 1.75 ;
      RECT  7.315 1.44 7.435 1.75 ;
      RECT  7.835 1.44 7.955 1.75 ;
      RECT  8.355 1.44 8.475 1.75 ;
      RECT  8.875 1.44 8.995 1.75 ;
      RECT  9.395 1.44 9.515 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.4 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  3.675 0.05 3.795 0.36 ;
      RECT  4.195 0.05 4.315 0.36 ;
      RECT  4.715 0.05 4.835 0.36 ;
      RECT  5.235 0.05 5.355 0.36 ;
      RECT  5.755 0.05 5.875 0.36 ;
      RECT  6.275 0.05 6.395 0.36 ;
      RECT  6.795 0.05 6.915 0.36 ;
      RECT  7.315 0.05 7.435 0.36 ;
      RECT  7.835 0.05 7.955 0.36 ;
      RECT  8.355 0.05 8.475 0.36 ;
      RECT  8.875 0.05 8.995 0.36 ;
      RECT  9.395 0.05 9.515 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.89 0.475 11.125 0.595 ;
      RECT  9.95 0.595 10.08 0.91 ;
      RECT  9.34 0.91 10.08 1.0 ;
      RECT  3.15 1.0 10.08 1.09 ;
      RECT  9.91 1.09 10.08 1.11 ;
      RECT  3.15 1.09 9.445 1.13 ;
      RECT  9.91 1.11 10.65 1.205 ;
      RECT  3.15 1.13 3.28 1.22 ;
      RECT  9.91 1.205 11.125 1.31 ;
      RECT  1.885 0.51 3.05 0.69 ;
      RECT  2.15 0.69 2.28 1.22 ;
      RECT  1.86 1.22 3.28 1.35 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.625 0.205 3.355 0.335 ;
      RECT  1.625 0.335 1.755 0.465 ;
      RECT  0.065 0.29 0.185 0.465 ;
      RECT  0.065 0.465 1.755 0.595 ;
      RECT  9.65 0.21 11.335 0.34 ;
      RECT  11.215 0.34 11.335 0.405 ;
      RECT  9.65 0.34 9.78 0.45 ;
      RECT  3.39 0.45 9.78 0.58 ;
      RECT  0.065 1.22 1.75 1.35 ;
      RECT  1.62 1.35 1.75 1.46 ;
      RECT  0.065 1.35 0.185 1.51 ;
      RECT  1.62 1.46 3.355 1.59 ;
      RECT  3.37 1.22 9.78 1.35 ;
      RECT  9.65 1.35 9.78 1.425 ;
      RECT  9.65 1.425 11.335 1.555 ;
      RECT  11.215 1.29 11.335 1.425 ;
  END
END SEN_MAJI3_T_6
#-----------------------------------------------------------------------
#      Cell        : SEN_MAJI3_T_8
#      Description : "3-input majority, inverted"
#      Equation    : X=!((A1&A2)|(A1&A3)|(A2&A3))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MAJI3_T_8
  CLASS CORE ;
  FOREIGN SEN_MAJI3_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 15.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.45 0.755 ;
      RECT  3.27 0.755 8.86 0.845 ;
      RECT  3.27 0.845 3.65 0.85 ;
      RECT  3.335 0.85 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5552 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.115 0.75 13.13 0.85 ;
      RECT  0.66 0.71 1.855 0.89 ;
      LAYER M2 ;
      RECT  1.31 0.75 10.855 0.85 ;
      LAYER V1 ;
      RECT  9.35 0.75 9.45 0.85 ;
      RECT  9.68 0.75 9.78 0.85 ;
      RECT  10.01 0.75 10.11 0.85 ;
      RECT  10.34 0.75 10.44 0.85 ;
      RECT  10.67 0.75 10.77 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5552 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  13.67 0.71 14.85 0.89 ;
      RECT  14.75 0.89 14.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 15.2 1.85 ;
      RECT  0.845 1.415 0.965 1.75 ;
      RECT  1.365 1.415 1.48 1.75 ;
      RECT  1.885 1.415 2.005 1.75 ;
      RECT  4.845 1.48 5.015 1.75 ;
      RECT  5.365 1.48 5.535 1.75 ;
      RECT  5.885 1.48 6.055 1.75 ;
      RECT  6.405 1.48 6.575 1.75 ;
      RECT  6.925 1.48 7.095 1.75 ;
      RECT  7.445 1.48 7.615 1.75 ;
      RECT  7.965 1.48 8.135 1.75 ;
      RECT  8.485 1.48 8.655 1.75 ;
      RECT  9.005 1.48 9.175 1.75 ;
      RECT  9.525 1.48 9.695 1.75 ;
      RECT  10.045 1.48 10.215 1.75 ;
      RECT  10.565 1.48 10.735 1.75 ;
      RECT  11.085 1.48 11.255 1.75 ;
      RECT  11.605 1.48 11.775 1.75 ;
      RECT  12.125 1.48 12.295 1.75 ;
      RECT  12.645 1.48 12.815 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 15.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
      RECT  14.65 1.75 14.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 15.2 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  1.885 0.05 2.005 0.36 ;
      RECT  4.825 0.05 4.945 0.36 ;
      RECT  5.345 0.05 5.465 0.36 ;
      RECT  5.865 0.05 5.985 0.36 ;
      RECT  6.385 0.05 6.505 0.36 ;
      RECT  6.905 0.05 7.025 0.36 ;
      RECT  7.425 0.05 7.545 0.36 ;
      RECT  7.945 0.05 8.065 0.36 ;
      RECT  8.465 0.05 8.585 0.36 ;
      RECT  9.03 0.05 9.15 0.36 ;
      RECT  9.55 0.05 9.67 0.36 ;
      RECT  10.07 0.05 10.19 0.36 ;
      RECT  10.59 0.05 10.71 0.36 ;
      RECT  11.11 0.05 11.23 0.36 ;
      RECT  11.63 0.05 11.75 0.36 ;
      RECT  12.15 0.05 12.27 0.36 ;
      RECT  12.67 0.05 12.79 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 15.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
      RECT  14.65 -0.05 14.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  13.165 0.465 14.92 0.595 ;
      RECT  13.28 0.595 13.45 0.94 ;
      RECT  4.15 0.94 13.45 1.11 ;
      RECT  4.15 1.11 4.32 1.205 ;
      RECT  13.19 1.11 14.65 1.205 ;
      RECT  2.38 0.45 4.11 0.57 ;
      RECT  2.945 0.57 3.115 1.11 ;
      RECT  2.405 1.11 3.115 1.205 ;
      RECT  2.405 1.205 4.32 1.29 ;
      RECT  13.19 1.205 14.92 1.305 ;
      RECT  2.945 1.29 4.32 1.375 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.1 0.205 4.395 0.345 ;
      RECT  2.1 0.345 2.24 0.465 ;
      RECT  0.065 0.41 0.185 0.465 ;
      RECT  0.065 0.465 2.24 0.605 ;
      RECT  12.905 0.19 15.115 0.36 ;
      RECT  12.905 0.36 13.075 0.45 ;
      RECT  4.565 0.45 13.075 0.62 ;
      RECT  0.065 1.17 2.27 1.31 ;
      RECT  0.065 1.31 0.185 1.365 ;
      RECT  2.13 1.31 2.27 1.465 ;
      RECT  2.13 1.465 4.395 1.605 ;
      RECT  4.53 1.205 13.075 1.375 ;
      RECT  12.905 1.375 13.075 1.44 ;
      RECT  12.905 1.44 15.13 1.61 ;
  END
END SEN_MAJI3_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_0P5
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_0P5
  CLASS CORE ;
  FOREIGN SEN_MUX2_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.705 1.66 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0399 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.41 1.495 0.58 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.705 1.39 1.835 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.42 0.05 0.55 0.39 ;
      RECT  1.74 0.05 1.86 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.265 2.12 0.45 ;
      RECT  1.95 0.45 2.05 1.39 ;
      RECT  1.95 1.39 2.12 1.56 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.11 0.14 1.65 0.23 ;
      RECT  1.56 0.23 1.65 0.505 ;
      RECT  1.11 0.23 1.215 1.46 ;
      RECT  1.56 0.505 1.85 0.595 ;
      RECT  1.75 0.595 1.85 0.91 ;
      RECT  1.355 0.32 1.47 0.535 ;
      RECT  1.355 0.535 1.46 1.46 ;
      RECT  0.74 0.19 0.84 1.225 ;
      RECT  0.14 0.18 0.26 1.315 ;
      RECT  0.14 1.315 1.02 1.405 ;
      RECT  0.93 0.515 1.02 1.315 ;
      RECT  0.93 1.405 1.02 1.55 ;
      RECT  0.93 1.55 1.375 1.66 ;
  END
END SEN_MUX2_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_1
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_1
  CLASS CORE ;
  FOREIGN SEN_MUX2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.46 0.725 0.56 0.91 ;
      RECT  0.35 0.91 0.56 1.0 ;
      RECT  0.35 1.0 0.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.65 0.73 ;
      RECT  1.55 0.73 1.67 0.925 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.063 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.68 0.16 1.28 0.25 ;
      RECT  0.68 0.25 0.78 0.26 ;
      RECT  1.19 0.25 1.28 0.82 ;
      RECT  0.26 0.26 0.78 0.35 ;
      RECT  0.26 0.35 0.36 0.62 ;
      RECT  0.235 0.62 0.36 0.79 ;
      LAYER M2 ;
      RECT  0.21 0.35 0.775 0.45 ;
      LAYER V1 ;
      RECT  0.26 0.35 0.36 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0828 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.575 0.485 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.745 1.44 1.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.32 0.05 0.49 0.17 ;
      RECT  1.745 0.05 1.86 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.13 0.69 ;
      RECT  2.025 0.69 2.13 1.11 ;
      RECT  1.95 1.11 2.13 1.2 ;
      RECT  1.95 1.2 2.05 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.37 0.17 0.54 ;
      RECT  0.055 0.54 0.145 1.395 ;
      RECT  0.055 1.395 0.92 1.485 ;
      RECT  0.83 0.715 0.92 1.395 ;
      RECT  0.83 1.485 0.92 1.555 ;
      RECT  0.055 1.485 0.175 1.59 ;
      RECT  0.83 1.555 1.51 1.655 ;
      RECT  0.65 0.44 0.85 0.55 ;
      RECT  0.65 0.55 0.74 1.21 ;
      RECT  1.76 0.78 1.935 0.95 ;
      RECT  1.76 0.95 1.86 1.24 ;
      RECT  0.95 0.34 1.05 0.525 ;
      RECT  0.95 0.525 1.1 0.615 ;
      RECT  1.01 0.615 1.1 1.24 ;
      RECT  1.01 1.24 1.86 1.35 ;
      RECT  1.37 0.37 1.46 1.04 ;
      RECT  1.37 1.04 1.65 1.15 ;
  END
END SEN_MUX2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_2
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_2
  CLASS CORE ;
  FOREIGN SEN_MUX2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.93 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 2.85 1.185 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.665 0.45 1.02 ;
      RECT  0.35 1.02 1.685 1.03 ;
      RECT  0.985 0.925 1.685 1.02 ;
      RECT  0.35 1.03 1.075 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1656 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.385 1.59 0.555 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  1.035 1.59 1.205 1.75 ;
      RECT  2.635 1.46 2.805 1.75 ;
      RECT  3.215 1.46 3.385 1.75 ;
      RECT  3.805 1.215 3.925 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.6 0.05 0.73 0.39 ;
      RECT  3.795 0.05 3.93 0.39 ;
      RECT  2.7 0.05 2.815 0.44 ;
      RECT  1.135 0.05 1.255 0.59 ;
      RECT  3.235 0.05 3.355 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.495 0.51 3.85 0.69 ;
      RECT  3.75 0.69 3.85 1.005 ;
      RECT  3.53 1.005 3.85 1.125 ;
      RECT  3.53 1.125 3.65 1.3 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.145 0.325 2.325 0.4 ;
      RECT  1.885 0.4 2.325 0.415 ;
      RECT  1.885 0.415 2.235 0.49 ;
      RECT  1.885 0.49 1.975 0.74 ;
      RECT  0.83 0.28 1.04 0.4 ;
      RECT  0.95 0.4 1.04 0.74 ;
      RECT  0.95 0.74 1.975 0.83 ;
      RECT  1.775 0.83 1.865 1.2 ;
      RECT  0.735 1.2 1.865 1.3 ;
      RECT  1.615 0.405 1.795 0.65 ;
      RECT  3.265 0.78 3.64 0.88 ;
      RECT  3.265 0.88 3.355 1.28 ;
      RECT  1.955 0.14 2.55 0.2 ;
      RECT  1.39 0.2 2.55 0.23 ;
      RECT  1.39 0.23 2.055 0.31 ;
      RECT  2.43 0.23 2.55 0.33 ;
      RECT  1.39 0.31 1.51 0.42 ;
      RECT  2.43 0.33 2.605 0.42 ;
      RECT  2.515 0.42 2.605 1.28 ;
      RECT  2.41 1.28 3.355 1.37 ;
      RECT  2.41 1.37 2.53 1.57 ;
      RECT  1.295 1.57 2.53 1.66 ;
      RECT  2.11 0.725 2.21 0.92 ;
      RECT  1.955 0.92 2.21 1.01 ;
      RECT  1.955 1.01 2.045 1.39 ;
      RECT  0.34 0.26 0.47 0.48 ;
      RECT  0.065 0.48 0.47 0.575 ;
      RECT  0.065 0.575 0.185 1.39 ;
      RECT  0.065 1.39 2.045 1.48 ;
      RECT  2.325 0.51 2.425 1.1 ;
      RECT  2.14 1.1 2.425 1.19 ;
      RECT  2.14 1.19 2.26 1.43 ;
      RECT  2.95 0.44 3.07 1.15 ;
      LAYER M2 ;
      RECT  1.615 0.55 3.105 0.65 ;
      LAYER V1 ;
      RECT  1.655 0.55 1.755 0.65 ;
      RECT  2.325 0.55 2.425 0.65 ;
      RECT  2.965 0.55 3.065 0.65 ;
  END
END SEN_MUX2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_3
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_3
  CLASS CORE ;
  FOREIGN SEN_MUX2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.79 1.115 0.91 ;
      RECT  0.55 0.91 1.115 1.09 ;
      RECT  0.55 1.09 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.189 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 3.92 0.89 ;
      RECT  3.55 0.89 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.189 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.605 1.45 0.695 ;
      RECT  0.55 0.695 0.65 0.7 ;
      RECT  1.35 0.695 1.45 0.76 ;
      RECT  0.35 0.7 0.65 0.795 ;
      RECT  1.35 0.76 2.035 0.89 ;
      RECT  0.35 0.795 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2484 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.57 1.585 0.74 1.75 ;
      RECT  1.11 1.585 1.28 1.75 ;
      RECT  3.635 1.59 3.805 1.75 ;
      RECT  4.2 1.495 4.37 1.75 ;
      RECT  4.74 1.215 4.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  1.08 0.05 1.25 0.315 ;
      RECT  0.06 0.05 0.185 0.365 ;
      RECT  4.74 0.05 4.87 0.385 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  3.68 0.05 3.81 0.4 ;
      RECT  4.215 0.05 4.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.46 0.51 5.125 0.69 ;
      RECT  4.95 0.69 5.125 1.0 ;
      RECT  4.46 1.0 5.125 1.12 ;
      RECT  4.95 1.12 5.125 1.49 ;
    END
    ANTENNADIFFAREA 0.4 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.59 0.18 3.545 0.27 ;
      RECT  2.09 0.27 2.28 0.305 ;
      RECT  1.59 0.27 1.775 0.325 ;
      RECT  3.425 0.27 3.545 0.49 ;
      RECT  3.425 0.49 4.1 0.595 ;
      RECT  4.01 0.595 4.1 1.04 ;
      RECT  3.75 1.04 4.1 1.16 ;
      RECT  3.75 1.16 3.85 1.18 ;
      RECT  2.75 1.18 3.85 1.29 ;
      RECT  0.82 0.415 1.76 0.515 ;
      RECT  1.66 0.515 1.76 0.58 ;
      RECT  1.66 0.58 2.845 0.67 ;
      RECT  2.62 0.54 2.845 0.58 ;
      RECT  2.135 0.67 2.225 1.015 ;
      RECT  1.4 1.015 2.225 1.105 ;
      RECT  1.4 1.105 1.51 1.21 ;
      RECT  0.81 1.21 1.51 1.3 ;
      RECT  2.315 0.78 2.89 0.87 ;
      RECT  2.315 0.87 2.405 1.2 ;
      RECT  1.6 1.2 2.405 1.29 ;
      RECT  1.6 1.29 1.7 1.405 ;
      RECT  0.155 0.455 0.47 0.555 ;
      RECT  0.155 0.555 0.255 1.21 ;
      RECT  0.155 1.21 0.445 1.3 ;
      RECT  0.325 1.3 0.445 1.405 ;
      RECT  0.325 1.405 1.7 1.495 ;
      RECT  4.25 0.795 4.81 0.885 ;
      RECT  4.25 0.885 4.35 1.31 ;
      RECT  3.95 1.31 4.35 1.4 ;
      RECT  2.37 0.36 3.09 0.4 ;
      RECT  1.85 0.4 3.09 0.45 ;
      RECT  1.85 0.45 2.545 0.49 ;
      RECT  2.98 0.45 3.09 0.98 ;
      RECT  2.495 0.98 3.09 1.07 ;
      RECT  2.495 1.07 2.61 1.4 ;
      RECT  1.79 1.4 4.05 1.5 ;
      RECT  1.79 1.5 1.905 1.62 ;
      RECT  3.18 0.405 3.29 0.92 ;
      LAYER M2 ;
      RECT  2.635 0.55 3.33 0.65 ;
      LAYER V1 ;
      RECT  2.675 0.55 2.775 0.65 ;
      RECT  3.19 0.55 3.29 0.65 ;
  END
END SEN_MUX2_3
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_4
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_4
  CLASS CORE ;
  FOREIGN SEN_MUX2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.02 0.78 1.4 0.905 ;
      RECT  1.02 0.905 1.25 0.91 ;
      RECT  0.55 0.91 1.25 1.09 ;
      RECT  0.55 1.09 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.65 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.785 0.6 1.58 0.69 ;
      RECT  0.785 0.69 0.875 0.71 ;
      RECT  1.49 0.69 1.58 0.8 ;
      RECT  0.35 0.71 0.875 0.8 ;
      RECT  0.35 0.8 0.45 1.09 ;
      RECT  1.49 0.8 2.44 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3285 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.57 1.59 0.74 1.75 ;
      RECT  1.11 1.59 1.28 1.75 ;
      RECT  1.65 1.59 1.82 1.75 ;
      RECT  3.845 1.585 4.015 1.75 ;
      RECT  4.385 1.585 4.555 1.75 ;
      RECT  4.97 1.41 5.1 1.75 ;
      RECT  5.495 1.21 5.615 1.75 ;
      RECT  6.015 1.21 6.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  3.85 0.05 4.02 0.215 ;
      RECT  1.355 0.05 1.525 0.31 ;
      RECT  4.45 0.05 4.58 0.38 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  5.49 0.05 5.62 0.39 ;
      RECT  1.9 0.05 2.02 0.42 ;
      RECT  0.825 0.05 0.995 0.505 ;
      RECT  4.975 0.05 5.095 0.59 ;
      RECT  6.015 0.05 6.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.21 0.51 5.87 0.69 ;
      RECT  5.75 0.69 5.87 1.0 ;
      RECT  5.21 1.0 5.87 1.12 ;
      RECT  5.75 1.12 5.87 1.49 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.135 0.18 3.76 0.27 ;
      RECT  2.135 0.27 2.795 0.305 ;
      RECT  3.67 0.27 3.76 0.31 ;
      RECT  2.135 0.305 2.25 0.48 ;
      RECT  3.67 0.31 4.11 0.4 ;
      RECT  4.01 0.4 4.11 0.47 ;
      RECT  4.01 0.47 4.86 0.59 ;
      RECT  4.75 0.59 4.86 1.01 ;
      RECT  4.55 1.01 4.86 1.125 ;
      RECT  4.55 1.125 4.65 1.2 ;
      RECT  3.095 1.2 4.65 1.29 ;
      RECT  1.095 0.4 1.785 0.49 ;
      RECT  1.69 0.49 1.785 0.6 ;
      RECT  1.69 0.6 3.335 0.69 ;
      RECT  3.08 0.55 3.335 0.6 ;
      RECT  2.53 0.69 2.63 1.015 ;
      RECT  1.75 1.015 2.63 1.105 ;
      RECT  1.75 1.105 1.85 1.205 ;
      RECT  0.81 1.205 1.85 1.305 ;
      RECT  3.685 0.49 3.815 0.87 ;
      RECT  5.0 0.795 5.64 0.885 ;
      RECT  5.0 0.885 5.09 1.215 ;
      RECT  4.75 1.215 5.09 1.305 ;
      RECT  4.75 1.305 4.85 1.4 ;
      RECT  3.42 1.4 4.85 1.45 ;
      RECT  2.885 0.36 3.575 0.4 ;
      RECT  2.365 0.4 3.575 0.45 ;
      RECT  2.365 0.45 3.0 0.49 ;
      RECT  3.48 0.45 3.575 1.0 ;
      RECT  2.91 1.0 3.575 1.09 ;
      RECT  2.91 1.09 3.005 1.45 ;
      RECT  2.155 1.45 4.85 1.49 ;
      RECT  2.155 1.49 3.56 1.57 ;
      RECT  2.72 0.8 3.39 0.89 ;
      RECT  2.72 0.89 2.82 1.2 ;
      RECT  1.95 1.2 2.82 1.29 ;
      RECT  1.95 1.29 2.05 1.405 ;
      RECT  0.065 0.36 0.185 0.495 ;
      RECT  0.065 0.495 0.695 0.59 ;
      RECT  0.585 0.36 0.695 0.495 ;
      RECT  0.115 0.59 0.225 1.21 ;
      RECT  0.115 1.21 0.45 1.3 ;
      RECT  0.315 1.3 0.45 1.405 ;
      RECT  0.315 1.405 2.05 1.5 ;
      LAYER M2 ;
      RECT  3.105 0.55 3.85 0.65 ;
      LAYER V1 ;
      RECT  3.15 0.55 3.25 0.65 ;
      RECT  3.7 0.55 3.8 0.65 ;
  END
END SEN_MUX2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_6
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_6
  CLASS CORE ;
  FOREIGN SEN_MUX2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.51 5.85 0.71 ;
      RECT  4.775 0.71 5.85 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2727 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.85 0.91 ;
      RECT  6.75 0.91 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2727 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.79 0.745 4.215 0.895 ;
      RECT  1.915 0.71 2.285 0.89 ;
      LAYER M2 ;
      RECT  1.91 0.75 3.97 0.85 ;
      LAYER V1 ;
      RECT  3.83 0.75 3.93 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3501 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.6 1.49 1.77 1.75 ;
      RECT  2.12 1.49 2.29 1.75 ;
      RECT  4.645 1.47 4.815 1.75 ;
      RECT  5.165 1.47 5.335 1.75 ;
      RECT  5.685 1.47 5.855 1.75 ;
      RECT  6.205 1.47 6.375 1.75 ;
      RECT  6.725 1.47 6.895 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  4.625 0.05 4.755 0.255 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  1.62 0.05 1.75 0.39 ;
      RECT  5.185 0.05 5.315 0.39 ;
      RECT  5.705 0.05 5.835 0.39 ;
      RECT  6.225 0.05 6.355 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.77 0.05 6.89 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.325 0.51 1.65 0.69 ;
      RECT  0.55 0.69 0.68 1.11 ;
      RECT  0.325 1.11 1.525 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.205 0.14 4.45 0.23 ;
      RECT  3.205 0.23 3.325 0.275 ;
      RECT  4.36 0.23 4.45 0.345 ;
      RECT  2.635 0.275 3.325 0.4 ;
      RECT  4.36 0.345 4.67 0.435 ;
      RECT  4.58 0.435 4.67 0.48 ;
      RECT  4.58 0.48 5.62 0.6 ;
      RECT  4.58 0.6 4.67 1.005 ;
      RECT  3.775 1.005 4.67 1.075 ;
      RECT  3.775 1.075 5.62 1.11 ;
      RECT  4.555 1.11 5.62 1.195 ;
      RECT  3.415 0.32 4.23 0.44 ;
      RECT  3.415 0.44 3.505 0.49 ;
      RECT  2.895 0.49 3.505 0.61 ;
      RECT  3.415 0.61 3.505 1.145 ;
      RECT  2.695 1.145 3.505 1.265 ;
      RECT  2.695 1.265 2.785 1.31 ;
      RECT  3.415 1.265 3.505 1.38 ;
      RECT  0.825 0.785 1.725 0.895 ;
      RECT  1.635 0.895 1.725 1.31 ;
      RECT  1.635 1.31 2.785 1.4 ;
      RECT  3.415 1.38 4.23 1.48 ;
      RECT  1.835 0.45 2.55 0.57 ;
      RECT  2.46 0.57 2.55 0.78 ;
      RECT  2.46 0.78 3.325 0.9 ;
      RECT  2.46 0.9 2.55 1.115 ;
      RECT  1.835 1.115 2.55 1.22 ;
      RECT  5.945 0.485 6.66 0.605 ;
      RECT  5.945 0.605 6.055 1.255 ;
      RECT  5.945 1.255 7.13 1.285 ;
      RECT  3.595 0.53 4.49 0.65 ;
      RECT  3.595 0.65 3.685 1.2 ;
      RECT  3.595 1.2 4.43 1.285 ;
      RECT  3.595 1.285 7.13 1.29 ;
      RECT  4.335 1.29 7.13 1.375 ;
      RECT  7.01 1.375 7.13 1.475 ;
      RECT  4.335 1.375 4.43 1.57 ;
      RECT  3.205 1.39 3.325 1.49 ;
      RECT  2.635 1.49 3.325 1.57 ;
      RECT  2.635 1.57 4.43 1.6 ;
      RECT  3.205 1.6 4.43 1.66 ;
  END
END SEN_MUX2_6
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_8
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_8
  CLASS CORE ;
  FOREIGN SEN_MUX2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.51 7.45 0.71 ;
      RECT  6.35 0.71 7.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3636 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.71 8.65 0.89 ;
      RECT  7.95 0.89 8.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3636 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.71 5.65 0.785 ;
      RECT  4.87 0.785 5.65 0.895 ;
      RECT  2.55 0.71 3.05 0.89 ;
      LAYER M2 ;
      RECT  2.71 0.75 5.69 0.85 ;
      LAYER V1 ;
      RECT  5.55 0.75 5.65 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.462 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.2 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.12 1.49 2.29 1.75 ;
      RECT  2.64 1.49 2.81 1.75 ;
      RECT  3.16 1.49 3.33 1.75 ;
      RECT  5.79 1.44 5.92 1.75 ;
      RECT  6.33 1.44 6.46 1.75 ;
      RECT  6.85 1.44 6.98 1.75 ;
      RECT  7.37 1.44 7.5 1.75 ;
      RECT  7.89 1.44 8.02 1.75 ;
      RECT  8.41 1.44 8.54 1.75 ;
      RECT  8.96 1.21 9.08 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.2 0.05 ;
      RECT  5.795 0.05 5.92 0.29 ;
      RECT  2.64 0.05 2.81 0.35 ;
      RECT  3.16 0.05 3.33 0.35 ;
      RECT  6.33 0.05 6.46 0.385 ;
      RECT  6.85 0.05 6.98 0.385 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  1.62 0.05 1.75 0.39 ;
      RECT  2.14 0.05 2.27 0.39 ;
      RECT  7.37 0.05 7.5 0.39 ;
      RECT  7.89 0.05 8.02 0.39 ;
      RECT  8.41 0.05 8.54 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  8.96 0.05 9.08 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.3 0.51 2.05 0.69 ;
      RECT  0.55 0.69 0.72 1.11 ;
      RECT  0.325 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.45 0.2 5.7 0.305 ;
      RECT  3.45 0.305 3.57 0.575 ;
      RECT  3.45 0.575 4.415 0.665 ;
      RECT  4.325 0.665 4.415 1.04 ;
      RECT  3.45 1.04 4.415 1.135 ;
      RECT  3.45 1.135 3.57 1.31 ;
      RECT  0.83 0.785 2.245 0.895 ;
      RECT  2.155 0.895 2.245 1.31 ;
      RECT  2.155 1.31 3.57 1.4 ;
      RECT  3.45 1.4 3.57 1.45 ;
      RECT  3.45 1.45 5.7 1.57 ;
      RECT  3.66 0.395 6.0 0.475 ;
      RECT  3.66 0.475 7.26 0.485 ;
      RECT  5.87 0.485 7.26 0.605 ;
      RECT  5.87 0.605 6.0 1.02 ;
      RECT  4.7 1.02 7.285 1.14 ;
      RECT  2.355 0.44 3.245 0.56 ;
      RECT  3.155 0.56 3.245 0.78 ;
      RECT  3.155 0.78 4.235 0.9 ;
      RECT  3.155 0.9 3.245 1.115 ;
      RECT  2.355 1.115 3.245 1.22 ;
      RECT  7.61 0.485 8.845 0.605 ;
      RECT  7.61 0.605 7.74 1.23 ;
      RECT  4.515 0.575 5.44 0.665 ;
      RECT  4.515 0.665 4.605 1.23 ;
      RECT  3.66 1.23 8.845 1.35 ;
  END
END SEN_MUX2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_DG_1
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_DG_1
  CLASS CORE ;
  FOREIGN SEN_MUX2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.71 0.65 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.7 1.25 0.83 ;
      RECT  1.15 0.83 1.3 1.01 ;
      RECT  1.15 1.01 1.25 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.165 1.14 0.255 ;
      RECT  0.55 0.255 0.65 0.5 ;
      RECT  0.35 0.5 0.65 0.59 ;
      RECT  0.35 0.59 0.45 0.91 ;
      RECT  0.26 0.91 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.46 0.46 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.35 1.21 1.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.345 0.05 1.475 0.36 ;
      RECT  0.33 0.05 0.46 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.61 0.34 1.73 1.11 ;
      RECT  1.55 1.11 1.73 1.2 ;
      RECT  1.55 1.2 1.65 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.835 0.45 1.52 0.54 ;
      RECT  1.43 0.54 1.52 0.93 ;
      RECT  0.835 0.54 0.925 1.405 ;
      RECT  0.065 0.335 0.17 1.28 ;
      RECT  0.065 1.28 0.665 1.37 ;
      RECT  0.575 1.37 0.665 1.565 ;
      RECT  0.575 1.565 1.1 1.66 ;
  END
END SEN_MUX2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_DG_12
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_DG_12
  CLASS CORE ;
  FOREIGN SEN_MUX2_DG_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.45 0.71 ;
      RECT  2.95 0.71 3.45 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.335 0.89 ;
      RECT  3.95 0.89 4.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.31 0.975 ;
      RECT  0.52 0.75 0.84 0.94 ;
      LAYER M2 ;
      RECT  0.66 0.75 2.29 0.85 ;
      LAYER V1 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  0.7 0.75 0.8 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2904 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.585 1.21 0.705 1.75 ;
      RECT  2.9 1.44 3.03 1.75 ;
      RECT  3.42 1.44 3.55 1.75 ;
      RECT  3.93 1.44 4.06 1.75 ;
      RECT  4.45 1.41 4.58 1.75 ;
      RECT  4.97 1.41 5.1 1.75 ;
      RECT  5.49 1.41 5.62 1.75 ;
      RECT  6.01 1.41 6.14 1.75 ;
      RECT  6.53 1.41 6.66 1.75 ;
      RECT  7.05 1.41 7.18 1.75 ;
      RECT  7.59 1.205 7.71 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  4.97 0.05 5.1 0.35 ;
      RECT  5.49 0.05 5.62 0.35 ;
      RECT  6.01 0.05 6.14 0.35 ;
      RECT  6.53 0.05 6.66 0.35 ;
      RECT  7.05 0.05 7.18 0.35 ;
      RECT  3.93 0.05 4.06 0.36 ;
      RECT  3.425 0.05 3.55 0.39 ;
      RECT  0.58 0.05 0.71 0.43 ;
      RECT  2.9 0.05 3.03 0.43 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  4.455 0.05 4.575 0.59 ;
      RECT  7.59 0.05 7.71 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.665 0.44 7.485 0.56 ;
      RECT  5.73 0.56 6.86 0.61 ;
      RECT  6.61 0.61 6.86 1.11 ;
      RECT  4.73 1.11 7.45 1.29 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.12 0.24 3.335 0.36 ;
      RECT  3.12 0.36 3.21 0.52 ;
      RECT  0.835 0.14 2.765 0.23 ;
      RECT  1.355 0.23 1.475 0.39 ;
      RECT  0.835 0.23 0.955 0.43 ;
      RECT  2.645 0.23 2.765 0.52 ;
      RECT  2.645 0.52 3.21 0.61 ;
      RECT  2.645 0.61 2.75 1.025 ;
      RECT  2.645 1.025 3.335 1.055 ;
      RECT  2.41 1.055 3.335 1.145 ;
      RECT  2.41 1.145 2.5 1.36 ;
      RECT  1.825 1.36 2.5 1.48 ;
      RECT  1.615 0.32 2.305 0.41 ;
      RECT  1.615 0.41 1.735 0.48 ;
      RECT  1.11 0.33 1.215 0.48 ;
      RECT  1.11 0.48 1.735 0.57 ;
      RECT  1.19 0.57 1.28 1.11 ;
      RECT  1.095 1.11 1.28 1.29 ;
      RECT  0.325 0.29 0.445 0.53 ;
      RECT  0.325 0.53 1.02 0.62 ;
      RECT  0.93 0.62 1.02 0.955 ;
      RECT  0.325 0.62 0.43 1.45 ;
      RECT  3.65 0.455 4.365 0.575 ;
      RECT  3.65 0.575 3.74 1.255 ;
      RECT  2.72 1.255 4.365 1.345 ;
      RECT  2.72 1.345 2.81 1.57 ;
      RECT  2.41 0.35 2.515 0.5 ;
      RECT  1.85 0.5 2.515 0.59 ;
      RECT  1.85 0.59 1.94 0.885 ;
      RECT  1.37 0.885 1.94 0.975 ;
      RECT  1.37 0.975 1.46 1.57 ;
      RECT  0.83 1.37 0.955 1.57 ;
      RECT  0.83 1.57 2.81 1.66 ;
      RECT  4.53 0.77 6.52 0.895 ;
      RECT  4.53 0.895 4.63 1.31 ;
      RECT  1.565 1.115 2.28 1.205 ;
      RECT  2.1 1.205 2.28 1.25 ;
      LAYER M2 ;
      RECT  1.14 1.15 4.67 1.25 ;
      LAYER V1 ;
      RECT  1.18 1.15 1.28 1.25 ;
      RECT  2.14 1.15 2.24 1.25 ;
      RECT  4.53 1.15 4.63 1.25 ;
  END
END SEN_MUX2_DG_12
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_DG_16
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_DG_16
  CLASS CORE ;
  FOREIGN SEN_MUX2_DG_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.45 0.71 ;
      RECT  3.75 0.71 4.45 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.84 0.71 5.25 0.89 ;
      RECT  5.15 0.89 5.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.21 0.71 2.65 0.89 ;
      RECT  0.52 0.71 0.84 0.89 ;
      LAYER M2 ;
      RECT  0.7 0.75 2.35 0.85 ;
      LAYER V1 ;
      RECT  2.21 0.75 2.31 0.85 ;
      RECT  0.74 0.75 0.84 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  0.585 1.21 0.705 1.75 ;
      RECT  3.29 1.44 3.4 1.75 ;
      RECT  3.79 1.44 3.92 1.75 ;
      RECT  4.31 1.44 4.44 1.75 ;
      RECT  4.83 1.44 4.96 1.75 ;
      RECT  5.35 1.41 5.48 1.75 ;
      RECT  5.87 1.41 6.0 1.75 ;
      RECT  6.39 1.41 6.52 1.75 ;
      RECT  6.91 1.41 7.04 1.75 ;
      RECT  7.445 1.41 7.575 1.75 ;
      RECT  7.975 1.41 8.105 1.75 ;
      RECT  8.495 1.41 8.625 1.75 ;
      RECT  9.015 1.41 9.145 1.75 ;
      RECT  9.56 1.21 9.68 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  5.87 0.05 6.0 0.345 ;
      RECT  6.39 0.05 6.52 0.345 ;
      RECT  6.91 0.05 7.04 0.345 ;
      RECT  7.455 0.05 7.585 0.345 ;
      RECT  7.975 0.05 8.105 0.345 ;
      RECT  8.495 0.05 8.625 0.345 ;
      RECT  9.015 0.05 9.145 0.345 ;
      RECT  3.29 0.05 3.4 0.36 ;
      RECT  3.79 0.05 3.92 0.36 ;
      RECT  4.31 0.05 4.44 0.36 ;
      RECT  4.83 0.05 4.96 0.36 ;
      RECT  0.585 0.05 0.705 0.585 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.355 0.05 5.475 0.59 ;
      RECT  9.56 0.05 9.68 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.615 0.435 9.45 0.565 ;
      RECT  5.615 0.565 8.05 0.605 ;
      RECT  7.73 0.605 8.05 1.11 ;
      RECT  5.62 1.11 9.45 1.29 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.615 0.14 3.2 0.23 ;
      RECT  1.615 0.23 1.735 0.32 ;
      RECT  3.11 0.23 3.2 0.45 ;
      RECT  1.04 0.32 1.735 0.44 ;
      RECT  3.11 0.45 4.225 0.54 ;
      RECT  3.11 0.54 3.2 0.84 ;
      RECT  3.535 0.54 3.64 1.045 ;
      RECT  2.74 0.84 3.2 0.93 ;
      RECT  2.74 0.93 2.83 1.36 ;
      RECT  3.535 1.045 4.225 1.155 ;
      RECT  2.085 1.36 2.83 1.48 ;
      RECT  1.85 0.32 3.02 0.41 ;
      RECT  1.85 0.41 1.94 0.53 ;
      RECT  2.915 0.41 3.02 0.54 ;
      RECT  0.795 0.53 1.94 0.62 ;
      RECT  1.44 0.62 1.54 1.145 ;
      RECT  1.225 1.145 1.54 1.16 ;
      RECT  0.795 1.16 1.54 1.25 ;
      RECT  4.575 0.455 5.265 0.575 ;
      RECT  4.575 0.575 4.695 1.255 ;
      RECT  3.11 1.255 5.265 1.345 ;
      RECT  3.11 1.345 3.2 1.57 ;
      RECT  2.03 0.5 2.825 0.59 ;
      RECT  2.03 0.59 2.12 0.885 ;
      RECT  1.63 0.885 2.12 0.975 ;
      RECT  1.63 0.975 1.72 1.44 ;
      RECT  1.045 1.44 1.72 1.56 ;
      RECT  1.63 1.56 1.72 1.57 ;
      RECT  1.63 1.57 3.2 1.66 ;
      RECT  5.43 0.775 7.605 0.895 ;
      RECT  5.43 0.895 5.53 1.31 ;
      RECT  1.035 0.755 1.325 0.93 ;
      RECT  1.035 0.93 1.125 0.98 ;
      RECT  0.325 0.29 0.43 0.98 ;
      RECT  0.325 0.98 1.125 1.07 ;
      RECT  0.325 1.07 0.43 1.45 ;
      RECT  1.825 1.115 2.54 1.205 ;
      RECT  2.36 1.205 2.54 1.25 ;
      RECT  2.92 1.03 3.02 1.47 ;
      LAYER M2 ;
      RECT  1.36 1.15 5.57 1.25 ;
      LAYER V1 ;
      RECT  1.4 1.15 1.5 1.25 ;
      RECT  2.4 1.15 2.5 1.25 ;
      RECT  2.92 1.15 3.02 1.25 ;
      RECT  5.43 1.15 5.53 1.25 ;
  END
END SEN_MUX2_DG_16
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_DG_2
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_DG_2
  CLASS CORE ;
  FOREIGN SEN_MUX2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.71 0.65 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.32 0.77 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.14 1.215 0.235 ;
      RECT  0.75 0.235 0.85 0.49 ;
      RECT  0.325 0.49 0.85 0.58 ;
      RECT  0.325 0.58 0.45 0.745 ;
      RECT  0.225 0.745 0.45 0.915 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.405 1.4 0.535 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.47 1.38 1.6 1.75 ;
      RECT  2.005 1.21 2.125 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.395 0.05 0.525 0.4 ;
      RECT  1.47 0.05 1.6 0.48 ;
      RECT  2.005 0.05 2.125 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.745 0.31 1.915 0.49 ;
      RECT  1.825 0.49 1.915 1.015 ;
      RECT  1.75 1.015 1.915 1.1 ;
      RECT  1.75 1.1 1.855 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.045 0.33 0.235 0.5 ;
      RECT  0.045 0.5 0.135 1.22 ;
      RECT  0.045 1.22 0.86 1.31 ;
      RECT  0.77 0.67 0.86 1.22 ;
      RECT  0.77 1.31 0.86 1.51 ;
      RECT  0.77 1.51 1.22 1.62 ;
      RECT  0.95 0.375 1.04 0.59 ;
      RECT  0.95 0.59 1.735 0.68 ;
      RECT  1.645 0.68 1.735 0.925 ;
      RECT  0.95 0.68 1.04 1.39 ;
  END
END SEN_MUX2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_DG_4
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_DG_4
  CLASS CORE ;
  FOREIGN SEN_MUX2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.65 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.05 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.605 2.28 0.935 ;
      RECT  1.15 0.51 1.25 0.735 ;
      RECT  1.15 0.735 1.33 0.925 ;
      LAYER M2 ;
      RECT  1.11 0.75 2.29 0.85 ;
      LAYER V1 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.105 1.21 1.225 1.75 ;
      RECT  2.73 1.44 2.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  2.73 0.05 2.86 0.375 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.51 1.015 0.615 ;
      RECT  0.34 0.615 0.45 1.11 ;
      RECT  0.34 1.11 0.85 1.18 ;
      RECT  0.34 1.18 1.015 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.17 0.19 2.325 0.4 ;
      RECT  2.17 0.4 2.28 0.49 ;
      RECT  2.98 0.225 3.115 0.465 ;
      RECT  2.75 0.465 3.115 0.555 ;
      RECT  2.75 0.555 2.84 1.26 ;
      RECT  2.49 1.26 3.115 1.35 ;
      RECT  2.49 1.35 2.58 1.465 ;
      RECT  2.995 1.35 3.115 1.535 ;
      RECT  1.635 1.465 2.58 1.585 ;
      RECT  2.37 0.49 2.645 0.58 ;
      RECT  2.37 0.58 2.46 1.03 ;
      RECT  2.29 1.03 2.46 1.14 ;
      RECT  2.29 1.14 2.4 1.275 ;
      RECT  1.655 0.235 1.87 0.405 ;
      RECT  1.78 0.405 1.87 1.275 ;
      RECT  1.78 1.275 2.4 1.365 ;
      RECT  1.42 0.21 1.525 0.755 ;
      RECT  1.42 0.755 1.69 0.925 ;
      RECT  1.42 0.925 1.525 1.56 ;
      RECT  0.55 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
      RECT  1.96 0.445 2.06 1.185 ;
      LAYER M2 ;
      RECT  2.14 0.35 3.12 0.45 ;
      RECT  0.91 0.95 2.1 1.05 ;
      LAYER V1 ;
      RECT  2.18 0.35 2.28 0.45 ;
      RECT  2.98 0.35 3.08 0.45 ;
      RECT  0.95 0.95 1.05 1.05 ;
      RECT  1.96 0.95 2.06 1.05 ;
  END
END SEN_MUX2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_DG_8
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_DG_8
  CLASS CORE ;
  FOREIGN SEN_MUX2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.51 4.65 0.71 ;
      RECT  4.15 0.71 4.65 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.685 5.05 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 3.85 0.785 ;
      RECT  3.39 0.785 3.85 0.895 ;
      RECT  2.23 0.58 2.33 1.0 ;
      LAYER M2 ;
      RECT  2.19 0.75 3.89 0.85 ;
      LAYER V1 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.23 0.75 2.33 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.455 1.75 1.75 ;
      RECT  2.145 1.43 2.27 1.75 ;
      RECT  3.975 1.41 4.1 1.75 ;
      RECT  4.49 1.41 4.62 1.75 ;
      RECT  5.015 1.215 5.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  3.975 0.05 4.1 0.36 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  1.62 0.05 1.75 0.39 ;
      RECT  2.14 0.05 2.27 0.39 ;
      RECT  4.49 0.05 4.62 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.015 0.05 5.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.325 0.51 2.05 0.69 ;
      RECT  0.75 0.69 0.92 1.11 ;
      RECT  0.325 1.11 1.75 1.27 ;
      RECT  0.325 1.27 2.05 1.29 ;
      RECT  1.66 1.29 2.05 1.36 ;
      RECT  1.885 1.36 2.05 1.49 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.645 0.2 3.88 0.305 ;
      RECT  2.645 0.305 2.735 0.57 ;
      RECT  2.645 0.57 2.855 0.66 ;
      RECT  2.765 0.66 2.855 1.25 ;
      RECT  1.01 0.79 2.095 0.89 ;
      RECT  2.005 0.89 2.095 1.09 ;
      RECT  2.005 1.09 2.33 1.18 ;
      RECT  2.24 1.18 2.33 1.25 ;
      RECT  2.24 1.25 2.855 1.34 ;
      RECT  2.76 1.34 2.855 1.44 ;
      RECT  2.76 1.44 3.88 1.56 ;
      RECT  2.885 0.395 3.885 0.475 ;
      RECT  2.885 0.475 4.405 0.485 ;
      RECT  3.795 0.485 4.405 0.58 ;
      RECT  3.96 0.58 4.405 0.595 ;
      RECT  3.96 0.595 4.05 1.0 ;
      RECT  3.4 1.0 4.405 1.12 ;
      RECT  2.945 0.575 3.62 0.665 ;
      RECT  2.945 0.665 3.035 1.21 ;
      RECT  2.945 1.21 4.86 1.3 ;
      RECT  4.755 0.39 4.86 1.21 ;
      RECT  2.42 0.45 2.51 0.75 ;
      RECT  2.42 0.75 2.675 0.925 ;
      RECT  2.42 0.925 2.52 1.16 ;
  END
END SEN_MUX2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_S_0P5
#      Description : "2-1 multiplexer, symmetric rise/fall"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_S_0P5
  CLASS CORE ;
  FOREIGN SEN_MUX2_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.705 1.66 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0396 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.41 1.495 0.58 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.715 1.39 1.845 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.42 0.05 0.55 0.39 ;
      RECT  1.74 0.05 1.86 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.265 2.12 0.435 ;
      RECT  1.95 0.435 2.05 1.39 ;
      RECT  1.95 1.39 2.12 1.56 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.11 0.14 1.65 0.23 ;
      RECT  1.56 0.23 1.65 0.505 ;
      RECT  1.11 0.23 1.215 1.46 ;
      RECT  1.56 0.505 1.85 0.595 ;
      RECT  1.75 0.595 1.85 0.88 ;
      RECT  1.355 0.32 1.47 0.535 ;
      RECT  1.355 0.535 1.46 1.46 ;
      RECT  0.74 0.18 0.84 1.225 ;
      RECT  0.14 0.18 0.26 1.315 ;
      RECT  0.14 1.315 1.02 1.405 ;
      RECT  0.93 0.515 1.02 1.315 ;
      RECT  0.93 1.405 1.02 1.55 ;
      RECT  0.93 1.55 1.38 1.66 ;
  END
END SEN_MUX2_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_S_1
#      Description : "2-1 multiplexer, symmetric rise/fall"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_S_1
  CLASS CORE ;
  FOREIGN SEN_MUX2_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0393 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.705 1.66 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0393 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.425 1.435 0.555 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.675 1.41 1.805 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  1.74 0.05 1.865 0.385 ;
      RECT  0.42 0.05 0.55 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.12 0.69 ;
      RECT  1.95 0.69 2.05 1.11 ;
      RECT  1.95 1.11 2.12 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.11 0.14 1.65 0.23 ;
      RECT  1.56 0.23 1.65 0.495 ;
      RECT  1.11 0.23 1.215 1.385 ;
      RECT  1.56 0.495 1.85 0.585 ;
      RECT  1.75 0.585 1.85 0.93 ;
      RECT  1.355 0.32 1.47 0.535 ;
      RECT  1.355 0.535 1.46 1.41 ;
      RECT  0.74 0.225 0.84 1.16 ;
      RECT  0.14 0.18 0.26 1.25 ;
      RECT  0.14 1.25 1.02 1.34 ;
      RECT  0.93 0.51 1.02 1.25 ;
      RECT  0.14 1.34 0.26 1.5 ;
      RECT  0.93 1.34 1.02 1.55 ;
      RECT  0.93 1.55 1.375 1.66 ;
  END
END SEN_MUX2_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_S_2
#      Description : "2-1 multiplexer, symmetric rise/fall"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_S_2
  CLASS CORE ;
  FOREIGN SEN_MUX2_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.47 0.75 0.56 0.9 ;
      RECT  0.47 0.9 0.85 1.015 ;
      RECT  0.35 1.015 0.85 1.105 ;
      RECT  0.35 1.105 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 1.01 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.235 0.5 0.74 0.59 ;
      RECT  0.65 0.59 0.74 0.7 ;
      RECT  0.235 0.59 0.335 0.925 ;
      RECT  0.65 0.7 1.25 0.79 ;
      RECT  1.15 0.79 1.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1278 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.59 0.47 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.86 1.57 0.985 1.75 ;
      RECT  2.37 1.515 2.5 1.75 ;
      RECT  2.88 1.46 3.05 1.75 ;
      RECT  3.425 1.41 3.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.845 0.05 1.015 0.19 ;
      RECT  2.39 0.05 2.5 0.225 ;
      RECT  0.31 0.05 0.44 0.39 ;
      RECT  3.425 0.05 3.545 0.39 ;
      RECT  2.905 0.05 3.025 0.605 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.31 3.275 0.505 ;
      RECT  3.15 0.505 3.45 0.595 ;
      RECT  3.35 0.595 3.45 1.0 ;
      RECT  3.15 1.0 3.45 1.09 ;
      RECT  3.15 1.09 3.27 1.505 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.25 0.14 2.3 0.23 ;
      RECT  2.21 0.23 2.3 0.315 ;
      RECT  2.21 0.315 2.76 0.405 ;
      RECT  2.65 0.405 2.76 1.1 ;
      RECT  2.495 1.1 2.76 1.135 ;
      RECT  1.93 1.135 2.76 1.19 ;
      RECT  1.93 1.19 2.585 1.225 ;
      RECT  1.93 1.225 2.02 1.39 ;
      RECT  0.55 0.3 0.92 0.41 ;
      RECT  0.83 0.41 0.92 0.515 ;
      RECT  0.83 0.515 1.94 0.605 ;
      RECT  1.85 0.605 1.94 0.685 ;
      RECT  1.385 0.605 1.48 1.21 ;
      RECT  0.56 1.21 1.48 1.3 ;
      RECT  1.57 0.775 1.935 0.865 ;
      RECT  1.57 0.865 1.66 1.39 ;
      RECT  0.055 0.19 0.19 0.41 ;
      RECT  0.055 0.41 0.145 1.39 ;
      RECT  0.055 1.39 1.66 1.48 ;
      RECT  0.055 1.48 0.175 1.59 ;
      RECT  2.87 0.795 3.25 0.885 ;
      RECT  2.87 0.885 2.96 1.28 ;
      RECT  2.715 1.28 2.96 1.315 ;
      RECT  2.15 1.315 2.96 1.37 ;
      RECT  2.15 1.37 2.805 1.405 ;
      RECT  2.15 1.405 2.24 1.57 ;
      RECT  1.01 0.335 2.12 0.425 ;
      RECT  2.03 0.425 2.12 0.52 ;
      RECT  2.03 0.52 2.21 0.69 ;
      RECT  2.03 0.69 2.12 0.955 ;
      RECT  1.75 0.955 2.12 1.045 ;
      RECT  1.75 1.045 1.84 1.57 ;
      RECT  1.08 1.57 2.24 1.66 ;
  END
END SEN_MUX2_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_S_4
#      Description : "2-1 multiplexer, symmetric rise/fall"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_S_4
  CLASS CORE ;
  FOREIGN SEN_MUX2_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.7 1.05 0.89 ;
      RECT  0.55 0.89 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.65 0.89 ;
      RECT  4.15 0.89 4.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.5 1.25 0.59 ;
      RECT  0.35 0.59 0.45 0.72 ;
      RECT  1.15 0.59 1.25 0.8 ;
      RECT  0.255 0.72 0.45 0.96 ;
      RECT  1.15 0.8 2.2 0.89 ;
      RECT  1.15 0.89 1.25 0.985 ;
      RECT  0.35 0.96 0.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2247 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.29 1.6 0.5 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.83 1.6 1.04 1.75 ;
      RECT  1.37 1.6 1.58 1.75 ;
      RECT  3.71 1.6 3.92 1.75 ;
      RECT  4.315 1.6 4.525 1.75 ;
      RECT  4.855 1.6 5.065 1.75 ;
      RECT  5.465 1.43 5.615 1.75 ;
      RECT  6.005 1.21 6.125 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  3.83 0.05 4.03 0.185 ;
      RECT  0.81 0.05 1.02 0.2 ;
      RECT  1.35 0.05 1.56 0.2 ;
      RECT  5.475 0.05 5.6 0.375 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  4.435 0.05 4.565 0.4 ;
      RECT  4.955 0.05 5.095 0.59 ;
      RECT  6.005 0.05 6.125 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.195 0.51 5.855 0.69 ;
      RECT  5.75 0.69 5.855 1.11 ;
      RECT  5.22 1.11 5.855 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.405 0.16 3.74 0.205 ;
      RECT  1.79 0.205 3.74 0.25 ;
      RECT  3.65 0.25 3.74 0.275 ;
      RECT  1.79 0.25 2.515 0.305 ;
      RECT  3.65 0.275 4.3 0.365 ;
      RECT  4.18 0.365 4.3 0.49 ;
      RECT  4.18 0.49 4.85 0.59 ;
      RECT  4.75 0.59 4.85 1.22 ;
      RECT  2.905 1.22 4.85 1.31 ;
      RECT  0.54 0.29 1.45 0.39 ;
      RECT  1.35 0.39 1.45 0.6 ;
      RECT  1.35 0.6 3.055 0.69 ;
      RECT  2.845 0.545 3.055 0.6 ;
      RECT  2.32 0.69 2.42 1.015 ;
      RECT  1.36 1.015 2.42 1.105 ;
      RECT  1.36 1.105 1.46 1.205 ;
      RECT  0.56 1.205 1.46 1.32 ;
      RECT  3.38 0.4 3.565 0.65 ;
      RECT  2.52 0.8 3.07 0.89 ;
      RECT  2.52 0.89 2.62 1.2 ;
      RECT  1.56 1.2 2.62 1.29 ;
      RECT  1.56 1.29 1.655 1.41 ;
      RECT  0.055 0.22 0.185 0.44 ;
      RECT  0.055 0.44 0.155 1.41 ;
      RECT  0.055 1.41 1.655 1.5 ;
      RECT  0.055 1.5 0.2 1.6 ;
      RECT  4.95 0.8 5.64 0.9 ;
      RECT  4.95 0.9 5.05 1.41 ;
      RECT  2.59 0.36 3.275 0.4 ;
      RECT  1.54 0.4 3.275 0.45 ;
      RECT  1.54 0.45 2.77 0.49 ;
      RECT  3.16 0.45 3.275 0.97 ;
      RECT  3.16 0.97 3.795 1.0 ;
      RECT  3.685 0.455 3.795 0.97 ;
      RECT  2.71 1.0 3.795 1.09 ;
      RECT  2.71 1.09 2.81 1.41 ;
      RECT  1.87 1.41 5.05 1.51 ;
      LAYER M2 ;
      RECT  2.8 0.55 3.65 0.65 ;
      LAYER V1 ;
      RECT  2.885 0.55 2.985 0.65 ;
      RECT  3.42 0.55 3.52 0.65 ;
  END
END SEN_MUX2_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_S_8
#      Description : "2-1 multiplexer, symmetric rise/fall"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_S_8
  CLASS CORE ;
  FOREIGN SEN_MUX2_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.65 0.795 1.63 0.885 ;
      RECT  0.65 0.885 0.95 1.09 ;
      LAYER M2 ;
      RECT  0.5 0.95 1.1 1.05 ;
      LAYER V1 ;
      RECT  0.65 0.95 0.75 1.05 ;
      RECT  0.85 0.95 0.95 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4536 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.71 6.83 0.9 ;
      LAYER M2 ;
      RECT  6.1 0.75 6.7 0.85 ;
      LAYER V1 ;
      RECT  6.25 0.75 6.35 0.85 ;
      RECT  6.45 0.75 6.55 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4536 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.5 0.45 0.615 ;
      RECT  0.35 0.615 1.85 0.705 ;
      RECT  0.35 0.705 0.45 0.755 ;
      RECT  1.75 0.705 1.85 0.81 ;
      RECT  0.255 0.755 0.45 0.925 ;
      RECT  1.75 0.81 3.23 0.91 ;
      RECT  0.35 0.925 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4017 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.42 0.45 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  0.86 1.63 1.07 1.75 ;
      RECT  1.535 1.455 1.66 1.75 ;
      RECT  2.02 1.48 2.19 1.75 ;
      RECT  5.95 1.495 6.12 1.75 ;
      RECT  6.47 1.495 6.64 1.75 ;
      RECT  6.98 1.495 7.17 1.75 ;
      RECT  7.535 1.235 7.655 1.75 ;
      RECT  8.05 1.425 8.18 1.75 ;
      RECT  8.57 1.43 8.7 1.75 ;
      RECT  9.09 1.43 9.22 1.75 ;
      RECT  9.615 1.21 9.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  8.03 0.05 8.2 0.305 ;
      RECT  8.54 0.05 8.73 0.305 ;
      RECT  9.07 0.05 9.24 0.305 ;
      RECT  0.81 0.05 1.0 0.31 ;
      RECT  1.33 0.05 1.52 0.31 ;
      RECT  1.85 0.05 2.05 0.31 ;
      RECT  6.99 0.05 7.16 0.32 ;
      RECT  6.47 0.05 6.64 0.33 ;
      RECT  5.975 0.05 6.1 0.345 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  7.51 0.05 7.68 0.52 ;
      RECT  9.615 0.05 9.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.795 0.295 7.915 0.4 ;
      RECT  7.795 0.4 9.52 0.52 ;
      RECT  8.35 0.31 8.45 0.4 ;
      RECT  9.35 0.31 9.52 0.4 ;
      RECT  9.35 0.52 9.52 1.11 ;
      RECT  8.805 1.11 9.52 1.2 ;
      RECT  7.77 1.2 9.52 1.29 ;
      RECT  7.77 1.29 8.98 1.33 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.585 0.145 5.875 0.26 ;
      RECT  2.585 0.26 3.815 0.31 ;
      RECT  5.715 0.26 5.875 0.435 ;
      RECT  5.715 0.435 7.405 0.61 ;
      RECT  7.125 0.61 8.675 0.71 ;
      RECT  8.485 0.71 8.675 1.0 ;
      RECT  7.195 1.0 8.675 1.11 ;
      RECT  7.195 1.11 7.425 1.22 ;
      RECT  5.7 1.22 7.425 1.38 ;
      RECT  5.7 1.38 5.85 1.46 ;
      RECT  4.63 1.46 5.85 1.53 ;
      RECT  4.12 1.53 5.85 1.645 ;
      RECT  0.56 0.4 2.275 0.525 ;
      RECT  2.125 0.525 2.275 0.6 ;
      RECT  2.125 0.6 5.375 0.69 ;
      RECT  4.11 0.55 5.375 0.6 ;
      RECT  5.255 0.69 5.375 1.0 ;
      RECT  3.865 1.0 5.375 1.11 ;
      RECT  3.865 1.11 3.995 1.115 ;
      RECT  3.62 1.115 3.995 1.21 ;
      RECT  1.32 1.21 3.995 1.26 ;
      RECT  1.32 1.26 3.74 1.35 ;
      RECT  1.32 1.35 1.445 1.42 ;
      RECT  0.58 1.42 1.445 1.51 ;
      RECT  0.58 1.51 0.705 1.63 ;
      RECT  3.34 0.8 5.145 0.91 ;
      RECT  3.34 0.91 3.46 1.0 ;
      RECT  1.14 1.0 3.46 1.12 ;
      RECT  1.14 1.12 1.23 1.21 ;
      RECT  0.065 0.29 0.2 0.51 ;
      RECT  0.065 0.51 0.155 1.21 ;
      RECT  0.065 1.21 1.23 1.33 ;
      RECT  0.065 1.33 0.185 1.62 ;
      RECT  6.94 0.8 8.375 0.91 ;
      RECT  6.94 0.91 7.06 1.01 ;
      RECT  2.365 0.17 2.495 0.42 ;
      RECT  2.365 0.42 5.62 0.45 ;
      RECT  3.9 0.35 5.62 0.42 ;
      RECT  2.365 0.45 4.0 0.51 ;
      RECT  5.465 0.45 5.62 1.01 ;
      RECT  5.465 1.01 7.06 1.13 ;
      RECT  5.465 1.13 5.6 1.2 ;
      RECT  4.085 1.2 5.6 1.35 ;
      RECT  3.885 1.35 5.6 1.365 ;
      RECT  3.885 1.365 4.435 1.44 ;
      RECT  3.885 1.44 4.03 1.45 ;
      RECT  2.51 1.45 4.03 1.61 ;
  END
END SEN_MUX2_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_G_1
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_G_1
  CLASS CORE ;
  FOREIGN SEN_MUX2_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.71 0.65 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.845 1.3 1.025 ;
      RECT  1.15 1.025 1.25 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.165 1.14 0.255 ;
      RECT  0.55 0.255 0.65 0.5 ;
      RECT  0.35 0.5 0.65 0.59 ;
      RECT  0.35 0.59 0.45 0.745 ;
      RECT  0.26 0.745 0.45 0.925 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.46 0.46 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.35 1.39 1.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.345 0.05 1.475 0.36 ;
      RECT  0.33 0.05 0.455 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.61 0.34 1.73 1.11 ;
      RECT  1.55 1.11 1.73 1.2 ;
      RECT  1.55 1.2 1.65 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.81 0.45 1.52 0.54 ;
      RECT  1.43 0.54 1.52 0.925 ;
      RECT  0.96 0.54 1.05 1.495 ;
      RECT  0.8 1.495 1.05 1.585 ;
      RECT  0.065 0.36 0.17 1.28 ;
      RECT  0.065 1.28 0.865 1.37 ;
      RECT  0.77 0.785 0.865 1.28 ;
  END
END SEN_MUX2_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_G_12
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_G_12
  CLASS CORE ;
  FOREIGN SEN_MUX2_G_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.51 6.25 0.71 ;
      RECT  5.125 0.71 6.25 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.73 0.71 7.45 0.89 ;
      RECT  7.35 0.89 7.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.07 0.75 3.25 0.785 ;
      RECT  3.07 0.785 3.77 0.89 ;
      RECT  0.35 0.71 1.105 0.89 ;
      LAYER M2 ;
      RECT  0.96 0.75 3.25 0.85 ;
      LAYER V1 ;
      RECT  3.11 0.75 3.21 0.85 ;
      RECT  1.005 0.75 1.105 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5832 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 11.0 1.85 ;
      RECT  0.845 1.21 0.965 1.75 ;
      RECT  4.59 1.45 4.7 1.75 ;
      RECT  5.09 1.45 5.22 1.75 ;
      RECT  5.61 1.45 5.74 1.75 ;
      RECT  6.13 1.45 6.26 1.75 ;
      RECT  6.65 1.45 6.78 1.75 ;
      RECT  7.17 1.45 7.3 1.75 ;
      RECT  7.69 1.41 7.82 1.75 ;
      RECT  8.21 1.415 8.34 1.75 ;
      RECT  8.73 1.41 8.86 1.75 ;
      RECT  9.25 1.41 9.38 1.75 ;
      RECT  9.77 1.41 9.9 1.75 ;
      RECT  10.29 1.41 10.42 1.75 ;
      RECT  10.815 1.21 10.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      RECT  8.21 0.05 8.34 0.35 ;
      RECT  8.73 0.05 8.86 0.35 ;
      RECT  9.25 0.05 9.38 0.35 ;
      RECT  9.77 0.05 9.9 0.35 ;
      RECT  10.29 0.05 10.42 0.35 ;
      RECT  4.59 0.05 4.7 0.385 ;
      RECT  5.09 0.05 5.22 0.385 ;
      RECT  5.61 0.05 5.74 0.385 ;
      RECT  6.13 0.05 6.26 0.385 ;
      RECT  6.65 0.05 6.78 0.385 ;
      RECT  7.17 0.05 7.3 0.385 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.845 0.05 0.965 0.59 ;
      RECT  7.695 0.05 7.815 0.59 ;
      RECT  10.815 0.05 10.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.955 0.44 10.725 0.56 ;
      RECT  7.955 0.56 9.86 0.61 ;
      RECT  9.62 0.61 9.86 1.11 ;
      RECT  7.95 1.11 10.675 1.29 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.39 0.18 4.5 0.255 ;
      RECT  1.305 0.255 4.5 0.27 ;
      RECT  1.305 0.27 2.52 0.375 ;
      RECT  4.41 0.27 4.5 0.475 ;
      RECT  4.41 0.475 6.045 0.595 ;
      RECT  4.41 0.595 4.945 0.605 ;
      RECT  4.81 0.605 4.945 0.8 ;
      RECT  3.97 0.8 4.945 0.93 ;
      RECT  4.81 0.93 4.945 1.03 ;
      RECT  3.97 0.93 4.1 1.34 ;
      RECT  4.81 1.03 6.045 1.15 ;
      RECT  2.865 1.34 4.1 1.46 ;
      RECT  2.63 0.365 4.32 0.47 ;
      RECT  2.63 0.47 2.76 0.52 ;
      RECT  4.215 0.47 4.32 0.59 ;
      RECT  1.055 0.52 2.76 0.62 ;
      RECT  2.19 0.62 2.76 0.65 ;
      RECT  2.19 0.65 2.32 1.145 ;
      RECT  2.005 1.145 2.32 1.16 ;
      RECT  1.055 1.16 2.32 1.265 ;
      RECT  6.39 0.48 7.605 0.6 ;
      RECT  6.39 0.6 6.52 1.24 ;
      RECT  4.38 1.24 7.58 1.36 ;
      RECT  4.38 1.36 4.5 1.55 ;
      RECT  2.85 0.56 4.125 0.66 ;
      RECT  2.85 0.66 2.98 0.845 ;
      RECT  2.41 0.845 2.98 0.975 ;
      RECT  2.41 0.975 2.525 1.44 ;
      RECT  1.305 1.44 2.525 1.55 ;
      RECT  1.305 1.55 4.5 1.56 ;
      RECT  2.41 1.56 4.5 1.66 ;
      RECT  1.285 0.79 2.1 0.895 ;
      RECT  1.285 0.895 1.375 0.98 ;
      RECT  0.64 0.98 1.375 1.07 ;
      RECT  0.64 1.07 0.73 1.16 ;
      RECT  0.065 0.48 0.755 0.6 ;
      RECT  0.065 0.6 0.185 1.16 ;
      RECT  0.065 1.16 0.73 1.28 ;
      RECT  7.67 0.76 9.495 0.895 ;
      RECT  7.67 0.895 7.77 1.29 ;
      RECT  4.19 1.02 4.44 1.135 ;
      RECT  4.19 1.135 4.29 1.45 ;
      RECT  2.63 1.115 3.84 1.205 ;
      RECT  3.14 1.205 3.32 1.25 ;
      LAYER M2 ;
      RECT  2.14 1.15 7.81 1.25 ;
      LAYER V1 ;
      RECT  2.18 1.15 2.28 1.25 ;
      RECT  3.18 1.15 3.28 1.25 ;
      RECT  4.19 1.15 4.29 1.25 ;
      RECT  7.67 1.15 7.77 1.25 ;
  END
END SEN_MUX2_G_12
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_G_16
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_G_16
  CLASS CORE ;
  FOREIGN SEN_MUX2_G_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.51 8.05 0.71 ;
      RECT  6.75 0.71 8.05 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.75 0.71 9.65 0.89 ;
      RECT  9.55 0.89 9.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.85 0.75 4.03 0.785 ;
      RECT  3.85 0.785 4.98 0.89 ;
      RECT  0.55 0.71 1.2 0.89 ;
      LAYER M2 ;
      RECT  1.06 0.75 4.03 0.85 ;
      LAYER V1 ;
      RECT  3.89 0.75 3.99 0.85 ;
      RECT  1.1 0.75 1.2 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 14.4 1.85 ;
      RECT  0.58 1.435 0.71 1.75 ;
      RECT  1.105 1.21 1.215 1.75 ;
      RECT  5.89 1.455 6.0 1.75 ;
      RECT  6.39 1.455 6.52 1.75 ;
      RECT  6.91 1.455 7.04 1.75 ;
      RECT  7.43 1.455 7.56 1.75 ;
      RECT  7.95 1.455 8.08 1.75 ;
      RECT  8.47 1.455 8.6 1.75 ;
      RECT  8.99 1.455 9.12 1.75 ;
      RECT  9.51 1.455 9.64 1.75 ;
      RECT  10.03 1.41 10.16 1.75 ;
      RECT  10.55 1.41 10.68 1.75 ;
      RECT  11.07 1.41 11.2 1.75 ;
      RECT  11.59 1.41 11.72 1.75 ;
      RECT  12.11 1.41 12.24 1.75 ;
      RECT  12.63 1.41 12.76 1.75 ;
      RECT  13.15 1.41 13.28 1.75 ;
      RECT  13.67 1.41 13.8 1.75 ;
      RECT  14.205 1.21 14.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 14.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 14.4 0.05 ;
      RECT  5.89 0.05 6.0 0.345 ;
      RECT  6.39 0.05 6.52 0.345 ;
      RECT  6.91 0.05 7.04 0.345 ;
      RECT  7.43 0.05 7.56 0.345 ;
      RECT  8.47 0.05 8.6 0.345 ;
      RECT  8.99 0.05 9.12 0.345 ;
      RECT  9.51 0.05 9.64 0.345 ;
      RECT  10.55 0.05 10.68 0.35 ;
      RECT  11.07 0.05 11.2 0.35 ;
      RECT  11.59 0.05 11.72 0.35 ;
      RECT  12.11 0.05 12.24 0.35 ;
      RECT  12.63 0.05 12.76 0.35 ;
      RECT  13.15 0.05 13.28 0.35 ;
      RECT  13.67 0.05 13.8 0.35 ;
      RECT  0.58 0.05 0.71 0.365 ;
      RECT  7.95 0.05 8.08 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.105 0.05 1.215 0.59 ;
      RECT  10.035 0.05 10.155 0.59 ;
      RECT  14.205 0.05 14.325 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 14.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.295 0.44 14.08 0.56 ;
      RECT  10.295 0.56 12.86 0.64 ;
      RECT  12.54 0.64 12.86 1.09 ;
      RECT  10.29 1.09 12.86 1.11 ;
      RECT  10.29 1.11 14.055 1.29 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.17 0.18 5.8 0.25 ;
      RECT  1.565 0.25 5.8 0.27 ;
      RECT  1.565 0.27 3.3 0.375 ;
      RECT  5.71 0.27 5.8 0.435 ;
      RECT  2.415 0.375 2.8 0.45 ;
      RECT  5.71 0.435 7.815 0.565 ;
      RECT  6.15 0.31 6.25 0.435 ;
      RECT  6.67 0.31 6.77 0.435 ;
      RECT  7.695 0.345 7.815 0.435 ;
      RECT  6.285 0.565 6.455 1.005 ;
      RECT  5.27 0.8 6.01 0.93 ;
      RECT  5.89 0.93 6.01 1.005 ;
      RECT  5.27 0.93 5.4 1.34 ;
      RECT  5.89 1.005 7.865 1.135 ;
      RECT  3.645 1.34 5.4 1.46 ;
      RECT  3.405 0.365 5.62 0.47 ;
      RECT  3.405 0.47 3.54 0.555 ;
      RECT  5.515 0.47 5.62 0.59 ;
      RECT  1.305 0.555 3.54 0.655 ;
      RECT  2.93 0.655 3.54 0.685 ;
      RECT  2.93 0.685 3.1 1.145 ;
      RECT  2.375 1.145 3.1 1.16 ;
      RECT  1.305 1.16 3.1 1.25 ;
      RECT  8.165 0.435 9.945 0.565 ;
      RECT  8.42 0.565 8.59 1.225 ;
      RECT  5.68 1.225 8.59 1.235 ;
      RECT  5.68 1.235 9.92 1.365 ;
      RECT  6.15 1.365 6.25 1.49 ;
      RECT  6.69 1.365 6.79 1.49 ;
      RECT  7.18 1.365 7.28 1.49 ;
      RECT  7.67 1.365 7.77 1.49 ;
      RECT  8.235 1.365 8.335 1.49 ;
      RECT  8.725 1.365 8.825 1.49 ;
      RECT  5.68 1.365 5.8 1.55 ;
      RECT  3.63 0.56 5.425 0.66 ;
      RECT  3.63 0.66 3.74 0.845 ;
      RECT  3.19 0.845 3.74 0.955 ;
      RECT  3.19 0.955 3.3 1.44 ;
      RECT  2.685 1.35 2.865 1.44 ;
      RECT  1.565 1.44 3.3 1.55 ;
      RECT  1.565 1.55 5.8 1.56 ;
      RECT  3.19 1.56 5.8 1.66 ;
      RECT  1.735 0.785 2.84 0.89 ;
      RECT  1.735 0.89 1.825 0.98 ;
      RECT  0.9 0.98 1.825 1.07 ;
      RECT  0.9 1.07 0.99 1.225 ;
      RECT  0.325 0.455 1.015 0.575 ;
      RECT  0.325 0.575 0.445 1.225 ;
      RECT  0.325 1.225 0.99 1.345 ;
      RECT  10.01 0.775 12.4 0.895 ;
      RECT  10.01 0.895 10.11 1.31 ;
      RECT  5.49 1.02 5.74 1.135 ;
      RECT  5.49 1.135 5.59 1.45 ;
      RECT  3.435 1.1 5.165 1.22 ;
      RECT  3.92 1.22 4.1 1.25 ;
      RECT  3.435 1.22 3.555 1.31 ;
      LAYER M2 ;
      RECT  2.415 0.35 6.81 0.45 ;
      RECT  2.92 1.15 10.15 1.25 ;
      RECT  2.685 1.35 8.865 1.45 ;
      LAYER V1 ;
      RECT  2.46 0.35 2.56 0.45 ;
      RECT  2.66 0.35 2.76 0.45 ;
      RECT  6.15 0.35 6.25 0.45 ;
      RECT  6.67 0.35 6.77 0.45 ;
      RECT  2.96 1.15 3.06 1.25 ;
      RECT  3.96 1.15 4.06 1.25 ;
      RECT  5.49 1.15 5.59 1.25 ;
      RECT  10.01 1.15 10.11 1.25 ;
      RECT  2.725 1.35 2.825 1.45 ;
      RECT  3.2 1.35 3.3 1.45 ;
      RECT  6.15 1.35 6.25 1.45 ;
      RECT  6.69 1.35 6.79 1.45 ;
      RECT  7.18 1.35 7.28 1.45 ;
      RECT  7.67 1.35 7.77 1.45 ;
      RECT  8.235 1.35 8.335 1.45 ;
      RECT  8.725 1.35 8.825 1.45 ;
  END
END SEN_MUX2_G_16
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_G_2
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_G_2
  CLASS CORE ;
  FOREIGN SEN_MUX2_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.6 ;
      RECT  0.55 0.6 0.85 0.69 ;
      RECT  0.55 0.69 0.65 0.95 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.27 1.65 0.71 ;
      RECT  1.55 0.71 1.85 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.56 0.14 1.45 0.23 ;
      RECT  0.56 0.23 0.66 0.395 ;
      RECT  1.35 0.23 1.45 0.93 ;
      RECT  0.35 0.395 0.66 0.485 ;
      RECT  0.35 0.485 0.45 0.75 ;
      RECT  0.26 0.75 0.45 0.93 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.445 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.875 1.235 1.995 1.75 ;
      RECT  2.395 1.415 2.525 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.3 0.05 0.47 0.305 ;
      RECT  2.395 0.05 2.525 0.39 ;
      RECT  1.875 0.05 1.995 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.135 0.29 2.255 0.48 ;
      RECT  2.135 0.48 2.45 0.57 ;
      RECT  2.35 0.57 2.45 1.235 ;
      RECT  2.135 1.235 2.45 1.325 ;
      RECT  2.135 1.325 2.255 1.51 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.04 0.39 1.25 0.5 ;
      RECT  1.15 0.5 1.25 1.055 ;
      RECT  1.04 1.055 2.245 1.145 ;
      RECT  2.155 0.725 2.245 1.055 ;
      RECT  0.81 0.79 1.04 0.89 ;
      RECT  0.81 0.89 0.9 1.06 ;
      RECT  0.555 1.06 0.9 1.15 ;
      RECT  0.555 1.15 0.645 1.26 ;
      RECT  0.065 0.21 0.17 1.26 ;
      RECT  0.065 1.26 0.645 1.35 ;
      RECT  0.065 1.35 0.185 1.53 ;
      RECT  0.785 1.24 1.765 1.35 ;
      RECT  0.535 1.445 1.525 1.56 ;
  END
END SEN_MUX2_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_G_3
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_G_3
  CLASS CORE ;
  FOREIGN SEN_MUX2_G_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.675 0.25 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.144 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  2.13 1.575 2.26 1.75 ;
      RECT  2.65 1.575 2.78 1.75 ;
      RECT  3.19 1.39 3.32 1.75 ;
      RECT  3.715 1.24 3.835 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  2.66 0.05 2.79 0.39 ;
      RECT  3.71 0.05 3.84 0.39 ;
      RECT  2.135 0.05 2.255 0.42 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  3.19 0.05 3.31 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.405 0.51 4.135 0.6 ;
      RECT  3.95 0.6 4.05 1.055 ;
      RECT  3.405 1.055 4.135 1.145 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.14 1.78 0.23 ;
      RECT  0.34 0.23 0.445 0.965 ;
      RECT  0.34 0.965 0.755 1.07 ;
      RECT  0.34 1.07 0.445 1.35 ;
      RECT  0.575 0.335 1.215 0.425 ;
      RECT  0.575 0.425 0.695 0.56 ;
      RECT  1.095 0.425 1.215 1.395 ;
      RECT  0.525 1.395 3.045 1.485 ;
      RECT  2.94 0.285 3.045 1.395 ;
      RECT  1.345 0.34 1.985 0.43 ;
      RECT  1.865 0.43 1.985 1.215 ;
      RECT  1.345 0.43 1.465 1.305 ;
      RECT  1.865 1.215 2.535 1.305 ;
      RECT  2.42 0.45 2.535 1.215 ;
      RECT  3.16 0.785 3.86 0.895 ;
      RECT  3.16 0.895 3.26 1.29 ;
      RECT  0.85 0.515 0.95 1.305 ;
      RECT  1.61 0.52 1.725 1.305 ;
      LAYER M2 ;
      RECT  0.81 1.15 3.3 1.25 ;
      LAYER V1 ;
      RECT  0.85 1.15 0.95 1.25 ;
      RECT  1.61 1.15 1.71 1.25 ;
      RECT  3.16 1.15 3.26 1.25 ;
  END
END SEN_MUX2_G_3
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_G_4
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_G_4
  CLASS CORE ;
  FOREIGN SEN_MUX2_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.735 ;
      RECT  1.95 0.735 2.15 0.925 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.5 2.65 0.735 ;
      RECT  2.55 0.735 2.7 0.925 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.4 0.75 1.58 0.795 ;
      RECT  1.4 0.795 1.755 0.895 ;
      RECT  0.15 0.685 0.25 1.105 ;
      LAYER M2 ;
      RECT  0.11 0.75 1.58 0.85 ;
      LAYER V1 ;
      RECT  1.44 0.75 1.54 0.85 ;
      RECT  0.15 0.75 0.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  1.93 1.44 2.06 1.75 ;
      RECT  2.455 1.21 2.575 1.75 ;
      RECT  2.97 1.41 3.1 1.75 ;
      RECT  3.495 1.24 3.615 1.75 ;
      RECT  4.015 1.21 4.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  3.49 0.05 3.62 0.36 ;
      RECT  1.93 0.05 2.06 0.39 ;
      RECT  2.45 0.05 2.575 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  2.975 0.05 3.095 0.59 ;
      RECT  4.015 0.05 4.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.185 0.455 3.86 0.545 ;
      RECT  3.75 0.545 3.86 1.055 ;
      RECT  3.185 1.055 3.86 1.145 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.665 0.23 2.88 0.32 ;
      RECT  2.79 0.32 2.88 1.015 ;
      RECT  2.72 1.015 2.88 1.1 ;
      RECT  2.72 1.1 2.82 1.49 ;
      RECT  0.85 0.17 0.95 0.35 ;
      RECT  0.695 0.35 0.95 0.45 ;
      RECT  1.04 0.24 1.785 0.36 ;
      RECT  1.04 0.36 1.13 0.55 ;
      RECT  0.525 0.55 1.13 0.64 ;
      RECT  0.67 0.64 0.76 1.105 ;
      RECT  0.59 1.105 0.76 1.29 ;
      RECT  2.18 0.31 2.34 0.49 ;
      RECT  2.25 0.49 2.34 1.235 ;
      RECT  1.305 1.235 2.34 1.35 ;
      RECT  1.22 0.45 1.525 0.57 ;
      RECT  1.22 0.57 1.31 0.81 ;
      RECT  0.85 0.81 1.31 0.9 ;
      RECT  0.85 0.9 0.95 1.51 ;
      RECT  0.34 0.325 0.43 0.755 ;
      RECT  0.34 0.755 0.58 0.925 ;
      RECT  0.34 0.925 0.43 1.41 ;
      RECT  2.97 0.79 3.64 0.89 ;
      RECT  2.97 0.89 3.07 1.31 ;
      RECT  1.105 1.0 1.785 1.12 ;
      RECT  1.105 1.12 1.205 1.31 ;
      LAYER M2 ;
      RECT  0.77 0.35 2.325 0.45 ;
      RECT  0.62 1.15 3.11 1.25 ;
      RECT  0.81 1.35 2.86 1.45 ;
      LAYER V1 ;
      RECT  0.81 0.35 0.91 0.45 ;
      RECT  2.185 0.35 2.285 0.45 ;
      RECT  0.66 1.15 0.76 1.25 ;
      RECT  1.105 1.15 1.205 1.25 ;
      RECT  2.97 1.15 3.07 1.25 ;
      RECT  0.85 1.35 0.95 1.45 ;
      RECT  2.72 1.35 2.82 1.45 ;
  END
END SEN_MUX2_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_G_6
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_G_6
  CLASS CORE ;
  FOREIGN SEN_MUX2_G_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.45 0.71 ;
      RECT  2.95 0.71 3.45 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.34 0.89 ;
      RECT  3.95 0.89 4.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.31 0.975 ;
      RECT  0.52 0.71 0.84 0.89 ;
      RECT  0.52 0.89 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.67 0.75 2.32 0.85 ;
      LAYER V1 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  0.74 0.75 0.84 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2904 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.19 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.585 1.21 0.705 1.75 ;
      RECT  2.9 1.44 3.03 1.75 ;
      RECT  3.42 1.44 3.55 1.75 ;
      RECT  3.93 1.44 4.06 1.75 ;
      RECT  4.45 1.43 4.58 1.75 ;
      RECT  4.97 1.41 5.1 1.75 ;
      RECT  5.49 1.41 5.62 1.75 ;
      RECT  6.015 1.21 6.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  3.93 0.05 4.06 0.36 ;
      RECT  2.9 0.05 3.025 0.385 ;
      RECT  3.425 0.05 3.55 0.385 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  4.97 0.05 5.1 0.39 ;
      RECT  5.49 0.05 5.62 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  4.455 0.05 4.575 0.59 ;
      RECT  6.015 0.05 6.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.715 0.51 5.86 0.69 ;
      RECT  5.73 0.69 5.86 1.11 ;
      RECT  4.73 1.11 5.86 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.12 0.255 3.335 0.345 ;
      RECT  3.12 0.345 3.21 0.475 ;
      RECT  0.85 0.14 2.75 0.23 ;
      RECT  0.85 0.23 0.94 0.39 ;
      RECT  1.37 0.23 1.46 0.39 ;
      RECT  2.66 0.23 2.75 0.475 ;
      RECT  2.66 0.475 3.21 0.565 ;
      RECT  2.66 0.565 2.75 1.055 ;
      RECT  2.41 1.055 3.335 1.145 ;
      RECT  2.41 1.145 2.5 1.36 ;
      RECT  1.825 1.36 2.5 1.48 ;
      RECT  1.59 0.32 2.305 0.41 ;
      RECT  1.59 0.41 1.68 0.48 ;
      RECT  1.11 0.32 1.2 0.48 ;
      RECT  1.11 0.48 1.68 0.57 ;
      RECT  1.19 0.57 1.28 1.11 ;
      RECT  1.095 1.11 1.28 1.29 ;
      RECT  0.34 0.29 0.43 0.53 ;
      RECT  0.34 0.53 1.02 0.62 ;
      RECT  0.93 0.62 1.02 0.96 ;
      RECT  0.34 0.62 0.43 1.45 ;
      RECT  3.65 0.455 4.365 0.545 ;
      RECT  3.65 0.545 3.74 1.255 ;
      RECT  2.72 1.255 4.365 1.345 ;
      RECT  2.72 1.345 2.81 1.57 ;
      RECT  2.41 0.335 2.5 0.5 ;
      RECT  1.85 0.5 2.5 0.59 ;
      RECT  1.85 0.59 1.94 0.885 ;
      RECT  1.37 0.885 1.94 0.975 ;
      RECT  1.37 0.975 1.46 1.57 ;
      RECT  0.83 1.37 0.955 1.57 ;
      RECT  0.83 1.57 2.81 1.66 ;
      RECT  4.53 0.785 5.64 0.895 ;
      RECT  4.53 0.895 4.63 1.31 ;
      RECT  1.565 1.115 2.28 1.205 ;
      RECT  2.1 1.205 2.28 1.25 ;
      LAYER M2 ;
      RECT  1.11 1.15 4.7 1.25 ;
      LAYER V1 ;
      RECT  1.18 1.15 1.28 1.25 ;
      RECT  2.14 1.15 2.24 1.25 ;
      RECT  4.53 1.15 4.63 1.25 ;
  END
END SEN_MUX2_G_6
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2_G_8
#      Description : "2-1 multiplexer"
#      Equation    : X=(S&D1)|(!S&D0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2_G_8
  CLASS CORE ;
  FOREIGN SEN_MUX2_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.45 0.71 ;
      RECT  3.75 0.71 4.45 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.84 0.71 5.25 0.89 ;
      RECT  5.15 0.89 5.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.19 0.71 2.29 0.785 ;
      RECT  2.19 0.785 2.63 0.89 ;
      RECT  0.52 0.71 0.84 0.89 ;
      LAYER M2 ;
      RECT  0.67 0.75 2.36 0.85 ;
      LAYER V1 ;
      RECT  2.19 0.75 2.29 0.85 ;
      RECT  0.74 0.75 0.84 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  0.58 1.39 0.71 1.75 ;
      RECT  3.27 1.44 3.38 1.75 ;
      RECT  3.77 1.44 3.9 1.75 ;
      RECT  4.29 1.44 4.42 1.75 ;
      RECT  4.81 1.44 4.94 1.75 ;
      RECT  5.33 1.41 5.46 1.75 ;
      RECT  5.85 1.41 5.98 1.75 ;
      RECT  6.37 1.41 6.5 1.75 ;
      RECT  6.89 1.41 7.02 1.75 ;
      RECT  7.415 1.21 7.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  4.81 0.05 4.94 0.36 ;
      RECT  3.27 0.05 3.38 0.385 ;
      RECT  3.77 0.05 3.9 0.385 ;
      RECT  4.29 0.05 4.42 0.385 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  5.85 0.05 5.98 0.39 ;
      RECT  6.37 0.05 6.5 0.39 ;
      RECT  6.89 0.05 7.02 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.335 0.05 5.455 0.59 ;
      RECT  7.415 0.05 7.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.51 7.275 0.69 ;
      RECT  6.68 0.69 6.85 1.11 ;
      RECT  5.61 1.11 7.285 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.09 0.14 3.18 0.23 ;
      RECT  1.09 0.23 1.18 0.385 ;
      RECT  1.61 0.23 1.7 0.385 ;
      RECT  3.09 0.23 3.18 0.475 ;
      RECT  3.09 0.475 4.205 0.565 ;
      RECT  3.09 0.565 3.18 0.84 ;
      RECT  3.53 0.565 3.62 1.055 ;
      RECT  2.72 0.84 3.18 0.93 ;
      RECT  2.72 0.93 2.81 1.36 ;
      RECT  3.53 1.055 4.205 1.145 ;
      RECT  2.065 1.36 2.81 1.48 ;
      RECT  1.8 0.32 3.0 0.41 ;
      RECT  1.8 0.41 1.89 0.53 ;
      RECT  2.895 0.41 3.0 0.54 ;
      RECT  0.765 0.53 1.89 0.62 ;
      RECT  1.42 0.62 1.52 1.145 ;
      RECT  1.205 1.145 1.52 1.16 ;
      RECT  0.765 1.16 1.52 1.25 ;
      RECT  4.57 0.455 5.245 0.545 ;
      RECT  4.57 0.545 4.66 1.255 ;
      RECT  3.09 1.255 5.245 1.345 ;
      RECT  3.09 1.345 3.18 1.57 ;
      RECT  2.01 0.5 2.805 0.59 ;
      RECT  2.01 0.59 2.1 0.885 ;
      RECT  1.61 0.885 2.1 0.975 ;
      RECT  1.61 0.975 1.7 1.57 ;
      RECT  1.07 1.37 1.195 1.57 ;
      RECT  1.07 1.57 3.18 1.66 ;
      RECT  5.41 0.785 6.57 0.895 ;
      RECT  5.41 0.895 5.51 1.29 ;
      RECT  1.015 0.755 1.305 0.93 ;
      RECT  1.015 0.93 1.105 0.98 ;
      RECT  0.325 0.29 0.43 0.98 ;
      RECT  0.325 0.98 1.105 1.07 ;
      RECT  0.325 1.07 0.43 1.45 ;
      RECT  1.805 1.115 2.52 1.205 ;
      RECT  2.34 1.205 2.52 1.25 ;
      RECT  2.9 1.03 3.0 1.47 ;
      LAYER M2 ;
      RECT  1.31 1.15 5.58 1.25 ;
      LAYER V1 ;
      RECT  1.38 1.15 1.48 1.25 ;
      RECT  2.38 1.15 2.48 1.25 ;
      RECT  2.9 1.15 3.0 1.25 ;
      RECT  5.41 1.15 5.51 1.25 ;
  END
END SEN_MUX2_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2AN2_DG_1
#      Description : "2-1 multiplexer w/and2 input"
#      Equation    : X=(S&D1)|(!S&D0A1&D0A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2AN2_DG_1
  CLASS CORE ;
  FOREIGN SEN_MUX2AN2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.415 1.85 0.505 ;
      RECT  0.75 0.505 0.875 0.89 ;
      RECT  1.75 0.505 1.85 1.035 ;
      RECT  1.59 1.035 1.85 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D0A1
  PIN D0A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D0A2
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.57 0.145 1.42 0.255 ;
      RECT  0.57 0.255 0.66 0.305 ;
      RECT  0.35 0.305 0.66 0.395 ;
      RECT  0.35 0.395 0.45 0.755 ;
      RECT  0.26 0.755 0.45 0.925 ;
      RECT  0.35 0.925 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.47 0.44 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.375 1.615 1.545 1.75 ;
      RECT  1.95 1.44 2.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.34 0.05 0.47 0.215 ;
      RECT  1.685 0.05 1.815 0.325 ;
      RECT  1.94 0.05 2.06 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.215 2.305 0.385 ;
      RECT  2.15 0.385 2.25 1.215 ;
      RECT  2.15 1.215 2.305 1.385 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.89 1.09 0.98 1.195 ;
      RECT  0.89 1.195 1.5 1.255 ;
      RECT  1.16 0.595 1.25 1.195 ;
      RECT  0.89 1.255 2.06 1.285 ;
      RECT  1.97 0.72 2.06 1.255 ;
      RECT  1.41 1.285 2.06 1.345 ;
      RECT  0.565 1.09 0.8 1.2 ;
      RECT  0.71 1.2 0.8 1.375 ;
      RECT  0.71 1.375 1.32 1.435 ;
      RECT  0.71 1.435 1.86 1.465 ;
      RECT  1.23 1.465 1.86 1.525 ;
      RECT  0.065 0.34 0.17 1.29 ;
      RECT  0.065 1.29 0.62 1.38 ;
      RECT  0.53 1.38 0.62 1.555 ;
      RECT  0.53 1.555 1.14 1.645 ;
  END
END SEN_MUX2AN2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2AN2_DG_2
#      Description : "2-1 multiplexer w/and2 input"
#      Equation    : X=(S&D1)|(!S&D0A1&D0A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2AN2_DG_2
  CLASS CORE ;
  FOREIGN SEN_MUX2AN2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.71 ;
      RECT  0.35 0.71 0.65 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0A1
  PIN D0A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0A2
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.9 ;
      RECT  1.35 0.9 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0927 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.375 0.455 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  1.415 1.63 1.585 1.75 ;
      RECT  2.27 1.45 2.44 1.75 ;
      RECT  2.815 1.21 2.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  1.105 0.05 1.22 0.36 ;
      RECT  2.81 0.05 2.94 0.385 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  2.31 0.05 2.42 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.29 2.675 0.475 ;
      RECT  2.55 0.475 2.85 0.565 ;
      RECT  2.75 0.565 2.85 1.03 ;
      RECT  2.55 1.03 2.85 1.12 ;
      RECT  2.55 1.12 2.66 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.635 0.24 2.22 0.36 ;
      RECT  2.13 0.36 2.22 0.48 ;
      RECT  2.13 0.48 2.445 0.57 ;
      RECT  2.355 0.57 2.445 0.785 ;
      RECT  2.355 0.785 2.66 0.895 ;
      RECT  2.355 0.895 2.445 1.27 ;
      RECT  0.755 0.24 1.015 0.36 ;
      RECT  0.755 0.36 0.845 1.015 ;
      RECT  0.755 1.015 0.945 1.105 ;
      RECT  0.855 1.105 0.945 1.27 ;
      RECT  0.855 1.27 2.445 1.36 ;
      RECT  0.945 0.45 2.04 0.54 ;
      RECT  1.935 0.54 2.04 0.62 ;
      RECT  0.945 0.54 1.055 0.925 ;
      RECT  1.55 0.54 1.64 1.16 ;
      RECT  0.07 1.195 0.71 1.285 ;
      RECT  0.07 1.285 0.19 1.415 ;
      RECT  0.59 1.285 0.71 1.45 ;
      RECT  0.59 1.45 1.955 1.54 ;
  END
END SEN_MUX2AN2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2AN2_DG_4
#      Description : "2-1 multiplexer w/and2 input"
#      Equation    : X=(S&D1)|(!S&D0A1&D0A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2AN2_DG_4
  CLASS CORE ;
  FOREIGN SEN_MUX2AN2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D0A1
  PIN D0A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D0A2
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.71 ;
      RECT  2.35 0.71 2.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.51 3.05 0.71 ;
      RECT  2.95 0.71 3.335 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.58 1.38 0.71 1.75 ;
      RECT  1.105 1.21 1.225 1.75 ;
      RECT  2.135 1.455 2.265 1.75 ;
      RECT  2.655 1.39 2.785 1.75 ;
      RECT  3.965 1.44 4.075 1.75 ;
      RECT  4.465 1.41 4.595 1.75 ;
      RECT  5.0 1.21 5.12 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.435 0.05 2.565 0.24 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  4.465 0.05 4.595 0.365 ;
      RECT  3.965 0.05 4.075 0.39 ;
      RECT  5.0 0.05 5.12 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.16 0.455 4.85 0.575 ;
      RECT  4.745 0.575 4.85 1.11 ;
      RECT  4.15 1.11 4.85 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.99 0.15 3.875 0.24 ;
      RECT  3.775 0.24 3.875 0.48 ;
      RECT  3.775 0.48 4.045 0.57 ;
      RECT  3.955 0.57 4.045 0.785 ;
      RECT  3.955 0.785 4.635 0.895 ;
      RECT  3.955 0.895 4.045 1.25 ;
      RECT  3.785 1.25 4.045 1.34 ;
      RECT  3.785 1.34 3.875 1.455 ;
      RECT  3.39 1.455 3.875 1.545 ;
      RECT  0.795 0.215 1.785 0.335 ;
      RECT  2.09 0.33 3.51 0.42 ;
      RECT  1.9 0.285 2.0 0.45 ;
      RECT  1.37 0.45 2.0 0.54 ;
      RECT  1.37 0.54 1.46 1.04 ;
      RECT  1.37 1.04 1.785 1.16 ;
      RECT  0.065 0.35 0.185 0.455 ;
      RECT  0.065 0.455 1.275 0.575 ;
      RECT  3.595 0.495 3.685 0.71 ;
      RECT  3.425 0.71 3.685 0.8 ;
      RECT  3.425 0.8 3.515 1.055 ;
      RECT  1.575 0.785 2.045 0.895 ;
      RECT  1.955 0.895 2.045 1.055 ;
      RECT  1.955 1.055 3.515 1.145 ;
      RECT  3.605 1.03 3.865 1.12 ;
      RECT  3.605 1.12 3.695 1.255 ;
      RECT  2.95 1.255 3.695 1.345 ;
      RECT  2.95 1.345 3.05 1.51 ;
      RECT  0.275 1.19 0.965 1.29 ;
      RECT  0.845 1.29 0.965 1.515 ;
      RECT  1.355 1.255 2.57 1.345 ;
      RECT  1.355 1.345 1.475 1.475 ;
      LAYER M2 ;
      RECT  1.83 0.35 3.95 0.45 ;
      RECT  0.78 1.35 3.12 1.45 ;
      LAYER V1 ;
      RECT  1.9 0.35 2.0 0.45 ;
      RECT  3.775 0.35 3.875 0.45 ;
      RECT  0.85 1.35 0.95 1.45 ;
      RECT  2.95 1.35 3.05 1.45 ;
  END
END SEN_MUX2AN2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2AN2_DG_8
#      Description : "2-1 multiplexer w/and2 input"
#      Equation    : X=(S&D1)|(!S&D0A1&D0A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2AN2_DG_8
  CLASS CORE ;
  FOREIGN SEN_MUX2AN2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D0A1
  PIN D0A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D0A2
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.075 0.795 4.85 0.905 ;
      RECT  4.55 0.905 4.85 1.09 ;
      RECT  4.75 1.09 4.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.71 6.45 0.795 ;
      RECT  5.35 0.795 6.45 0.905 ;
      RECT  5.55 0.905 5.65 1.09 ;
      RECT  5.35 0.905 5.45 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.58 1.38 0.71 1.75 ;
      RECT  1.1 1.38 1.23 1.75 ;
      RECT  1.62 1.38 1.75 1.75 ;
      RECT  2.14 1.39 2.255 1.75 ;
      RECT  3.68 1.415 3.81 1.75 ;
      RECT  4.2 1.43 4.33 1.75 ;
      RECT  4.72 1.39 4.85 1.75 ;
      RECT  6.525 1.415 6.65 1.75 ;
      RECT  7.04 1.41 7.17 1.75 ;
      RECT  7.56 1.41 7.69 1.75 ;
      RECT  8.08 1.41 8.21 1.75 ;
      RECT  8.615 1.21 8.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  3.92 0.05 4.09 0.305 ;
      RECT  4.44 0.05 4.61 0.305 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.835 0.05 0.97 0.385 ;
      RECT  6.54 0.05 6.65 0.39 ;
      RECT  7.04 0.05 7.17 0.39 ;
      RECT  7.56 0.05 7.69 0.39 ;
      RECT  8.08 0.05 8.21 0.39 ;
      RECT  8.615 0.05 8.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.51 8.465 0.69 ;
      RECT  7.87 0.69 8.05 1.11 ;
      RECT  6.75 1.11 8.465 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.93 0.215 6.45 0.305 ;
      RECT  6.35 0.305 6.45 0.48 ;
      RECT  6.35 0.48 6.635 0.57 ;
      RECT  6.545 0.57 6.635 0.785 ;
      RECT  6.545 0.785 7.77 0.895 ;
      RECT  6.545 0.895 6.635 1.225 ;
      RECT  6.345 1.225 6.635 1.315 ;
      RECT  6.345 1.315 6.435 1.455 ;
      RECT  5.445 1.455 6.435 1.545 ;
      RECT  1.315 0.205 3.345 0.32 ;
      RECT  3.685 0.265 3.805 0.395 ;
      RECT  3.685 0.395 6.05 0.485 ;
      RECT  3.435 0.285 3.555 0.44 ;
      RECT  2.34 0.44 3.555 0.56 ;
      RECT  2.34 0.56 2.455 1.14 ;
      RECT  2.34 1.14 3.345 1.26 ;
      RECT  0.065 0.29 0.185 0.475 ;
      RECT  0.065 0.475 2.25 0.575 ;
      RECT  2.145 0.575 2.25 0.67 ;
      RECT  6.155 0.425 6.26 0.575 ;
      RECT  3.65 0.575 6.26 0.675 ;
      RECT  3.65 0.675 3.755 0.785 ;
      RECT  4.99 0.675 5.09 1.16 ;
      RECT  2.765 0.785 3.755 0.895 ;
      RECT  6.165 1.015 6.445 1.135 ;
      RECT  6.165 1.135 6.255 1.255 ;
      RECT  4.95 1.255 6.255 1.345 ;
      RECT  4.95 1.345 5.05 1.49 ;
      RECT  0.275 1.18 2.05 1.285 ;
      RECT  1.95 1.285 2.05 1.51 ;
      RECT  3.435 1.2 4.635 1.32 ;
      RECT  3.435 1.32 3.555 1.455 ;
      RECT  2.345 1.455 3.555 1.545 ;
      LAYER M2 ;
      RECT  3.37 0.35 6.52 0.45 ;
      RECT  1.88 1.35 5.12 1.45 ;
      LAYER V1 ;
      RECT  3.445 0.35 3.545 0.45 ;
      RECT  6.35 0.35 6.45 0.45 ;
      RECT  1.95 1.35 2.05 1.45 ;
      RECT  4.95 1.35 5.05 1.45 ;
  END
END SEN_MUX2AN2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2OR2B_DG_1
#      Description : "2-1 multiplexer w/or2b input"
#      Equation    : X=(S&D1)|(!S&(!D0A|D0B))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2OR2B_DG_1
  CLASS CORE ;
  FOREIGN SEN_MUX2OR2B_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END D0A
  PIN D0B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D0B
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.63 2.25 1.145 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.745 0.49 1.98 0.69 ;
      RECT  1.745 0.69 1.85 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.39 0.45 1.75 ;
      RECT  0.0 1.75 2.8 1.85 ;
      RECT  1.02 1.6 1.19 1.75 ;
      RECT  2.29 1.415 2.42 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      RECT  0.4 0.05 0.53 0.225 ;
      RECT  0.95 0.05 1.08 0.225 ;
      RECT  2.29 0.05 2.42 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.29 2.675 0.485 ;
      RECT  2.55 0.485 2.65 0.645 ;
      RECT  2.55 0.645 2.665 0.705 ;
      RECT  2.565 0.705 2.665 0.99 ;
      RECT  2.55 0.99 2.665 1.04 ;
      RECT  2.55 1.04 2.65 1.31 ;
      RECT  2.55 1.31 2.69 1.49 ;
    END
    ANTENNADIFFAREA 0.182 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.51 0.21 1.63 0.32 ;
      RECT  0.62 0.32 1.63 0.44 ;
      RECT  1.72 0.24 2.16 0.36 ;
      RECT  2.07 0.36 2.16 0.45 ;
      RECT  2.07 0.45 2.46 0.54 ;
      RECT  2.37 0.54 2.46 0.755 ;
      RECT  2.37 0.755 2.475 0.925 ;
      RECT  2.37 0.925 2.46 1.235 ;
      RECT  2.055 1.235 2.46 1.325 ;
      RECT  2.055 1.325 2.145 1.36 ;
      RECT  1.805 1.36 2.145 1.45 ;
      RECT  1.805 1.45 1.925 1.58 ;
      RECT  0.085 0.315 0.445 0.42 ;
      RECT  0.355 0.42 0.445 0.53 ;
      RECT  0.355 0.53 0.945 0.62 ;
      RECT  0.855 0.62 0.945 0.98 ;
      RECT  0.355 0.62 0.445 1.21 ;
      RECT  0.065 1.21 0.445 1.3 ;
      RECT  0.065 1.3 0.185 1.61 ;
      RECT  1.2 0.54 1.645 0.66 ;
      RECT  1.555 0.66 1.645 1.14 ;
      RECT  1.265 1.14 1.645 1.26 ;
      RECT  0.745 1.39 1.715 1.51 ;
  END
END SEN_MUX2OR2B_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2OR2B_DG_2
#      Description : "2-1 multiplexer w/or2b input"
#      Equation    : X=(S&D1)|(!S&(!D0A|D0B))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2OR2B_DG_2
  CLASS CORE ;
  FOREIGN SEN_MUX2OR2B_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.675 0.25 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END D0A
  PIN D0B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0B
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.66 2.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.76 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0927 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.43 0.45 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.07 1.615 1.24 1.75 ;
      RECT  2.49 1.44 2.62 1.75 ;
      RECT  3.015 1.21 3.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.88 0.05 1.01 0.225 ;
      RECT  2.49 0.05 2.62 0.39 ;
      RECT  3.01 0.05 3.14 0.39 ;
      RECT  0.32 0.05 0.445 0.405 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.31 2.875 0.51 ;
      RECT  2.75 0.51 3.05 0.6 ;
      RECT  2.95 0.6 3.05 1.02 ;
      RECT  2.75 1.02 3.05 1.11 ;
      RECT  2.75 1.11 2.86 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.535 0.315 1.595 0.405 ;
      RECT  1.685 0.31 1.805 0.48 ;
      RECT  1.685 0.48 2.66 0.57 ;
      RECT  2.57 0.57 2.66 0.785 ;
      RECT  2.57 0.785 2.845 0.895 ;
      RECT  2.57 0.895 2.66 1.26 ;
      RECT  1.945 1.26 2.66 1.35 ;
      RECT  1.945 1.35 2.065 1.51 ;
      RECT  0.065 0.21 0.185 0.495 ;
      RECT  0.065 0.495 0.845 0.585 ;
      RECT  0.755 0.585 0.845 1.23 ;
      RECT  0.065 1.23 0.845 1.32 ;
      RECT  0.065 1.32 0.185 1.61 ;
      RECT  1.105 0.55 1.47 0.67 ;
      RECT  1.38 0.67 1.47 0.745 ;
      RECT  1.38 0.745 2.195 0.855 ;
      RECT  1.38 0.855 1.485 1.345 ;
      RECT  1.685 1.065 1.805 1.435 ;
      RECT  0.795 1.435 1.805 1.525 ;
  END
END SEN_MUX2OR2B_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2OR2B_DG_4
#      Description : "2-1 multiplexer w/or2b input"
#      Equation    : X=(S&D1)|(!S&(!D0A|D0B))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2OR2B_DG_4
  CLASS CORE ;
  FOREIGN SEN_MUX2OR2B_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.55 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D0A
  PIN D0B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D0B
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.82 4.25 0.94 ;
      RECT  3.75 0.94 3.85 1.09 ;
      RECT  4.15 0.94 4.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.115 0.71 3.45 0.9 ;
      RECT  1.945 0.75 2.755 0.85 ;
      RECT  1.945 0.85 2.055 1.09 ;
      LAYER M2 ;
      RECT  2.52 0.75 3.29 0.85 ;
      LAYER V1 ;
      RECT  3.15 0.75 3.25 0.85 ;
      RECT  2.59 0.75 2.69 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.39 0.45 1.75 ;
      RECT  0.0 1.75 5.4 1.85 ;
      RECT  1.71 1.43 1.83 1.75 ;
      RECT  3.615 1.44 3.745 1.75 ;
      RECT  4.135 1.39 4.265 1.75 ;
      RECT  4.655 1.39 4.785 1.75 ;
      RECT  5.215 1.21 5.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      RECT  3.615 0.05 3.745 0.36 ;
      RECT  4.665 0.05 4.795 0.365 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.765 0.05 1.89 0.39 ;
      RECT  1.1 0.05 1.21 0.41 ;
      RECT  4.14 0.05 4.26 0.545 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.215 0.05 5.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.36 0.455 5.05 0.545 ;
      RECT  4.95 0.545 5.05 1.11 ;
      RECT  4.35 1.11 5.05 1.29 ;
    END
    ANTENNADIFFAREA 0.47 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.065 0.14 2.34 0.23 ;
      RECT  2.065 0.23 2.155 0.48 ;
      RECT  1.305 0.14 1.415 0.32 ;
      RECT  1.305 0.32 1.675 0.41 ;
      RECT  3.06 0.455 4.05 0.545 ;
      RECT  0.275 0.5 1.975 0.57 ;
      RECT  0.275 0.57 2.76 0.62 ;
      RECT  1.885 0.62 2.76 0.66 ;
      RECT  3.555 0.64 4.445 0.73 ;
      RECT  4.355 0.73 4.445 0.785 ;
      RECT  3.555 0.73 3.645 1.03 ;
      RECT  4.355 0.785 4.83 0.895 ;
      RECT  2.865 0.255 3.525 0.345 ;
      RECT  2.865 0.345 2.955 0.385 ;
      RECT  2.28 0.385 2.955 0.48 ;
      RECT  2.865 0.48 2.955 1.03 ;
      RECT  2.28 1.03 3.645 1.12 ;
      RECT  0.6 1.03 1.275 1.12 ;
      RECT  0.6 1.12 0.69 1.19 ;
      RECT  0.065 1.19 0.69 1.3 ;
      RECT  0.065 1.3 0.185 1.41 ;
      RECT  0.795 1.25 3.28 1.34 ;
      RECT  3.37 1.255 4.05 1.345 ;
      RECT  3.37 1.345 3.46 1.455 ;
      RECT  2.54 1.455 3.46 1.545 ;
      RECT  1.12 1.48 1.62 1.57 ;
      RECT  1.92 1.48 2.445 1.57 ;
  END
END SEN_MUX2OR2B_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX2OR2B_DG_8
#      Description : "2-1 multiplexer w/or2b input"
#      Equation    : X=(S&D1)|(!S&(!D0A|D0B))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX2OR2B_DG_8
  CLASS CORE ;
  FOREIGN SEN_MUX2OR2B_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 2.65 0.99 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0A
  PIN D0B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D0B
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.84 0.815 6.65 0.925 ;
      RECT  6.15 0.925 6.25 1.09 ;
      RECT  6.55 0.925 6.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.505 0.71 5.05 0.89 ;
      RECT  2.75 0.51 2.85 0.71 ;
      RECT  2.75 0.71 2.93 0.9 ;
      RECT  2.75 0.9 2.85 1.09 ;
      LAYER M2 ;
      RECT  2.76 0.75 4.92 0.85 ;
      LAYER V1 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  2.83 0.75 2.93 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.39 0.45 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.84 1.39 0.97 1.75 ;
      RECT  2.65 1.495 2.82 1.75 ;
      RECT  5.49 1.43 5.62 1.75 ;
      RECT  6.01 1.43 6.14 1.75 ;
      RECT  6.53 1.415 6.66 1.75 ;
      RECT  7.05 1.39 7.18 1.75 ;
      RECT  7.57 1.39 7.7 1.75 ;
      RECT  8.09 1.39 8.22 1.75 ;
      RECT  8.615 1.21 8.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  7.05 0.05 7.18 0.345 ;
      RECT  5.5 0.05 5.62 0.36 ;
      RECT  6.01 0.05 6.14 0.36 ;
      RECT  0.58 0.05 0.71 0.37 ;
      RECT  1.1 0.05 1.23 0.37 ;
      RECT  1.62 0.05 1.75 0.37 ;
      RECT  7.57 0.05 7.7 0.39 ;
      RECT  8.09 0.05 8.22 0.39 ;
      RECT  2.675 0.05 2.795 0.41 ;
      RECT  6.535 0.05 6.655 0.545 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  8.615 0.05 8.735 0.59 ;
      RECT  2.145 0.05 2.265 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.745 0.435 7.15 0.51 ;
      RECT  6.745 0.51 8.475 0.545 ;
      RECT  7.05 0.545 8.475 0.69 ;
      RECT  7.88 0.69 8.05 1.11 ;
      RECT  6.75 1.11 8.475 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.365 0.24 2.585 0.36 ;
      RECT  2.365 0.36 2.455 0.785 ;
      RECT  1.485 0.785 2.455 0.895 ;
      RECT  2.365 0.895 2.455 1.08 ;
      RECT  2.365 1.08 2.565 1.19 ;
      RECT  2.885 0.24 3.11 0.36 ;
      RECT  3.02 0.36 3.11 0.785 ;
      RECT  3.02 0.785 4.03 0.895 ;
      RECT  3.02 0.895 3.11 0.99 ;
      RECT  2.94 0.99 3.11 1.16 ;
      RECT  3.395 0.35 4.135 0.45 ;
      RECT  1.95 0.29 2.05 0.47 ;
      RECT  0.275 0.47 2.05 0.59 ;
      RECT  4.46 0.455 6.445 0.545 ;
      RECT  5.415 0.635 6.905 0.725 ;
      RECT  6.815 0.725 6.905 0.785 ;
      RECT  5.415 0.725 5.525 1.04 ;
      RECT  6.815 0.785 7.76 0.895 ;
      RECT  4.225 0.24 5.41 0.36 ;
      RECT  4.225 0.36 4.345 0.54 ;
      RECT  3.2 0.29 3.305 0.54 ;
      RECT  3.2 0.54 4.345 0.64 ;
      RECT  4.24 0.64 4.345 1.04 ;
      RECT  3.2 1.04 5.525 1.16 ;
      RECT  3.2 1.16 3.305 1.225 ;
      RECT  2.145 1.04 2.265 1.18 ;
      RECT  0.065 1.18 2.265 1.29 ;
      RECT  0.065 1.29 0.185 1.51 ;
      RECT  5.275 1.25 6.445 1.34 ;
      RECT  5.275 1.34 5.365 1.495 ;
      RECT  3.39 1.495 5.365 1.585 ;
      RECT  2.43 1.315 5.18 1.405 ;
      RECT  2.43 1.405 2.52 1.455 ;
      RECT  1.315 1.455 2.52 1.575 ;
      LAYER M2 ;
      RECT  1.88 0.35 3.63 0.45 ;
      LAYER V1 ;
      RECT  1.95 0.35 2.05 0.45 ;
      RECT  3.46 0.35 3.56 0.45 ;
  END
END SEN_MUX2OR2B_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX3_DG_1
#      Description : "3-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX3_DG_1
  CLASS CORE ;
  FOREIGN SEN_MUX3_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.69 0.595 0.885 ;
      RECT  0.35 0.885 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.485 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END D2
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.685 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.625 ;
      RECT  1.35 0.625 1.5 0.8 ;
      RECT  1.35 0.8 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.205 1.2 1.4 1.32 ;
      RECT  1.31 1.32 1.4 1.75 ;
      RECT  0.33 1.4 0.46 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  2.665 1.41 2.795 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  2.665 0.05 2.795 0.345 ;
      RECT  1.25 0.05 1.38 0.385 ;
      RECT  0.32 0.05 0.45 0.405 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.31 3.06 1.49 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.49 0.215 2.05 0.335 ;
      RECT  1.96 0.335 2.05 0.895 ;
      RECT  1.59 0.335 1.68 1.18 ;
      RECT  1.96 0.895 2.1 1.065 ;
      RECT  1.49 1.18 1.68 1.27 ;
      RECT  0.735 0.24 1.05 0.36 ;
      RECT  0.95 0.36 1.05 1.215 ;
      RECT  0.78 1.215 1.05 1.305 ;
      RECT  0.78 1.305 0.96 1.45 ;
      RECT  2.37 0.215 2.505 0.385 ;
      RECT  2.37 0.385 2.46 1.59 ;
      RECT  0.065 0.2 0.185 0.495 ;
      RECT  0.065 0.495 0.835 0.585 ;
      RECT  0.065 0.585 0.185 1.22 ;
      RECT  0.065 1.22 0.655 1.31 ;
      RECT  0.565 1.31 0.655 1.555 ;
      RECT  0.565 1.555 1.085 1.645 ;
      RECT  2.14 0.19 2.24 0.605 ;
      RECT  2.14 0.605 2.28 0.695 ;
      RECT  2.19 0.695 2.28 1.185 ;
      RECT  2.03 1.185 2.28 1.275 ;
      RECT  2.03 1.275 2.15 1.61 ;
      RECT  2.75 0.435 2.85 0.98 ;
      RECT  1.77 0.455 1.87 1.605 ;
      LAYER M2 ;
      RECT  2.1 0.55 2.89 0.65 ;
      RECT  0.78 1.35 1.91 1.45 ;
      LAYER V1 ;
      RECT  2.14 0.55 2.24 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  0.82 1.35 0.92 1.45 ;
      RECT  1.77 1.35 1.87 1.45 ;
  END
END SEN_MUX3_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX3_DG_2
#      Description : "3-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX3_DG_2
  CLASS CORE ;
  FOREIGN SEN_MUX3_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.84 ;
      RECT  0.35 0.84 0.65 0.93 ;
      RECT  0.55 0.93 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.51 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END D2
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 1.04 0.35 1.255 ;
      RECT  0.26 1.255 0.85 1.345 ;
      RECT  0.75 0.815 0.85 1.255 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0603 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  1.38 1.39 1.51 1.75 ;
      RECT  3.1 1.44 3.23 1.75 ;
      RECT  3.62 1.44 3.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  1.38 0.05 1.51 0.24 ;
      RECT  3.62 0.05 3.745 0.365 ;
      RECT  3.1 0.05 3.23 0.39 ;
      RECT  0.32 0.05 0.45 0.43 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.315 0.455 3.65 0.575 ;
      RECT  3.55 0.575 3.65 1.225 ;
      RECT  3.34 1.225 3.65 1.345 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.9 0.14 2.755 0.23 ;
      RECT  1.9 0.23 1.99 0.33 ;
      RECT  0.74 0.33 1.99 0.42 ;
      RECT  1.455 0.42 1.545 1.18 ;
      RECT  1.9 0.42 1.99 1.185 ;
      RECT  1.15 1.18 1.545 1.27 ;
      RECT  1.15 1.27 1.25 1.44 ;
      RECT  0.79 1.44 1.25 1.56 ;
      RECT  2.845 0.2 2.965 0.32 ;
      RECT  2.08 0.32 2.965 0.41 ;
      RECT  2.08 0.41 2.185 0.6 ;
      RECT  2.725 0.41 2.845 1.16 ;
      RECT  0.065 0.27 0.185 0.53 ;
      RECT  0.065 0.53 1.045 0.62 ;
      RECT  0.665 0.62 0.835 0.67 ;
      RECT  0.955 0.62 1.045 1.25 ;
      RECT  0.065 0.62 0.17 1.61 ;
      RECT  3.155 0.795 3.44 0.885 ;
      RECT  3.155 0.885 3.245 1.25 ;
      RECT  2.34 0.5 2.445 1.25 ;
      RECT  2.34 1.25 3.245 1.34 ;
      RECT  1.665 0.51 1.785 1.57 ;
      RECT  1.665 1.57 2.585 1.66 ;
      RECT  2.495 1.43 2.585 1.57 ;
  END
END SEN_MUX3_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX3_DG_3
#      Description : "3-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX3_DG_3
  CLASS CORE ;
  FOREIGN SEN_MUX3_DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.515 0.71 0.65 0.965 ;
      RECT  0.55 0.965 0.65 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.05 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END D2
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.255 1.11 ;
      RECT  0.75 0.91 0.85 1.49 ;
      RECT  0.26 0.635 0.36 1.09 ;
      LAYER M2 ;
      RECT  0.19 0.95 1.32 1.05 ;
      LAYER V1 ;
      RECT  1.15 0.95 1.25 1.05 ;
      RECT  0.75 0.95 0.85 1.05 ;
      RECT  0.26 0.95 0.36 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0759 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.605 ;
      RECT  2.35 0.605 2.535 0.775 ;
      RECT  2.35 0.775 2.45 0.89 ;
      RECT  1.55 0.51 1.65 0.71 ;
      RECT  1.55 0.71 2.05 0.89 ;
      LAYER M2 ;
      RECT  1.91 0.75 2.52 0.85 ;
      LAYER V1 ;
      RECT  2.35 0.75 2.45 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0759 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.39 0.46 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  1.49 1.44 1.62 1.75 ;
      RECT  3.02 1.455 3.19 1.75 ;
      RECT  3.56 1.44 3.69 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  1.49 0.05 1.6 0.24 ;
      RECT  0.315 0.05 0.485 0.36 ;
      RECT  3.04 0.05 3.17 0.36 ;
      RECT  3.56 0.05 3.69 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.32 0.29 3.45 0.455 ;
      RECT  3.32 0.455 3.945 0.545 ;
      RECT  3.825 0.19 3.945 0.455 ;
      RECT  3.75 0.545 3.85 1.255 ;
      RECT  3.32 1.255 3.945 1.345 ;
      RECT  3.32 1.345 3.45 1.51 ;
      RECT  3.825 1.345 3.945 1.61 ;
    END
    ANTENNADIFFAREA 0.356 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.295 0.23 2.95 0.32 ;
      RECT  2.86 0.32 2.95 0.45 ;
      RECT  2.86 0.45 3.23 0.54 ;
      RECT  3.14 0.54 3.23 0.795 ;
      RECT  3.14 0.795 3.64 0.885 ;
      RECT  3.14 0.885 3.23 1.255 ;
      RECT  2.295 1.255 3.23 1.345 ;
      RECT  1.69 0.255 2.19 0.33 ;
      RECT  0.955 0.33 2.19 0.345 ;
      RECT  0.955 0.345 1.78 0.42 ;
      RECT  2.1 0.345 2.19 0.43 ;
      RECT  0.955 0.42 1.045 1.26 ;
      RECT  0.955 1.26 2.205 1.35 ;
      RECT  0.075 0.23 0.17 0.45 ;
      RECT  0.075 0.45 0.845 0.54 ;
      RECT  0.755 0.54 0.845 0.815 ;
      RECT  0.075 0.54 0.17 1.59 ;
      RECT  1.87 0.435 1.96 0.52 ;
      RECT  1.87 0.52 2.245 0.61 ;
      RECT  2.155 0.61 2.245 0.995 ;
      RECT  1.79 0.995 2.565 1.085 ;
      RECT  1.79 1.085 1.88 1.17 ;
      RECT  2.655 0.41 2.745 1.16 ;
  END
END SEN_MUX3_DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX3_DG_4
#      Description : "3-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX3_DG_4
  CLASS CORE ;
  FOREIGN SEN_MUX3_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.61 2.45 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D2
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
      RECT  0.15 0.71 0.275 1.09 ;
      LAYER M2 ;
      RECT  0.105 0.75 1.52 0.85 ;
      LAYER V1 ;
      RECT  1.35 0.75 1.45 0.85 ;
      RECT  0.175 0.75 0.275 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.75 0.93 ;
      RECT  2.55 0.93 2.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.97 1.42 2.1 1.75 ;
      RECT  2.48 1.39 2.61 1.75 ;
      RECT  3.77 1.415 3.9 1.75 ;
      RECT  4.29 1.415 4.42 1.75 ;
      RECT  4.815 1.21 4.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  2.48 0.05 2.61 0.235 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  1.835 0.05 1.965 0.39 ;
      RECT  3.77 0.05 3.9 0.39 ;
      RECT  4.29 0.05 4.42 0.39 ;
      RECT  4.815 0.05 4.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.035 0.29 4.155 0.48 ;
      RECT  4.035 0.48 4.675 0.59 ;
      RECT  4.55 0.29 4.675 0.48 ;
      RECT  4.55 0.59 4.675 1.215 ;
      RECT  4.05 1.215 4.675 1.305 ;
      RECT  4.05 1.305 4.14 1.44 ;
      RECT  4.55 1.305 4.675 1.515 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.015 0.165 3.115 0.325 ;
      RECT  2.155 0.325 3.115 0.415 ;
      RECT  2.155 0.415 2.255 1.255 ;
      RECT  2.155 1.255 2.37 1.345 ;
      RECT  3.525 0.15 3.645 0.35 ;
      RECT  3.4 0.35 3.645 0.45 ;
      RECT  0.065 0.165 0.185 0.53 ;
      RECT  0.065 0.53 1.02 0.62 ;
      RECT  0.93 0.62 1.02 0.955 ;
      RECT  0.365 0.62 0.455 1.235 ;
      RECT  0.065 1.235 0.455 1.325 ;
      RECT  0.065 1.325 0.185 1.53 ;
      RECT  2.72 0.505 3.19 0.595 ;
      RECT  3.09 0.595 3.19 0.92 ;
      RECT  2.84 0.92 3.19 1.01 ;
      RECT  2.84 1.01 2.93 1.455 ;
      RECT  2.7 1.455 2.93 1.545 ;
      RECT  3.68 0.55 3.89 0.65 ;
      RECT  3.68 0.65 3.78 1.055 ;
      RECT  3.5 1.055 3.78 1.145 ;
      RECT  3.87 0.795 4.46 0.885 ;
      RECT  3.87 0.885 3.96 1.235 ;
      RECT  3.28 0.535 3.37 1.235 ;
      RECT  3.28 1.235 3.96 1.325 ;
      RECT  3.46 0.54 3.58 0.965 ;
      RECT  1.11 0.285 1.21 1.29 ;
      RECT  1.3 1.205 1.885 1.325 ;
      RECT  1.3 1.325 1.39 1.39 ;
      RECT  0.795 1.39 1.39 1.48 ;
      RECT  0.585 1.415 0.705 1.57 ;
      RECT  0.585 1.57 1.585 1.66 ;
      RECT  1.48 1.415 1.585 1.57 ;
      RECT  3.02 1.1 3.12 1.6 ;
      LAYER M2 ;
      RECT  1.04 0.35 3.63 0.45 ;
      RECT  2.115 0.55 3.92 0.65 ;
      RECT  3.02 0.75 3.63 0.85 ;
      RECT  1.07 1.15 3.19 1.25 ;
      LAYER V1 ;
      RECT  1.11 0.35 1.21 0.45 ;
      RECT  3.44 0.35 3.54 0.45 ;
      RECT  2.155 0.55 2.255 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  3.09 0.75 3.19 0.85 ;
      RECT  3.46 0.75 3.56 0.85 ;
      RECT  1.11 1.15 1.21 1.25 ;
      RECT  3.02 1.15 3.12 1.25 ;
  END
END SEN_MUX3_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX3_DG_6
#      Description : "3-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX3_DG_6
  CLASS CORE ;
  FOREIGN SEN_MUX3_DG_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.905 ;
      RECT  0.95 0.905 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  2.15 0.91 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.615 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END D2
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.61 3.05 1.31 ;
      RECT  1.55 0.91 1.65 1.36 ;
      RECT  0.15 0.51 0.25 1.29 ;
      LAYER M2 ;
      RECT  0.08 1.15 3.12 1.25 ;
      LAYER V1 ;
      RECT  2.95 1.15 3.05 1.25 ;
      RECT  1.55 1.15 1.65 1.25 ;
      RECT  0.15 1.15 0.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.144 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.51 4.05 0.79 ;
      RECT  3.95 0.79 4.19 0.96 ;
      RECT  3.95 0.96 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.144 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.83 1.455 0.96 1.75 ;
      RECT  2.14 1.44 2.25 1.75 ;
      RECT  3.505 1.455 3.635 1.75 ;
      RECT  4.02 1.21 4.14 1.75 ;
      RECT  6.06 1.21 6.165 1.75 ;
      RECT  6.56 1.39 6.69 1.75 ;
      RECT  7.08 1.39 7.21 1.75 ;
      RECT  7.615 1.21 7.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  2.18 0.05 2.27 0.255 ;
      RECT  0.83 0.05 0.96 0.345 ;
      RECT  3.505 0.05 3.635 0.345 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  4.02 0.05 4.145 0.39 ;
      RECT  6.56 0.05 6.69 0.42 ;
      RECT  7.08 0.05 7.21 0.42 ;
      RECT  6.06 0.05 6.165 0.59 ;
      RECT  7.615 0.05 7.735 0.59 ;
      RECT  2.1 0.255 2.27 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.305 0.51 7.465 0.69 ;
      RECT  7.12 0.69 7.25 1.11 ;
      RECT  6.28 1.11 7.465 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.11 0.14 1.72 0.23 ;
      RECT  1.63 0.23 1.72 0.385 ;
      RECT  1.11 0.23 1.2 0.435 ;
      RECT  0.545 0.435 1.2 0.525 ;
      RECT  2.49 0.14 3.105 0.23 ;
      RECT  2.49 0.23 2.58 0.255 ;
      RECT  3.015 0.23 3.105 0.47 ;
      RECT  2.36 0.255 2.58 0.345 ;
      RECT  2.36 0.345 2.45 0.435 ;
      RECT  1.865 0.205 1.985 0.435 ;
      RECT  1.865 0.435 2.45 0.525 ;
      RECT  4.28 0.145 5.45 0.245 ;
      RECT  4.28 0.245 4.4 1.51 ;
      RECT  3.745 0.235 3.915 0.355 ;
      RECT  3.745 0.355 3.835 0.435 ;
      RECT  3.265 0.315 3.355 0.435 ;
      RECT  3.265 0.435 3.835 0.525 ;
      RECT  3.265 0.525 3.355 1.275 ;
      RECT  3.265 1.275 3.85 1.29 ;
      RECT  3.75 1.09 3.85 1.275 ;
      RECT  3.265 1.29 3.89 1.365 ;
      RECT  3.77 1.365 3.89 1.51 ;
      RECT  1.29 0.35 1.47 0.45 ;
      RECT  1.37 0.45 1.46 1.34 ;
      RECT  2.745 0.35 2.925 0.45 ;
      RECT  2.745 0.45 2.845 1.335 ;
      RECT  4.985 0.35 5.63 0.45 ;
      RECT  4.985 0.45 5.075 0.97 ;
      RECT  4.985 0.97 5.79 1.06 ;
      RECT  5.7 1.06 5.79 1.35 ;
      RECT  4.75 1.35 5.79 1.47 ;
      RECT  5.165 0.54 5.97 0.66 ;
      RECT  5.88 0.66 5.97 0.785 ;
      RECT  5.88 0.785 7.01 0.895 ;
      RECT  5.88 0.895 5.97 1.56 ;
      RECT  4.545 0.37 4.66 1.56 ;
      RECT  4.545 1.56 5.97 1.66 ;
      RECT  1.55 0.51 1.65 0.71 ;
      RECT  1.55 0.71 1.86 0.8 ;
      RECT  4.805 0.37 4.895 1.15 ;
      RECT  4.805 1.15 5.605 1.26 ;
      RECT  2.55 0.49 2.65 1.165 ;
      RECT  1.95 1.255 2.61 1.345 ;
      RECT  1.95 1.345 2.05 1.415 ;
      RECT  2.52 1.345 2.61 1.455 ;
      RECT  1.865 1.415 2.05 1.585 ;
      RECT  2.52 1.455 3.17 1.545 ;
      RECT  0.54 1.24 1.265 1.36 ;
      RECT  1.175 1.36 1.265 1.46 ;
      RECT  1.175 1.46 1.76 1.58 ;
      RECT  0.34 0.29 0.45 1.41 ;
      LAYER M2 ;
      RECT  1.26 0.35 5.33 0.45 ;
      RECT  0.31 0.55 2.72 0.65 ;
      RECT  3.68 1.15 5.085 1.25 ;
      LAYER V1 ;
      RECT  1.33 0.35 1.43 0.45 ;
      RECT  2.785 0.35 2.885 0.45 ;
      RECT  5.19 0.35 5.29 0.45 ;
      RECT  0.35 0.55 0.45 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  2.55 0.55 2.65 0.65 ;
      RECT  3.75 1.15 3.85 1.25 ;
      RECT  4.945 1.15 5.045 1.25 ;
  END
END SEN_MUX3_DG_6
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX4_0P5
#      Description : "4-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX4_0P5
  CLASS CORE ;
  FOREIGN SEN_MUX4_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.86 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0264 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.625 0.71 2.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0264 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.515 0.685 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0264 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.67 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0264 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 1.85 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.215 0.91 4.45 1.14 ;
      RECT  4.35 1.14 4.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0396 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.58 1.19 0.71 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  1.67 1.43 1.795 1.75 ;
      RECT  2.74 1.185 2.87 1.75 ;
      RECT  4.35 1.415 4.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  1.62 0.05 1.79 0.17 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  4.35 0.05 4.48 0.6 ;
      RECT  2.74 0.05 2.87 0.605 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.615 0.405 4.72 0.71 ;
      RECT  4.55 0.71 4.72 0.8 ;
      RECT  4.55 0.8 4.65 1.2 ;
      RECT  4.55 1.2 4.72 1.29 ;
      RECT  4.615 1.29 4.72 1.53 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.01 0.14 4.1 0.22 ;
      RECT  3.58 0.22 4.1 0.31 ;
      RECT  3.58 0.31 3.67 1.39 ;
      RECT  1.88 0.14 2.53 0.235 ;
      RECT  1.88 0.235 1.97 0.26 ;
      RECT  1.335 0.26 1.97 0.38 ;
      RECT  1.335 0.38 1.425 1.455 ;
      RECT  1.335 1.455 1.58 1.575 ;
      RECT  0.055 0.31 0.24 0.49 ;
      RECT  0.055 0.49 0.175 1.38 ;
      RECT  0.805 0.435 1.04 0.56 ;
      RECT  0.95 0.56 1.04 1.23 ;
      RECT  0.805 1.23 1.04 1.35 ;
      RECT  4.03 0.405 4.175 0.575 ;
      RECT  4.03 0.575 4.12 1.23 ;
      RECT  4.03 1.23 4.2 1.32 ;
      RECT  4.11 1.32 4.2 1.56 ;
      RECT  3.4 1.56 4.2 1.66 ;
      RECT  2.985 0.46 3.23 0.58 ;
      RECT  3.14 0.58 3.23 1.235 ;
      RECT  2.985 1.235 3.23 1.355 ;
      RECT  1.53 0.505 2.06 0.61 ;
      RECT  1.94 0.61 2.06 0.7 ;
      RECT  1.53 0.61 1.62 1.25 ;
      RECT  1.53 1.25 2.035 1.34 ;
      RECT  1.945 1.34 2.035 1.57 ;
      RECT  1.945 1.57 2.53 1.66 ;
      RECT  2.43 0.43 2.535 1.215 ;
      RECT  2.43 1.215 2.6 1.305 ;
      RECT  2.165 0.435 2.28 1.35 ;
      RECT  2.165 1.35 2.345 1.45 ;
      RECT  3.825 0.435 3.94 1.35 ;
      RECT  3.76 1.35 3.94 1.45 ;
      RECT  3.32 0.29 3.42 1.39 ;
      RECT  0.33 0.42 0.425 1.4 ;
      RECT  1.13 0.41 1.235 1.51 ;
      LAYER M2 ;
      RECT  0.07 0.35 3.49 0.45 ;
      RECT  1.09 1.35 3.97 1.45 ;
      LAYER V1 ;
      RECT  0.14 0.35 0.24 0.45 ;
      RECT  3.32 0.35 3.42 0.45 ;
      RECT  1.13 1.35 1.23 1.45 ;
      RECT  2.205 1.35 2.305 1.45 ;
      RECT  3.8 1.35 3.9 1.45 ;
  END
END SEN_MUX4_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX4_3
#      Description : "4-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX4_3
  CLASS CORE ;
  FOREIGN SEN_MUX4_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.7 3.65 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.45 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.06 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.805 0.71 7.05 0.915 ;
      RECT  6.95 0.915 7.05 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.093 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 8.0 1.85 ;
      RECT  1.095 1.42 1.225 1.75 ;
      RECT  2.66 1.415 2.79 1.75 ;
      RECT  3.41 1.48 3.58 1.75 ;
      RECT  5.02 1.45 5.15 1.75 ;
      RECT  6.92 1.215 7.04 1.75 ;
      RECT  7.515 1.415 7.645 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      RECT  1.095 0.05 1.225 0.345 ;
      RECT  5.0 0.05 5.17 0.35 ;
      RECT  2.66 0.05 2.79 0.36 ;
      RECT  3.43 0.05 3.56 0.36 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  7.515 0.05 7.645 0.415 ;
      RECT  6.935 0.05 7.055 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.51 7.92 0.69 ;
      RECT  7.75 0.69 7.85 1.11 ;
      RECT  7.15 1.11 7.92 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.93 0.14 2.51 0.23 ;
      RECT  1.93 0.23 2.02 0.315 ;
      RECT  2.42 0.23 2.51 0.45 ;
      RECT  1.85 0.315 2.02 0.42 ;
      RECT  2.42 0.45 3.045 0.54 ;
      RECT  2.94 0.54 3.045 1.225 ;
      RECT  2.355 1.225 3.045 1.315 ;
      RECT  5.39 0.14 6.715 0.235 ;
      RECT  6.61 0.235 6.715 1.315 ;
      RECT  4.2 0.15 4.87 0.27 ;
      RECT  4.78 0.27 4.87 0.44 ;
      RECT  4.78 0.44 5.455 0.56 ;
      RECT  4.78 0.56 4.87 1.24 ;
      RECT  4.78 1.24 5.455 1.36 ;
      RECT  3.91 0.19 4.08 0.36 ;
      RECT  3.91 0.36 4.01 1.135 ;
      RECT  3.91 1.135 4.06 1.225 ;
      RECT  3.97 1.225 4.06 1.41 ;
      RECT  3.705 0.165 3.8 0.45 ;
      RECT  3.175 0.45 3.8 0.54 ;
      RECT  3.175 0.54 3.28 1.3 ;
      RECT  3.175 1.3 3.815 1.39 ;
      RECT  3.695 1.39 3.815 1.5 ;
      RECT  3.695 1.5 4.37 1.59 ;
      RECT  4.2 1.48 4.37 1.5 ;
      RECT  0.065 0.345 0.185 0.51 ;
      RECT  0.065 0.51 0.51 0.6 ;
      RECT  0.41 0.6 0.51 1.23 ;
      RECT  0.065 1.23 0.51 1.32 ;
      RECT  0.065 1.32 0.185 1.45 ;
      RECT  5.765 0.395 5.975 0.515 ;
      RECT  5.765 0.515 5.855 1.35 ;
      RECT  5.765 1.35 5.975 1.475 ;
      RECT  6.285 0.35 6.48 0.52 ;
      RECT  6.36 0.52 6.48 1.38 ;
      RECT  0.835 0.435 1.535 0.555 ;
      RECT  0.835 0.555 0.955 1.24 ;
      RECT  0.835 1.24 1.485 1.33 ;
      RECT  1.365 1.33 1.485 1.5 ;
      RECT  1.365 1.5 2.04 1.59 ;
      RECT  1.87 1.465 2.04 1.5 ;
      RECT  1.84 0.51 2.06 0.705 ;
      RECT  1.855 0.85 2.03 0.95 ;
      RECT  1.93 0.95 2.03 1.29 ;
      RECT  4.1 0.51 4.2 1.01 ;
      RECT  4.29 0.57 4.39 1.31 ;
      RECT  0.6 0.29 0.7 1.315 ;
      RECT  1.63 0.165 1.75 1.41 ;
      RECT  2.15 0.32 2.255 1.51 ;
      RECT  4.51 0.375 4.61 1.52 ;
      RECT  6.1 0.37 6.195 1.56 ;
      RECT  6.1 1.56 6.7 1.565 ;
      RECT  5.57 0.37 5.675 1.565 ;
      RECT  5.57 1.565 6.7 1.66 ;
      LAYER M2 ;
      RECT  1.61 0.35 6.5 0.45 ;
      RECT  0.37 0.55 4.24 0.65 ;
      RECT  0.56 1.15 4.43 1.25 ;
      RECT  2.115 1.35 5.945 1.45 ;
      LAYER V1 ;
      RECT  1.65 0.35 1.75 0.45 ;
      RECT  3.91 0.35 4.01 0.45 ;
      RECT  6.325 0.35 6.425 0.45 ;
      RECT  0.41 0.55 0.51 0.65 ;
      RECT  1.9 0.55 2.0 0.65 ;
      RECT  4.1 0.55 4.2 0.65 ;
      RECT  0.6 1.15 0.7 1.25 ;
      RECT  1.93 1.15 2.03 1.25 ;
      RECT  4.29 1.15 4.39 1.25 ;
      RECT  2.155 1.35 2.255 1.45 ;
      RECT  4.51 1.35 4.61 1.45 ;
      RECT  5.805 1.35 5.905 1.45 ;
  END
END SEN_MUX4_3
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX4_D_1
#      Description : "4-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX4_D_1
  CLASS CORE ;
  FOREIGN SEN_MUX4_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.5 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.485 2.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.48 2.25 0.755 ;
      RECT  2.15 0.755 2.33 0.925 ;
      RECT  2.15 0.925 2.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.525 3.45 0.755 ;
      RECT  3.22 0.755 3.45 0.925 ;
      RECT  3.35 0.925 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0636 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.145 0.14 4.38 0.23 ;
      RECT  4.145 0.23 4.25 0.35 ;
      RECT  4.07 0.35 4.25 0.45 ;
      LAYER M2 ;
      RECT  4.07 0.35 4.745 0.45 ;
      LAYER V1 ;
      RECT  4.11 0.35 4.21 0.45 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.835 1.475 1.015 1.75 ;
      RECT  2.06 1.44 2.19 1.75 ;
      RECT  3.28 1.495 3.455 1.75 ;
      RECT  4.525 1.44 4.655 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  2.045 0.05 2.185 0.385 ;
      RECT  4.525 0.05 4.655 0.385 ;
      RECT  0.075 0.05 0.205 0.39 ;
      RECT  0.86 0.05 0.99 0.39 ;
      RECT  3.305 0.05 3.435 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.31 4.91 0.495 ;
      RECT  4.75 0.495 4.85 1.11 ;
      RECT  4.75 1.11 4.895 1.295 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.465 0.235 3.085 0.335 ;
      RECT  2.985 0.335 3.085 0.925 ;
      RECT  2.465 0.335 2.565 0.955 ;
      RECT  1.14 0.285 1.52 0.415 ;
      RECT  1.14 0.415 1.36 0.495 ;
      RECT  3.7 0.35 3.945 0.45 ;
      RECT  3.805 0.45 3.945 0.585 ;
      RECT  3.855 0.585 3.945 1.28 ;
      RECT  3.755 1.28 3.945 1.45 ;
      RECT  4.345 0.48 4.455 0.585 ;
      RECT  4.345 0.585 4.66 0.69 ;
      RECT  4.57 0.69 4.66 1.24 ;
      RECT  4.31 1.24 4.66 1.34 ;
      RECT  4.31 1.34 4.41 1.565 ;
      RECT  2.95 1.295 3.655 1.395 ;
      RECT  2.95 1.395 3.05 1.44 ;
      RECT  3.56 1.395 3.655 1.565 ;
      RECT  2.55 1.44 3.05 1.56 ;
      RECT  3.56 1.565 4.41 1.66 ;
      RECT  4.04 0.54 4.21 0.63 ;
      RECT  4.04 0.63 4.145 0.89 ;
      RECT  4.04 0.89 4.46 1.06 ;
      RECT  4.04 1.06 4.15 1.47 ;
      RECT  3.54 0.55 3.715 0.65 ;
      RECT  3.585 0.65 3.675 0.76 ;
      RECT  3.585 0.76 3.75 0.93 ;
      RECT  3.585 0.93 3.675 1.19 ;
      RECT  2.695 0.43 2.895 0.69 ;
      RECT  1.465 0.51 1.635 0.94 ;
      RECT  1.725 0.725 1.825 1.17 ;
      RECT  1.725 1.17 1.885 1.26 ;
      RECT  1.795 1.26 2.79 1.35 ;
      RECT  2.7 0.79 2.79 1.26 ;
      RECT  1.795 1.35 1.885 1.55 ;
      RECT  0.355 0.37 0.485 0.59 ;
      RECT  0.395 0.59 0.485 0.73 ;
      RECT  0.395 0.73 0.53 0.95 ;
      RECT  0.395 0.95 0.485 1.17 ;
      RECT  0.355 1.17 0.485 1.295 ;
      RECT  0.355 1.295 1.335 1.385 ;
      RECT  1.24 0.63 1.335 1.295 ;
      RECT  1.24 1.385 1.335 1.55 ;
      RECT  1.24 1.55 1.885 1.64 ;
      RECT  0.62 0.31 0.72 1.19 ;
      RECT  1.455 1.05 1.56 1.35 ;
      RECT  1.455 1.35 1.705 1.45 ;
      LAYER M2 ;
      RECT  1.22 0.35 3.9 0.45 ;
      RECT  0.58 0.55 2.605 0.65 ;
      RECT  2.74 0.55 4.495 0.65 ;
      RECT  1.455 1.35 3.935 1.45 ;
      LAYER V1 ;
      RECT  1.26 0.35 1.36 0.45 ;
      RECT  3.76 0.35 3.86 0.45 ;
      RECT  0.62 0.55 0.72 0.65 ;
      RECT  1.465 0.55 1.565 0.65 ;
      RECT  2.465 0.55 2.565 0.65 ;
      RECT  2.78 0.55 2.88 0.65 ;
      RECT  4.355 0.55 4.455 0.65 ;
      RECT  1.565 1.35 1.665 1.45 ;
      RECT  3.795 1.35 3.895 1.45 ;
  END
END SEN_MUX4_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX4_D_2
#      Description : "4-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX4_D_2
  CLASS CORE ;
  FOREIGN SEN_MUX4_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.5 1.25 0.7 ;
      RECT  1.15 0.7 1.65 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.525 0.51 3.85 0.69 ;
      RECT  3.695 0.69 3.85 0.8 ;
      RECT  3.695 0.8 4.055 0.97 ;
      LAYER M2 ;
      RECT  3.3 0.55 4.1 0.65 ;
      LAYER V1 ;
      RECT  3.525 0.55 3.625 0.65 ;
      RECT  3.725 0.55 3.825 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.65 0.69 ;
      RECT  4.35 0.69 4.45 0.9 ;
      LAYER M2 ;
      RECT  4.31 0.55 5.1 0.65 ;
      LAYER V1 ;
      RECT  4.35 0.55 4.45 0.65 ;
      RECT  4.55 0.55 4.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.48 0.71 7.05 0.89 ;
      RECT  6.95 0.89 7.05 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1272 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.49 0.25 1.32 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.7 7.85 0.925 ;
      RECT  7.55 0.925 7.85 1.1 ;
      RECT  7.55 1.1 7.65 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1896 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.585 1.215 0.705 1.75 ;
      RECT  1.12 1.215 1.225 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  3.56 1.41 3.675 1.75 ;
      RECT  4.065 1.21 4.185 1.75 ;
      RECT  4.585 1.21 4.705 1.75 ;
      RECT  6.385 1.21 6.505 1.75 ;
      RECT  6.9 1.41 7.03 1.75 ;
      RECT  7.42 1.41 7.55 1.75 ;
      RECT  8.91 0.97 9.015 1.75 ;
      RECT  9.415 1.41 9.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  3.47 0.05 3.64 0.195 ;
      RECT  4.36 0.05 4.53 0.21 ;
      RECT  6.51 0.05 6.64 0.36 ;
      RECT  1.1 0.05 1.23 0.38 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  9.42 0.05 9.545 0.39 ;
      RECT  1.62 0.05 1.75 0.41 ;
      RECT  7.28 0.05 7.41 0.41 ;
      RECT  0.585 0.05 0.705 0.59 ;
      RECT  8.905 0.05 9.025 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.15 0.5 9.285 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.875 0.16 2.515 0.25 ;
      RECT  1.875 0.25 1.995 0.41 ;
      RECT  2.395 0.25 2.515 0.465 ;
      RECT  2.395 0.465 3.33 0.555 ;
      RECT  2.91 0.345 3.035 0.465 ;
      RECT  3.24 0.555 3.33 1.0 ;
      RECT  3.175 1.0 3.33 1.09 ;
      RECT  3.175 1.09 3.29 1.21 ;
      RECT  2.655 1.21 3.29 1.3 ;
      RECT  3.11 1.3 3.29 1.45 ;
      RECT  2.655 1.3 2.775 1.46 ;
      RECT  2.11 1.46 2.775 1.575 ;
      RECT  2.655 0.16 3.295 0.25 ;
      RECT  3.175 0.25 3.295 0.285 ;
      RECT  2.655 0.25 2.775 0.375 ;
      RECT  3.175 0.285 3.935 0.375 ;
      RECT  3.815 0.19 3.935 0.285 ;
      RECT  5.735 0.16 6.365 0.25 ;
      RECT  5.735 0.25 5.855 0.36 ;
      RECT  6.265 0.25 6.365 0.45 ;
      RECT  6.265 0.45 6.92 0.55 ;
      RECT  4.065 0.19 4.185 0.3 ;
      RECT  4.065 0.3 5.37 0.4 ;
      RECT  7.545 0.25 8.045 0.34 ;
      RECT  7.545 0.34 7.66 0.5 ;
      RECT  7.03 0.37 7.145 0.5 ;
      RECT  7.03 0.5 7.66 0.59 ;
      RECT  7.14 0.59 7.23 1.14 ;
      RECT  7.14 1.14 7.28 1.34 ;
      RECT  0.32 0.215 0.46 0.39 ;
      RECT  0.37 0.39 0.46 0.945 ;
      RECT  0.37 0.945 0.85 1.01 ;
      RECT  0.75 0.715 0.85 0.945 ;
      RECT  0.34 1.01 0.85 1.05 ;
      RECT  0.75 1.05 0.85 1.09 ;
      RECT  0.34 1.05 0.485 1.31 ;
      RECT  5.48 0.29 5.59 0.47 ;
      RECT  5.48 0.47 6.115 0.53 ;
      RECT  5.99 0.355 6.115 0.47 ;
      RECT  4.91 0.53 6.115 0.56 ;
      RECT  4.91 0.56 5.725 0.65 ;
      RECT  5.625 0.65 5.725 1.55 ;
      RECT  5.095 1.415 5.215 1.55 ;
      RECT  5.095 1.55 6.255 1.64 ;
      RECT  6.135 1.37 6.255 1.55 ;
      RECT  1.365 0.37 1.485 0.5 ;
      RECT  1.365 0.5 2.255 0.59 ;
      RECT  2.135 0.34 2.255 0.5 ;
      RECT  7.8 0.43 8.455 0.52 ;
      RECT  7.8 0.52 7.91 0.61 ;
      RECT  8.31 0.52 8.455 0.65 ;
      RECT  8.31 0.65 8.4 0.87 ;
      RECT  8.25 0.87 8.4 0.96 ;
      RECT  8.25 0.96 8.34 1.37 ;
      RECT  8.2 1.37 8.34 1.54 ;
      RECT  7.675 1.41 7.8 1.54 ;
      RECT  7.675 1.54 8.82 1.63 ;
      RECT  8.73 0.775 8.82 1.54 ;
      RECT  8.55 0.545 8.74 0.655 ;
      RECT  8.55 0.655 8.64 1.305 ;
      RECT  8.43 1.305 8.64 1.41 ;
      RECT  2.4 0.645 3.15 0.735 ;
      RECT  2.4 0.735 2.49 0.8 ;
      RECT  2.995 0.735 3.15 0.91 ;
      RECT  1.875 0.8 2.49 0.89 ;
      RECT  1.875 0.89 2.0 1.01 ;
      RECT  0.82 0.48 1.03 0.59 ;
      RECT  0.94 0.59 1.03 1.01 ;
      RECT  0.94 1.01 2.0 1.1 ;
      RECT  0.94 1.1 1.03 1.19 ;
      RECT  0.795 1.19 1.03 1.3 ;
      RECT  8.0 0.61 8.18 0.805 ;
      RECT  8.0 0.805 8.09 1.215 ;
      RECT  7.91 1.215 8.09 1.45 ;
      RECT  4.775 0.75 5.165 0.85 ;
      RECT  5.02 0.85 5.165 1.11 ;
      RECT  5.86 0.65 6.075 0.89 ;
      RECT  4.325 1.01 4.93 1.1 ;
      RECT  4.835 1.1 4.93 1.21 ;
      RECT  4.325 1.1 4.44 1.385 ;
      RECT  4.835 1.21 5.475 1.3 ;
      RECT  5.355 1.3 5.475 1.43 ;
      RECT  4.835 1.3 4.955 1.6 ;
      RECT  2.715 0.85 2.905 1.12 ;
      RECT  5.255 0.74 5.465 1.12 ;
      RECT  5.875 1.03 6.765 1.12 ;
      RECT  6.645 1.12 6.765 1.25 ;
      RECT  5.875 1.12 6.0 1.42 ;
      RECT  1.34 1.2 2.54 1.3 ;
      RECT  1.34 1.3 1.51 1.325 ;
      RECT  1.875 1.3 2.0 1.57 ;
      RECT  3.38 1.21 3.86 1.3 ;
      RECT  3.765 1.3 3.86 1.4 ;
      RECT  3.38 1.3 3.47 1.56 ;
      RECT  3.765 1.4 3.92 1.62 ;
      RECT  2.915 1.4 3.02 1.56 ;
      RECT  2.915 1.56 3.47 1.65 ;
      LAYER M2 ;
      RECT  5.37 0.55 8.73 0.65 ;
      RECT  2.94 0.75 6.12 0.85 ;
      RECT  0.51 0.95 5.445 1.05 ;
      RECT  3.11 1.35 8.09 1.45 ;
      LAYER V1 ;
      RECT  5.45 0.55 5.55 0.65 ;
      RECT  8.59 0.55 8.69 0.65 ;
      RECT  3.015 0.75 3.115 0.85 ;
      RECT  4.815 0.75 4.915 0.85 ;
      RECT  5.025 0.75 5.125 0.85 ;
      RECT  5.915 0.75 6.015 0.85 ;
      RECT  0.55 0.95 0.65 1.05 ;
      RECT  0.75 0.95 0.85 1.05 ;
      RECT  2.775 0.95 2.875 1.05 ;
      RECT  5.275 0.95 5.375 1.05 ;
      RECT  3.15 1.35 3.25 1.45 ;
      RECT  7.95 1.35 8.05 1.45 ;
  END
END SEN_MUX4_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUX4_D_4
#      Description : "4-1 multiplexer"
#      Equation    : X=((D0&!S0&!S1)|(D1&S0&!S1)|(D2&!S0&S1)|(D3&S0&S1))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUX4_D_4
  CLASS CORE ;
  FOREIGN SEN_MUX4_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 16.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.5 2.25 0.7 ;
      RECT  2.15 0.7 2.85 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.415 0.755 7.185 0.9 ;
      RECT  7.085 0.9 7.185 1.3 ;
      LAYER M2 ;
      RECT  6.835 1.15 7.435 1.25 ;
      LAYER V1 ;
      RECT  7.085 1.15 7.185 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 ;
  END D1
  PIN D2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.42 0.51 7.785 0.69 ;
      RECT  7.485 0.69 7.785 0.9 ;
      LAYER M2 ;
      RECT  7.38 0.55 7.97 0.65 ;
      LAYER V1 ;
      RECT  7.42 0.55 7.52 0.65 ;
      RECT  7.62 0.55 7.72 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 ;
  END D2
  PIN D3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.22 0.71 12.05 0.89 ;
      RECT  11.95 0.89 12.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2544 ;
  END D3
  PIN S0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.7 0.9 ;
      RECT  0.15 0.9 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END S0
  PIN S1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.55 0.7 13.25 0.9 ;
      RECT  13.15 0.9 13.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3792 ;
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 16.2 1.85 ;
      RECT  0.585 1.21 0.705 1.75 ;
      RECT  1.105 1.21 1.225 1.75 ;
      RECT  1.625 1.215 1.745 1.75 ;
      RECT  2.145 1.21 2.265 1.75 ;
      RECT  2.66 1.435 2.79 1.75 ;
      RECT  3.18 1.41 3.31 1.75 ;
      RECT  5.97 1.41 6.1 1.75 ;
      RECT  6.49 1.41 6.62 1.75 ;
      RECT  7.01 1.41 7.14 1.75 ;
      RECT  7.535 1.21 7.655 1.75 ;
      RECT  8.05 1.41 8.18 1.75 ;
      RECT  10.825 1.415 10.955 1.75 ;
      RECT  11.345 1.415 11.475 1.75 ;
      RECT  11.91 1.21 12.03 1.75 ;
      RECT  12.46 1.21 12.58 1.75 ;
      RECT  12.975 1.17 13.085 1.75 ;
      RECT  14.975 1.44 15.105 1.75 ;
      RECT  15.495 1.41 15.625 1.75 ;
      RECT  16.015 1.41 16.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 16.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
      RECT  14.65 1.75 14.75 1.85 ;
      RECT  15.25 1.75 15.35 1.85 ;
      RECT  15.85 1.75 15.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 16.2 0.05 ;
      RECT  7.555 0.05 7.725 0.21 ;
      RECT  6.29 0.05 6.42 0.38 ;
      RECT  6.81 0.05 6.94 0.38 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.62 0.05 1.75 0.385 ;
      RECT  8.155 0.05 8.285 0.385 ;
      RECT  2.14 0.05 2.27 0.39 ;
      RECT  2.66 0.05 2.79 0.39 ;
      RECT  3.18 0.05 3.31 0.39 ;
      RECT  12.49 0.05 12.62 0.39 ;
      RECT  13.01 0.05 13.14 0.39 ;
      RECT  15.495 0.05 15.625 0.39 ;
      RECT  16.015 0.05 16.14 0.39 ;
      RECT  11.265 0.05 11.395 0.41 ;
      RECT  11.785 0.05 11.915 0.41 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.105 0.05 1.225 0.59 ;
      RECT  14.98 0.05 15.1 0.68 ;
      LAYER M2 ;
      RECT  0.0 -0.05 16.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
      RECT  14.65 -0.05 14.75 0.05 ;
      RECT  15.25 -0.05 15.35 0.05 ;
      RECT  15.85 -0.05 15.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  15.215 0.51 15.875 0.69 ;
      RECT  15.75 0.69 15.875 1.11 ;
      RECT  15.24 1.11 15.875 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.63 0.16 4.795 0.25 ;
      RECT  3.63 0.25 3.75 0.385 ;
      RECT  4.15 0.25 4.27 0.385 ;
      RECT  4.665 0.25 4.795 0.435 ;
      RECT  4.665 0.435 5.92 0.545 ;
      RECT  5.82 0.545 5.92 0.98 ;
      RECT  5.34 0.98 5.92 1.07 ;
      RECT  5.34 1.07 5.43 1.21 ;
      RECT  4.67 1.21 5.43 1.3 ;
      RECT  5.18 1.3 5.36 1.45 ;
      RECT  4.67 1.3 4.79 1.485 ;
      RECT  3.635 1.41 3.745 1.485 ;
      RECT  3.635 1.485 4.79 1.595 ;
      RECT  13.725 0.16 14.89 0.25 ;
      RECT  14.755 0.25 14.89 0.39 ;
      RECT  13.725 0.25 13.83 0.6 ;
      RECT  14.23 0.25 14.345 0.95 ;
      RECT  13.975 0.95 14.955 1.04 ;
      RECT  14.835 1.04 14.955 1.12 ;
      RECT  13.975 1.04 14.09 1.54 ;
      RECT  13.445 1.425 13.565 1.54 ;
      RECT  13.445 1.54 14.605 1.63 ;
      RECT  14.49 1.425 14.605 1.54 ;
      RECT  9.92 0.2 11.13 0.31 ;
      RECT  11.01 0.31 11.13 0.5 ;
      RECT  11.01 0.5 12.16 0.59 ;
      RECT  12.055 0.17 12.16 0.5 ;
      RECT  4.94 0.2 6.155 0.315 ;
      RECT  6.035 0.315 6.155 0.49 ;
      RECT  6.035 0.49 7.22 0.6 ;
      RECT  7.05 0.6 7.22 0.64 ;
      RECT  8.42 0.225 9.63 0.325 ;
      RECT  8.42 0.325 8.54 0.5 ;
      RECT  7.26 0.17 7.38 0.3 ;
      RECT  7.26 0.3 8.02 0.39 ;
      RECT  7.9 0.39 8.02 0.5 ;
      RECT  7.9 0.5 8.54 0.59 ;
      RECT  13.25 0.23 13.635 0.345 ;
      RECT  13.25 0.345 13.34 0.49 ;
      RECT  12.25 0.49 13.34 0.59 ;
      RECT  12.25 0.59 12.455 0.68 ;
      RECT  12.355 0.68 12.455 1.01 ;
      RECT  12.21 1.01 12.835 1.1 ;
      RECT  12.21 1.1 12.315 1.26 ;
      RECT  12.725 1.1 12.835 1.26 ;
      RECT  2.4 0.37 2.525 0.485 ;
      RECT  2.4 0.485 4.01 0.5 ;
      RECT  3.89 0.375 4.01 0.485 ;
      RECT  2.4 0.5 4.535 0.59 ;
      RECT  4.41 0.375 4.535 0.5 ;
      RECT  9.685 0.455 10.92 0.485 ;
      RECT  8.655 0.485 10.92 0.56 ;
      RECT  8.655 0.56 9.91 0.59 ;
      RECT  9.545 0.59 9.91 0.655 ;
      RECT  9.545 0.655 9.655 1.55 ;
      RECT  8.5 1.415 8.62 1.55 ;
      RECT  8.5 1.55 10.7 1.64 ;
      RECT  9.02 1.415 9.14 1.55 ;
      RECT  10.06 1.415 10.18 1.55 ;
      RECT  10.58 1.415 10.7 1.55 ;
      RECT  0.3 0.485 0.99 0.595 ;
      RECT  0.89 0.595 0.99 0.71 ;
      RECT  0.89 0.71 1.85 0.89 ;
      RECT  0.89 0.89 1.2 1.015 ;
      RECT  0.34 1.015 1.2 1.095 ;
      RECT  0.34 1.095 0.965 1.105 ;
      RECT  0.34 1.105 0.445 1.27 ;
      RECT  0.845 1.105 0.965 1.27 ;
      RECT  5.345 0.645 5.715 0.665 ;
      RECT  4.645 0.665 5.715 0.755 ;
      RECT  4.645 0.755 4.735 0.8 ;
      RECT  5.345 0.755 5.715 0.89 ;
      RECT  3.0 0.8 4.735 0.89 ;
      RECT  3.0 0.89 3.09 1.01 ;
      RECT  1.34 0.49 2.03 0.59 ;
      RECT  1.94 0.59 2.03 1.01 ;
      RECT  1.375 1.01 3.09 1.1 ;
      RECT  1.375 1.1 1.48 1.28 ;
      RECT  1.885 1.1 2.01 1.28 ;
      RECT  13.465 0.54 13.575 0.715 ;
      RECT  13.465 0.715 14.1 0.805 ;
      RECT  13.98 0.5 14.1 0.715 ;
      RECT  13.79 0.805 13.88 1.215 ;
      RECT  13.185 1.215 13.88 1.315 ;
      RECT  13.185 1.315 13.285 1.63 ;
      RECT  10.205 0.65 10.74 0.75 ;
      RECT  10.205 0.75 10.575 0.89 ;
      RECT  14.49 0.4 14.615 0.77 ;
      RECT  14.49 0.77 15.15 0.86 ;
      RECT  15.05 0.86 15.15 1.225 ;
      RECT  14.2 1.225 15.15 1.325 ;
      RECT  14.2 1.325 14.72 1.33 ;
      RECT  9.06 0.73 9.45 0.84 ;
      RECT  9.06 0.84 9.36 1.09 ;
      RECT  8.275 0.75 8.665 0.85 ;
      RECT  8.475 0.85 8.665 0.93 ;
      RECT  8.475 0.93 8.845 1.045 ;
      RECT  8.475 1.045 8.665 1.05 ;
      RECT  4.845 0.85 5.215 1.09 ;
      RECT  3.385 1.01 4.53 1.1 ;
      RECT  3.385 1.1 3.48 1.205 ;
      RECT  4.41 1.1 4.53 1.39 ;
      RECT  3.89 1.1 4.01 1.395 ;
      RECT  2.38 1.205 3.48 1.305 ;
      RECT  7.275 1.01 8.36 1.1 ;
      RECT  8.245 1.1 8.36 1.195 ;
      RECT  7.275 1.1 7.395 1.24 ;
      RECT  7.8 1.1 7.915 1.27 ;
      RECT  8.245 1.195 9.455 1.3 ;
      RECT  5.52 1.16 6.905 1.25 ;
      RECT  5.52 1.25 5.61 1.4 ;
      RECT  5.45 1.4 5.61 1.56 ;
      RECT  4.945 1.4 5.065 1.56 ;
      RECT  4.945 1.56 5.61 1.65 ;
      RECT  9.745 1.2 11.78 1.315 ;
      RECT  5.7 1.35 5.88 1.65 ;
      LAYER M2 ;
      RECT  9.43 0.55 14.74 0.65 ;
      RECT  5.305 0.75 10.56 0.85 ;
      RECT  0.85 0.95 9.4 1.05 ;
      RECT  5.08 1.35 13.325 1.45 ;
      LAYER V1 ;
      RECT  9.55 0.55 9.65 0.65 ;
      RECT  9.77 0.55 9.87 0.65 ;
      RECT  14.49 0.55 14.59 0.65 ;
      RECT  5.345 0.75 5.445 0.85 ;
      RECT  5.555 0.75 5.655 0.85 ;
      RECT  8.315 0.75 8.415 0.85 ;
      RECT  8.525 0.75 8.625 0.85 ;
      RECT  10.22 0.75 10.32 0.85 ;
      RECT  10.42 0.75 10.52 0.85 ;
      RECT  0.89 0.95 0.99 1.05 ;
      RECT  1.1 0.95 1.2 1.05 ;
      RECT  4.885 0.95 4.985 1.05 ;
      RECT  5.085 0.95 5.185 1.05 ;
      RECT  9.06 0.95 9.16 1.05 ;
      RECT  9.26 0.95 9.36 1.05 ;
      RECT  5.22 1.35 5.32 1.45 ;
      RECT  5.74 1.35 5.84 1.45 ;
      RECT  13.185 1.35 13.285 1.45 ;
  END
END SEN_MUX4_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_0P75
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_0P75
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.32 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.14 1.65 0.23 ;
      RECT  0.55 0.23 0.65 0.51 ;
      RECT  1.55 0.23 1.65 0.71 ;
      RECT  0.35 0.51 0.65 0.6 ;
      RECT  0.35 0.6 0.45 0.795 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  0.26 0.795 0.45 0.975 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0759 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.445 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.81 1.21 1.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  1.81 0.05 1.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.07 0.32 1.25 0.5 ;
      RECT  1.15 0.5 1.25 1.055 ;
      RECT  1.045 1.055 1.25 1.145 ;
    END
    ANTENNADIFFAREA 0.192 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.8 1.125 0.925 1.24 ;
      RECT  0.8 1.24 1.72 1.33 ;
      RECT  0.065 0.195 0.17 1.26 ;
      RECT  0.065 1.26 0.645 1.35 ;
      RECT  0.555 0.74 0.645 1.26 ;
      RECT  0.065 1.35 0.185 1.635 ;
      RECT  0.55 1.445 1.51 1.56 ;
  END
END SEN_MUXI2_DG_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_1
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_1
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.32 0.85 0.71 ;
      RECT  0.75 0.71 1.05 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.14 1.65 0.23 ;
      RECT  0.55 0.23 0.65 0.51 ;
      RECT  1.55 0.23 1.65 0.71 ;
      RECT  0.35 0.51 0.65 0.6 ;
      RECT  0.35 0.6 0.45 0.725 ;
      RECT  1.55 0.71 1.85 0.91 ;
      RECT  0.26 0.725 0.45 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0927 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.445 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.81 1.21 1.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  1.81 0.05 1.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.07 0.32 1.25 0.5 ;
      RECT  1.15 0.5 1.25 1.055 ;
      RECT  1.02 1.055 1.25 1.145 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.195 0.17 1.26 ;
      RECT  0.065 1.26 0.645 1.35 ;
      RECT  0.555 0.72 0.645 1.26 ;
      RECT  0.065 1.35 0.185 1.635 ;
      RECT  0.76 1.24 1.72 1.33 ;
      RECT  0.535 1.445 1.5 1.56 ;
  END
END SEN_MUXI2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_10
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_10
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.45 0.745 ;
      RECT  3.35 0.745 6.09 0.85 ;
      RECT  4.45 0.71 6.09 0.745 ;
      RECT  4.41 0.85 6.09 0.89 ;
      RECT  3.35 0.85 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.73 0.71 8.25 0.74 ;
      RECT  6.73 0.74 9.45 0.84 ;
      RECT  9.35 0.71 9.45 0.74 ;
      RECT  6.73 0.84 8.25 0.89 ;
      RECT  9.35 0.84 9.45 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.75 0.51 11.85 0.71 ;
      RECT  9.75 0.71 11.85 0.89 ;
      RECT  0.79 0.51 0.89 0.71 ;
      RECT  0.35 0.71 0.89 0.9 ;
      LAYER M2 ;
      RECT  0.75 0.55 11.89 0.65 ;
      LAYER V1 ;
      RECT  11.75 0.55 11.85 0.65 ;
      RECT  0.79 0.55 0.89 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.81 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.44 0.46 1.75 ;
      RECT  0.0 1.75 12.0 1.85 ;
      RECT  0.88 1.44 1.01 1.75 ;
      RECT  1.405 1.255 1.525 1.75 ;
      RECT  1.925 1.255 2.045 1.75 ;
      RECT  2.445 1.255 2.565 1.75 ;
      RECT  2.96 1.425 3.09 1.75 ;
      RECT  3.48 1.425 3.61 1.75 ;
      RECT  9.19 1.495 9.36 1.75 ;
      RECT  9.71 1.495 9.88 1.75 ;
      RECT  10.25 1.455 10.38 1.75 ;
      RECT  10.77 1.455 10.9 1.75 ;
      RECT  11.29 1.455 11.42 1.75 ;
      RECT  11.815 1.21 11.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.0 0.05 ;
      RECT  1.38 0.05 1.55 0.305 ;
      RECT  1.9 0.05 2.07 0.305 ;
      RECT  2.42 0.05 2.59 0.305 ;
      RECT  2.94 0.05 3.11 0.305 ;
      RECT  9.71 0.05 9.88 0.305 ;
      RECT  10.23 0.05 10.4 0.305 ;
      RECT  10.75 0.05 10.92 0.305 ;
      RECT  11.27 0.05 11.44 0.305 ;
      RECT  3.46 0.05 3.63 0.32 ;
      RECT  9.19 0.05 9.36 0.32 ;
      RECT  0.33 0.05 0.46 0.36 ;
      RECT  11.81 0.05 11.94 0.39 ;
      RECT  0.88 0.05 1.01 0.42 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.72 0.17 9.09 0.26 ;
      RECT  4.76 0.26 9.09 0.3 ;
      RECT  4.24 0.26 4.41 0.305 ;
      RECT  3.72 0.26 3.89 0.32 ;
      RECT  4.76 0.3 8.57 0.32 ;
      RECT  8.92 0.3 9.09 0.32 ;
      RECT  5.28 0.32 8.05 0.345 ;
      RECT  6.3 0.345 6.51 0.98 ;
      RECT  3.695 0.98 9.09 1.02 ;
      RECT  8.395 0.93 9.09 0.98 ;
      RECT  8.92 1.02 9.09 1.105 ;
      RECT  3.695 1.02 8.53 1.12 ;
      RECT  4.77 1.12 8.53 1.155 ;
    END
    ANTENNADIFFAREA 2.274 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.12 0.41 4.675 0.445 ;
      RECT  1.12 0.445 6.19 0.575 ;
      RECT  2.68 0.575 6.19 0.62 ;
      RECT  3.505 0.62 4.4 0.63 ;
      RECT  8.655 0.41 11.66 0.45 ;
      RECT  6.62 0.45 11.66 0.58 ;
      RECT  6.62 0.58 9.62 0.62 ;
      RECT  0.98 0.79 2.795 0.89 ;
      RECT  0.98 0.89 1.07 1.23 ;
      RECT  0.595 0.35 0.7 0.455 ;
      RECT  0.05 0.455 0.7 0.575 ;
      RECT  0.05 0.575 0.14 1.23 ;
      RECT  0.05 1.23 1.07 1.35 ;
      RECT  1.16 0.995 3.26 1.165 ;
      RECT  3.05 1.165 3.26 1.215 ;
      RECT  3.05 1.215 3.61 1.245 ;
      RECT  3.05 1.245 8.79 1.335 ;
      RECT  8.69 1.11 8.79 1.245 ;
      RECT  8.89 1.195 11.675 1.365 ;
      RECT  8.89 1.365 10.135 1.405 ;
      RECT  8.89 1.405 9.1 1.445 ;
      RECT  3.98 1.445 9.1 1.62 ;
      RECT  6.085 1.62 9.1 1.64 ;
      LAYER M2 ;
      RECT  3.08 1.15 8.86 1.25 ;
      LAYER V1 ;
      RECT  3.15 1.15 3.25 1.25 ;
      RECT  8.69 1.15 8.79 1.25 ;
  END
END SEN_MUXI2_DG_10
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_12
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_12
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.71 6.25 0.79 ;
      RECT  3.95 0.79 6.25 0.88 ;
      RECT  5.015 0.88 6.25 0.89 ;
      RECT  3.95 0.88 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.75 0.71 9.05 0.79 ;
      RECT  8.75 0.79 11.05 0.88 ;
      RECT  8.75 0.88 9.945 0.89 ;
      RECT  10.95 0.88 11.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  13.88 0.51 13.98 0.71 ;
      RECT  11.78 0.71 13.98 0.89 ;
      RECT  0.79 0.51 0.89 0.71 ;
      RECT  0.35 0.71 0.89 0.89 ;
      LAYER M2 ;
      RECT  0.75 0.55 14.02 0.65 ;
      LAYER V1 ;
      RECT  13.88 0.55 13.98 0.65 ;
      RECT  0.79 0.55 0.89 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.972 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.415 0.46 1.75 ;
      RECT  0.0 1.75 14.2 1.85 ;
      RECT  0.88 1.415 1.01 1.75 ;
      RECT  1.405 1.255 1.525 1.75 ;
      RECT  1.925 1.255 2.045 1.75 ;
      RECT  2.445 1.255 2.565 1.75 ;
      RECT  2.94 1.48 3.11 1.75 ;
      RECT  3.46 1.48 3.63 1.75 ;
      RECT  3.98 1.48 4.15 1.75 ;
      RECT  10.81 1.44 10.92 1.75 ;
      RECT  11.31 1.455 11.44 1.75 ;
      RECT  11.83 1.455 11.96 1.75 ;
      RECT  12.35 1.455 12.48 1.75 ;
      RECT  12.87 1.455 13.0 1.75 ;
      RECT  13.39 1.455 13.52 1.75 ;
      RECT  13.935 1.21 14.055 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 14.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
      RECT  11.85 1.75 11.95 1.85 ;
      RECT  12.45 1.75 12.55 1.85 ;
      RECT  13.05 1.75 13.15 1.85 ;
      RECT  13.65 1.75 13.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 14.2 0.05 ;
      RECT  3.46 0.05 3.63 0.32 ;
      RECT  3.98 0.05 4.15 0.32 ;
      RECT  10.77 0.05 10.94 0.32 ;
      RECT  11.29 0.05 11.46 0.32 ;
      RECT  11.81 0.05 11.98 0.32 ;
      RECT  0.34 0.05 0.46 0.36 ;
      RECT  12.35 0.05 12.48 0.36 ;
      RECT  12.87 0.05 13.0 0.36 ;
      RECT  13.39 0.05 13.52 0.36 ;
      RECT  0.88 0.05 1.01 0.385 ;
      RECT  1.4 0.05 1.53 0.385 ;
      RECT  1.92 0.05 2.05 0.385 ;
      RECT  2.44 0.05 2.57 0.385 ;
      RECT  2.955 0.05 3.09 0.385 ;
      RECT  13.93 0.05 14.06 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 14.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
      RECT  11.85 -0.05 11.95 0.05 ;
      RECT  12.45 -0.05 12.55 0.05 ;
      RECT  13.05 -0.05 13.15 0.05 ;
      RECT  13.65 -0.05 13.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.255 0.17 10.665 0.32 ;
      RECT  5.295 0.32 9.625 0.34 ;
      RECT  6.895 0.34 9.625 0.345 ;
      RECT  6.895 0.345 8.03 0.38 ;
      RECT  7.35 0.38 7.56 0.895 ;
      RECT  6.75 0.895 8.05 0.91 ;
      RECT  6.34 0.91 8.65 0.98 ;
      RECT  4.255 0.97 4.88 0.98 ;
      RECT  4.255 0.98 10.665 1.06 ;
      RECT  10.06 0.97 10.665 0.98 ;
      RECT  4.255 1.06 4.425 1.105 ;
      RECT  4.775 1.06 10.145 1.105 ;
      RECT  10.495 1.06 10.665 1.105 ;
    END
    ANTENNADIFFAREA 2.74 ;
  END X
  OBS
      LAYER M1 ;
      RECT  9.21 0.435 12.24 0.46 ;
      RECT  9.21 0.46 13.76 0.48 ;
      RECT  13.67 0.435 13.76 0.46 ;
      RECT  7.675 0.48 13.76 0.605 ;
      RECT  7.675 0.605 11.68 0.61 ;
      RECT  9.17 0.61 11.68 0.63 ;
      RECT  7.675 0.61 7.765 0.65 ;
      RECT  9.725 0.63 11.68 0.68 ;
      RECT  3.195 0.43 5.73 0.49 ;
      RECT  1.12 0.49 7.245 0.62 ;
      RECT  1.12 0.62 5.78 0.63 ;
      RECT  7.155 0.62 7.245 0.66 ;
      RECT  1.12 0.63 5.21 0.64 ;
      RECT  2.68 0.64 5.21 0.68 ;
      RECT  0.98 0.785 3.085 0.885 ;
      RECT  0.98 0.885 1.07 1.235 ;
      RECT  0.61 0.325 0.7 0.455 ;
      RECT  0.05 0.455 0.7 0.545 ;
      RECT  0.05 0.545 0.14 1.235 ;
      RECT  0.05 1.235 1.07 1.325 ;
      RECT  1.16 1.035 3.3 1.165 ;
      RECT  2.705 1.165 3.3 1.205 ;
      RECT  1.16 1.165 1.25 1.25 ;
      RECT  3.05 1.205 3.3 1.215 ;
      RECT  3.05 1.215 3.89 1.345 ;
      RECT  3.61 1.15 3.79 1.215 ;
      RECT  4.51 1.15 4.69 1.215 ;
      RECT  4.51 1.215 10.405 1.345 ;
      RECT  10.225 1.15 10.405 1.215 ;
      RECT  10.505 1.195 11.715 1.235 ;
      RECT  10.505 1.235 13.825 1.35 ;
      RECT  11.025 1.35 13.825 1.365 ;
      RECT  10.505 1.35 10.715 1.455 ;
      RECT  11.025 1.365 11.205 1.45 ;
      RECT  11.545 1.365 11.725 1.45 ;
      RECT  4.24 1.35 4.42 1.455 ;
      RECT  4.24 1.455 10.715 1.64 ;
      LAYER M2 ;
      RECT  3.11 1.15 10.405 1.25 ;
      RECT  4.24 1.35 11.745 1.45 ;
      LAYER V1 ;
      RECT  3.15 1.15 3.25 1.25 ;
      RECT  3.65 1.15 3.75 1.25 ;
      RECT  4.55 1.15 4.65 1.25 ;
      RECT  10.265 1.15 10.365 1.25 ;
      RECT  4.28 1.35 4.38 1.45 ;
      RECT  10.55 1.35 10.65 1.45 ;
      RECT  11.065 1.35 11.165 1.45 ;
      RECT  11.585 1.35 11.685 1.45 ;
  END
END SEN_MUXI2_DG_12
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_2
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_2
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.94 0.71 2.65 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.51 3.05 0.71 ;
      RECT  2.75 0.71 3.05 0.9 ;
      RECT  0.35 0.49 0.45 0.735 ;
      RECT  0.26 0.735 0.45 0.925 ;
      LAYER M2 ;
      RECT  0.31 0.55 3.09 0.65 ;
      LAYER V1 ;
      RECT  2.95 0.55 3.05 0.65 ;
      RECT  0.35 0.55 0.45 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.162 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.82 1.495 0.99 1.75 ;
      RECT  2.43 1.435 2.56 1.75 ;
      RECT  2.99 1.21 3.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.855 0.05 0.985 0.36 ;
      RECT  2.45 0.05 2.575 0.36 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  2.985 0.05 3.115 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.085 0.24 2.36 0.36 ;
      RECT  1.75 0.36 1.85 1.03 ;
      RECT  1.06 1.03 2.355 1.15 ;
    END
    ANTENNADIFFAREA 0.569 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.94 0.45 2.855 0.54 ;
      RECT  1.94 0.54 2.03 0.62 ;
      RECT  0.56 0.455 1.54 0.545 ;
      RECT  0.555 0.72 0.645 1.045 ;
      RECT  0.355 1.045 0.645 1.135 ;
      RECT  0.355 1.135 0.445 1.3 ;
      RECT  0.065 0.185 0.17 1.3 ;
      RECT  0.065 1.3 0.445 1.39 ;
      RECT  0.065 1.39 0.185 1.53 ;
      RECT  1.32 1.255 2.88 1.345 ;
      RECT  0.535 1.255 1.17 1.365 ;
      RECT  1.08 1.365 1.17 1.455 ;
      RECT  1.08 1.455 2.07 1.565 ;
  END
END SEN_MUXI2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_3
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_3
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.71 ;
      RECT  1.35 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.51 3.05 0.71 ;
      RECT  2.35 0.71 3.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.85 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
      RECT  0.15 0.71 0.25 1.13 ;
      LAYER M2 ;
      RECT  0.11 0.95 3.29 1.05 ;
      LAYER V1 ;
      RECT  3.15 0.95 3.25 1.05 ;
      RECT  0.15 0.95 0.25 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.845 1.235 0.965 1.75 ;
      RECT  3.435 1.45 3.565 1.75 ;
      RECT  3.98 1.21 4.1 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  0.84 0.05 0.97 0.36 ;
      RECT  3.44 0.05 3.565 0.385 ;
      RECT  3.98 0.05 4.1 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.565 0.45 2.825 0.56 ;
      RECT  2.15 0.56 2.25 1.04 ;
      RECT  1.565 1.04 2.825 1.16 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.345 0.215 3.35 0.335 ;
      RECT  3.26 0.335 3.35 0.475 ;
      RECT  3.26 0.475 3.87 0.595 ;
      RECT  1.08 0.24 2.045 0.36 ;
      RECT  1.08 0.36 1.17 0.45 ;
      RECT  0.54 0.45 1.17 0.56 ;
      RECT  0.065 0.245 0.185 0.45 ;
      RECT  0.065 0.45 0.45 0.54 ;
      RECT  0.36 0.54 0.45 0.79 ;
      RECT  0.36 0.79 1.02 0.89 ;
      RECT  0.36 0.89 0.45 1.26 ;
      RECT  0.065 1.26 0.45 1.35 ;
      RECT  0.065 1.35 0.185 1.525 ;
      RECT  0.54 1.055 1.225 1.145 ;
      RECT  1.105 1.145 1.225 1.45 ;
      RECT  1.105 1.45 3.085 1.56 ;
      RECT  1.315 1.25 3.87 1.36 ;
  END
END SEN_MUXI2_DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_4
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_4
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 2.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.985 0.51 5.085 0.71 ;
      RECT  4.35 0.71 5.085 0.89 ;
      RECT  0.23 0.51 0.33 0.93 ;
      LAYER M2 ;
      RECT  0.19 0.55 5.125 0.65 ;
      LAYER V1 ;
      RECT  4.985 0.55 5.085 0.65 ;
      RECT  0.23 0.55 0.33 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.44 0.45 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.845 1.21 0.965 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  3.965 1.44 4.095 1.75 ;
      RECT  4.485 1.45 4.615 1.75 ;
      RECT  5.01 1.21 5.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  0.84 0.05 0.97 0.36 ;
      RECT  1.36 0.05 1.485 0.36 ;
      RECT  3.97 0.05 4.095 0.36 ;
      RECT  4.485 0.05 4.615 0.36 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  5.005 0.05 5.135 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.575 0.25 3.875 0.36 ;
      RECT  2.75 0.36 2.85 1.04 ;
      RECT  1.575 1.04 3.85 1.16 ;
    END
    ANTENNADIFFAREA 0.994 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.56 0.45 2.575 0.56 ;
      RECT  2.94 0.455 4.895 0.56 ;
      RECT  2.94 0.56 3.045 0.65 ;
      RECT  0.42 0.79 1.135 0.89 ;
      RECT  0.42 0.89 0.51 1.26 ;
      RECT  0.05 0.225 0.185 0.42 ;
      RECT  0.05 0.42 0.14 1.26 ;
      RECT  0.05 1.26 0.51 1.35 ;
      RECT  0.05 1.35 0.185 1.525 ;
      RECT  0.6 1.03 1.225 1.12 ;
      RECT  0.6 1.12 0.69 1.25 ;
      RECT  1.105 1.12 1.225 1.25 ;
      RECT  1.105 1.25 3.615 1.35 ;
      RECT  3.75 1.25 4.92 1.35 ;
      RECT  3.75 1.35 3.84 1.45 ;
      RECT  1.835 1.45 3.84 1.56 ;
  END
END SEN_MUXI2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_5
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_5
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  2.15 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 4.85 0.71 ;
      RECT  3.75 0.71 4.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.26 0.71 5.96 0.89 ;
      RECT  5.26 0.89 5.36 1.09 ;
      RECT  0.15 0.71 0.51 0.89 ;
      RECT  0.41 0.89 0.51 1.13 ;
      LAYER M2 ;
      RECT  0.37 0.95 5.4 1.05 ;
      LAYER V1 ;
      RECT  5.26 0.95 5.36 1.05 ;
      RECT  0.41 0.95 0.51 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.405 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.215 0.185 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  1.105 1.235 1.225 1.75 ;
      RECT  1.625 1.255 1.745 1.75 ;
      RECT  5.155 1.455 5.275 1.75 ;
      RECT  5.675 1.45 5.795 1.75 ;
      RECT  6.215 1.215 6.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  0.065 0.05 0.185 0.36 ;
      RECT  0.585 0.05 0.705 0.36 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  1.625 0.05 1.745 0.36 ;
      RECT  5.155 0.05 5.275 0.36 ;
      RECT  5.675 0.05 5.795 0.36 ;
      RECT  6.215 0.05 6.335 0.56 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.365 0.45 4.575 0.56 ;
      RECT  2.365 0.56 2.455 0.62 ;
      RECT  3.34 0.56 3.45 1.04 ;
      RECT  2.325 1.04 4.575 1.16 ;
    END
    ANTENNADIFFAREA 1.08 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.625 0.215 5.065 0.335 ;
      RECT  4.975 0.335 5.065 0.475 ;
      RECT  4.975 0.475 6.085 0.595 ;
      RECT  1.86 0.24 3.275 0.36 ;
      RECT  1.86 0.36 1.95 0.45 ;
      RECT  0.82 0.45 1.95 0.56 ;
      RECT  0.325 0.27 0.445 0.45 ;
      RECT  0.325 0.45 0.71 0.54 ;
      RECT  0.62 0.54 0.71 0.79 ;
      RECT  0.62 0.79 1.55 0.89 ;
      RECT  0.62 0.89 0.71 1.26 ;
      RECT  0.325 1.26 0.71 1.35 ;
      RECT  0.325 1.35 0.445 1.5 ;
      RECT  0.82 1.055 2.005 1.145 ;
      RECT  1.885 1.145 2.005 1.45 ;
      RECT  1.885 1.45 4.835 1.56 ;
      RECT  2.095 1.0 2.21 1.25 ;
      RECT  2.095 1.25 6.08 1.36 ;
      RECT  4.895 1.0 5.015 1.25 ;
  END
END SEN_MUXI2_DG_5
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_6
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_6
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 3.85 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.325 0.71 6.05 0.89 ;
      RECT  5.95 0.89 6.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.325 0.51 7.45 0.71 ;
      RECT  6.35 0.71 7.45 0.89 ;
      RECT  0.49 0.51 0.59 0.93 ;
      LAYER M2 ;
      RECT  0.45 0.55 7.465 0.65 ;
      LAYER V1 ;
      RECT  7.325 0.55 7.425 0.65 ;
      RECT  0.49 0.55 0.59 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4848 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.105 1.255 1.225 1.75 ;
      RECT  1.625 1.255 1.745 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  5.785 1.44 5.915 1.75 ;
      RECT  6.305 1.45 6.435 1.75 ;
      RECT  6.825 1.45 6.955 1.75 ;
      RECT  7.37 1.21 7.49 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  5.785 0.05 5.915 0.36 ;
      RECT  6.305 0.05 6.435 0.36 ;
      RECT  6.825 0.05 6.955 0.36 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  7.365 0.05 7.495 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.38 0.215 5.67 0.345 ;
      RECT  3.94 0.345 4.07 1.0 ;
      RECT  2.355 1.0 5.7 1.13 ;
    END
    ANTENNADIFFAREA 1.426 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.795 0.45 3.85 0.58 ;
      RECT  4.2 0.455 7.235 0.585 ;
      RECT  0.68 0.79 1.715 0.89 ;
      RECT  0.68 0.89 0.77 1.26 ;
      RECT  0.31 0.25 0.445 0.42 ;
      RECT  0.31 0.42 0.4 1.26 ;
      RECT  0.31 1.26 0.77 1.35 ;
      RECT  0.31 1.35 0.445 1.5 ;
      RECT  0.86 1.035 2.01 1.165 ;
      RECT  1.88 1.165 2.01 1.22 ;
      RECT  0.86 1.165 0.95 1.25 ;
      RECT  1.88 1.22 5.44 1.35 ;
      RECT  5.565 1.22 7.24 1.35 ;
      RECT  5.565 1.35 5.695 1.475 ;
      RECT  2.615 1.475 5.695 1.605 ;
  END
END SEN_MUXI2_DG_6
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_DG_8
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_DG_8
  CLASS CORE ;
  FOREIGN SEN_MUXI2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 4.85 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.335 0.71 7.45 0.89 ;
      RECT  7.35 0.89 7.45 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.35 0.51 9.45 0.71 ;
      RECT  7.95 0.71 9.45 0.89 ;
      RECT  0.49 0.51 0.59 0.955 ;
      LAYER M2 ;
      RECT  0.45 0.55 9.49 0.65 ;
      LAYER V1 ;
      RECT  9.35 0.55 9.45 0.65 ;
      RECT  0.49 0.55 0.59 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.648 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  1.105 1.255 1.225 1.75 ;
      RECT  1.625 1.255 1.745 1.75 ;
      RECT  2.12 1.48 2.29 1.75 ;
      RECT  2.64 1.475 2.81 1.75 ;
      RECT  7.33 1.455 7.455 1.75 ;
      RECT  7.845 1.455 7.975 1.75 ;
      RECT  8.365 1.455 8.495 1.75 ;
      RECT  8.885 1.455 9.015 1.75 ;
      RECT  9.41 1.21 9.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  2.66 0.05 2.79 0.36 ;
      RECT  7.325 0.05 7.455 0.36 ;
      RECT  7.845 0.05 7.975 0.36 ;
      RECT  8.365 0.05 8.495 0.36 ;
      RECT  8.885 0.05 9.015 0.36 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  9.405 0.05 9.535 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.89 0.205 7.22 0.345 ;
      RECT  4.95 0.345 5.12 0.985 ;
      RECT  2.865 0.985 7.25 1.105 ;
      RECT  2.865 1.105 6.7 1.125 ;
    END
    ANTENNADIFFAREA 1.844 ;
  END X
  OBS
      LAYER M1 ;
      RECT  9.165 0.41 9.255 0.45 ;
      RECT  5.23 0.45 9.255 0.58 ;
      RECT  6.785 0.58 7.735 0.62 ;
      RECT  0.795 0.45 4.84 0.58 ;
      RECT  2.38 0.58 3.325 0.62 ;
      RECT  4.75 0.58 4.84 0.62 ;
      RECT  0.68 0.79 2.24 0.89 ;
      RECT  0.68 0.89 0.77 1.26 ;
      RECT  0.31 0.25 0.445 0.42 ;
      RECT  0.31 0.42 0.4 1.26 ;
      RECT  0.31 1.26 0.77 1.35 ;
      RECT  0.31 1.35 0.445 1.5 ;
      RECT  0.86 1.035 2.46 1.165 ;
      RECT  2.29 1.165 2.46 1.215 ;
      RECT  0.86 1.165 0.95 1.25 ;
      RECT  2.29 1.215 6.98 1.385 ;
      RECT  7.07 1.195 8.25 1.235 ;
      RECT  7.07 1.235 9.295 1.365 ;
      RECT  7.07 1.365 7.24 1.49 ;
      RECT  3.125 1.49 7.24 1.62 ;
      RECT  4.705 1.62 7.24 1.66 ;
  END
END SEN_MUXI2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_S_0P5
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_S_0P5
  CLASS CORE ;
  FOREIGN SEN_MUXI2_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.65 0.69 ;
      RECT  0.55 0.69 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.25 0.91 0.45 1.09 ;
      RECT  0.35 1.09 0.45 1.25 ;
      RECT  0.35 1.25 0.65 1.34 ;
      RECT  0.55 1.34 0.65 1.555 ;
      RECT  0.55 1.555 1.25 1.66 ;
      RECT  1.15 0.71 1.25 1.555 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.43 0.44 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.61 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.365 0.05 0.535 0.21 ;
      RECT  1.61 0.05 1.74 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.485 1.24 0.605 ;
      RECT  0.95 0.605 1.05 1.465 ;
    END
    ANTENNADIFFAREA 0.132 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.915 0.15 1.025 0.3 ;
      RECT  0.055 0.3 1.025 0.39 ;
      RECT  0.055 0.39 0.16 1.625 ;
      RECT  0.75 0.48 0.86 1.04 ;
      RECT  0.56 1.04 0.86 1.16 ;
      RECT  1.35 0.38 1.45 1.505 ;
  END
END SEN_MUXI2_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_S_1
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_S_1
  CLASS CORE ;
  FOREIGN SEN_MUXI2_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.65 0.69 ;
      RECT  0.55 0.69 0.65 0.945 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0501 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0501 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.25 0.8 0.45 0.97 ;
      RECT  0.35 0.97 0.45 1.265 ;
      RECT  0.35 1.265 0.65 1.355 ;
      RECT  0.55 1.355 0.65 1.555 ;
      RECT  0.55 1.555 1.25 1.66 ;
      RECT  1.15 0.71 1.25 1.555 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0723 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.445 0.44 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.62 1.41 1.75 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.235 0.05 0.365 0.225 ;
      RECT  1.595 0.05 1.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.31 1.25 0.49 ;
      RECT  0.95 0.49 1.05 1.415 ;
    END
    ANTENNADIFFAREA 0.24 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.68 0.14 0.79 0.32 ;
      RECT  0.055 0.32 0.79 0.41 ;
      RECT  0.055 0.41 0.16 1.635 ;
      RECT  0.745 0.5 0.86 1.055 ;
      RECT  0.55 1.055 0.86 1.175 ;
      RECT  1.35 0.265 1.45 1.215 ;
      RECT  1.35 1.215 1.495 1.385 ;
  END
END SEN_MUXI2_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_S_2
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_S_2
  CLASS CORE ;
  FOREIGN SEN_MUXI2_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.705 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.055 0.89 ;
      RECT  0.55 0.71 0.85 0.89 ;
      LAYER M2 ;
      RECT  0.51 0.75 2.09 0.85 ;
      LAYER V1 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1443 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.61 1.435 0.74 1.75 ;
      RECT  2.49 1.415 2.62 1.75 ;
      RECT  3.015 1.21 3.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  2.75 0.05 2.88 0.385 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  0.61 0.05 0.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.19 0.25 1.85 0.34 ;
      RECT  1.725 0.34 1.85 0.465 ;
      RECT  1.19 0.34 1.31 1.165 ;
      RECT  1.725 0.465 2.405 0.585 ;
      RECT  2.15 0.585 2.25 1.015 ;
      RECT  1.7 1.015 2.405 1.135 ;
    END
    ANTENNADIFFAREA 0.476 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.96 0.235 2.615 0.355 ;
      RECT  2.495 0.355 2.615 0.51 ;
      RECT  2.495 0.51 3.135 0.6 ;
      RECT  3.015 0.245 3.135 0.51 ;
      RECT  2.495 0.6 2.6 1.205 ;
      RECT  2.495 1.205 2.925 1.225 ;
      RECT  2.265 1.225 2.925 1.325 ;
      RECT  2.265 1.325 2.375 1.47 ;
      RECT  1.405 1.47 2.375 1.59 ;
      RECT  0.86 0.34 1.1 0.46 ;
      RECT  1.01 0.46 1.1 1.04 ;
      RECT  0.86 1.04 1.1 1.16 ;
      RECT  1.465 0.455 1.585 1.225 ;
      RECT  1.465 1.225 2.155 1.255 ;
      RECT  0.34 0.21 0.46 1.255 ;
      RECT  0.34 1.255 2.155 1.345 ;
  END
END SEN_MUXI2_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_S_3
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_S_3
  CLASS CORE ;
  FOREIGN SEN_MUXI2_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.54 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1578 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.65 0.89 ;
      RECT  3.55 0.89 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1578 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.66 0.89 ;
      RECT  0.81 0.71 1.11 0.89 ;
      LAYER M2 ;
      RECT  0.77 0.75 2.09 0.85 ;
      LAYER V1 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  0.81 0.75 0.91 0.85 ;
      RECT  1.01 0.75 1.11 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2172 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.225 0.45 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.845 1.415 0.975 1.75 ;
      RECT  3.215 1.435 3.345 1.75 ;
      RECT  3.77 1.21 3.89 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  0.59 0.05 0.72 0.39 ;
      RECT  1.125 0.05 1.255 0.39 ;
      RECT  3.215 0.05 3.345 0.39 ;
      RECT  3.76 0.05 3.89 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.655 0.425 1.775 0.475 ;
      RECT  1.655 0.475 2.85 0.595 ;
      RECT  2.75 0.595 2.85 1.015 ;
      RECT  1.605 1.015 2.85 1.135 ;
      RECT  1.605 1.135 1.725 1.24 ;
    END
    ANTENNADIFFAREA 0.624 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.395 0.215 2.09 0.335 ;
      RECT  1.395 0.335 1.515 1.235 ;
      RECT  0.34 0.37 0.45 0.5 ;
      RECT  0.34 0.5 0.72 0.59 ;
      RECT  0.63 0.59 0.72 1.015 ;
      RECT  0.07 1.015 0.72 1.135 ;
      RECT  0.59 1.135 0.72 1.235 ;
      RECT  0.07 1.135 0.19 1.24 ;
      RECT  0.59 1.235 1.515 1.325 ;
      RECT  1.395 1.325 1.515 1.445 ;
      RECT  1.395 1.445 2.56 1.565 ;
      RECT  2.38 0.215 3.075 0.335 ;
      RECT  2.95 0.335 3.075 0.49 ;
      RECT  2.95 0.49 3.605 0.58 ;
      RECT  3.485 0.23 3.605 0.49 ;
      RECT  2.95 0.58 3.05 1.225 ;
      RECT  1.82 1.225 3.63 1.345 ;
      RECT  0.86 0.22 0.98 0.49 ;
      RECT  0.86 0.49 1.305 0.58 ;
      RECT  1.2 0.58 1.305 1.025 ;
      RECT  1.095 1.025 1.305 1.145 ;
  END
END SEN_MUXI2_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_S_4
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_S_4
  CLASS CORE ;
  FOREIGN SEN_MUXI2_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.805 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 4.85 0.89 ;
      RECT  4.75 0.89 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 3.65 0.89 ;
      RECT  1.15 0.71 1.45 0.89 ;
      LAYER M2 ;
      RECT  1.11 0.75 2.29 0.85 ;
      LAYER V1 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2886 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.585 1.415 0.715 1.75 ;
      RECT  1.105 1.415 1.235 1.75 ;
      RECT  3.93 1.48 4.1 1.75 ;
      RECT  4.49 1.415 4.62 1.75 ;
      RECT  5.015 1.21 5.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  0.325 0.05 0.455 0.345 ;
      RECT  0.845 0.05 0.975 0.345 ;
      RECT  1.365 0.05 1.495 0.39 ;
      RECT  4.23 0.05 4.36 0.39 ;
      RECT  4.75 0.05 4.88 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.9 0.43 2.015 0.48 ;
      RECT  1.9 0.48 3.86 0.6 ;
      RECT  3.745 0.6 3.86 1.07 ;
      RECT  2.27 1.07 3.86 1.185 ;
    END
    ANTENNADIFFAREA 0.702 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.59 0.22 2.82 0.34 ;
      RECT  1.72 0.34 1.81 1.235 ;
      RECT  0.07 0.34 0.19 0.435 ;
      RECT  0.07 0.435 1.02 0.56 ;
      RECT  0.93 0.56 1.02 1.205 ;
      RECT  0.305 1.205 1.02 1.235 ;
      RECT  0.305 1.235 1.81 1.325 ;
      RECT  1.72 1.325 1.81 1.48 ;
      RECT  1.72 1.48 3.79 1.6 ;
      RECT  2.91 0.235 4.095 0.355 ;
      RECT  3.975 0.355 4.095 0.51 ;
      RECT  3.975 0.51 5.135 0.6 ;
      RECT  4.495 0.255 4.615 0.51 ;
      RECT  5.015 0.21 5.135 0.51 ;
      RECT  3.975 0.6 4.075 1.195 ;
      RECT  3.975 1.195 4.9 1.275 ;
      RECT  2.01 1.275 4.9 1.315 ;
      RECT  2.01 1.315 4.075 1.39 ;
      RECT  1.11 0.31 1.23 0.53 ;
      RECT  1.11 0.53 1.63 0.62 ;
      RECT  1.54 0.62 1.63 1.025 ;
      RECT  1.32 1.025 1.63 1.145 ;
  END
END SEN_MUXI2_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_S_6
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_S_6
  CLASS CORE ;
  FOREIGN SEN_MUXI2_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.05 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3156 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.94 0.71 6.85 0.89 ;
      RECT  6.75 0.89 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3156 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 5.08 0.89 ;
      RECT  4.98 0.89 5.08 1.09 ;
      RECT  1.345 0.63 1.745 0.74 ;
      RECT  1.645 0.74 1.745 1.09 ;
      LAYER M2 ;
      RECT  1.605 0.95 5.12 1.05 ;
      LAYER V1 ;
      RECT  4.98 0.95 5.08 1.05 ;
      RECT  1.645 0.95 1.745 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4284 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.59 1.215 0.71 1.75 ;
      RECT  1.115 1.215 1.235 1.75 ;
      RECT  1.615 1.445 1.785 1.75 ;
      RECT  2.145 1.445 2.315 1.75 ;
      RECT  5.25 1.44 5.38 1.75 ;
      RECT  5.775 1.21 5.895 1.75 ;
      RECT  6.295 1.21 6.415 1.75 ;
      RECT  6.815 1.21 6.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  1.635 0.05 1.765 0.36 ;
      RECT  0.585 0.05 0.715 0.385 ;
      RECT  1.105 0.05 1.235 0.385 ;
      RECT  5.77 0.05 5.9 0.385 ;
      RECT  6.29 0.05 6.42 0.385 ;
      RECT  6.81 0.05 6.94 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.11 0.225 3.84 0.355 ;
      RECT  3.71 0.355 3.84 0.46 ;
      RECT  3.71 0.46 5.4 0.59 ;
      RECT  3.71 0.59 3.85 1.02 ;
      RECT  2.62 1.02 4.88 1.14 ;
    END
    ANTENNADIFFAREA 1.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.93 0.235 5.64 0.355 ;
      RECT  5.51 0.355 5.64 0.485 ;
      RECT  5.51 0.485 6.675 0.595 ;
      RECT  6.035 0.26 6.155 0.485 ;
      RECT  6.555 0.26 6.675 0.485 ;
      RECT  5.51 0.595 5.64 1.0 ;
      RECT  5.51 1.0 6.66 1.12 ;
      RECT  5.51 1.12 5.635 1.23 ;
      RECT  6.555 1.12 6.66 1.23 ;
      RECT  2.85 1.23 5.635 1.35 ;
      RECT  1.38 0.28 1.5 0.45 ;
      RECT  1.38 0.45 2.295 0.54 ;
      RECT  1.9 0.3 2.02 0.45 ;
      RECT  2.195 0.54 2.295 1.015 ;
      RECT  1.85 1.015 2.295 1.135 ;
      RECT  2.395 0.455 3.6 0.575 ;
      RECT  2.395 0.575 2.525 1.225 ;
      RECT  0.305 0.485 1.25 0.605 ;
      RECT  1.15 0.605 1.25 0.995 ;
      RECT  1.15 0.995 1.505 1.005 ;
      RECT  0.34 1.005 1.505 1.125 ;
      RECT  1.375 1.125 1.505 1.225 ;
      RECT  0.34 1.125 0.45 1.29 ;
      RECT  1.375 1.225 2.525 1.355 ;
      RECT  2.405 1.355 2.525 1.44 ;
      RECT  2.405 1.44 4.65 1.56 ;
      RECT  2.615 0.735 3.51 0.89 ;
      LAYER M2 ;
      RECT  2.155 0.75 2.995 0.85 ;
      LAYER V1 ;
      RECT  2.195 0.75 2.295 0.85 ;
      RECT  2.655 0.75 2.755 0.85 ;
      RECT  2.855 0.75 2.955 0.85 ;
  END
END SEN_MUXI2_S_6
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_S_8
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_S_8
  CLASS CORE ;
  FOREIGN SEN_MUXI2_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.07 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 8.65 0.89 ;
      RECT  8.55 0.89 8.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 5.85 0.89 ;
      RECT  1.76 0.63 2.25 0.71 ;
      RECT  1.76 0.71 2.46 0.74 ;
      RECT  2.15 0.74 2.46 0.89 ;
      LAYER M2 ;
      RECT  2.11 0.75 4.09 0.85 ;
      LAYER V1 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  3.95 0.75 4.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  2.35 0.75 2.45 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5661 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.59 1.23 0.71 1.75 ;
      RECT  1.11 1.23 1.23 1.75 ;
      RECT  1.63 1.23 1.75 1.75 ;
      RECT  2.135 1.465 2.305 1.75 ;
      RECT  2.675 1.465 2.845 1.75 ;
      RECT  6.48 1.24 6.6 1.75 ;
      RECT  7.0 1.24 7.12 1.75 ;
      RECT  7.53 1.24 7.65 1.75 ;
      RECT  8.05 1.24 8.17 1.75 ;
      RECT  8.59 1.21 8.71 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  1.895 0.05 2.025 0.36 ;
      RECT  2.415 0.05 2.54 0.36 ;
      RECT  7.375 0.05 7.505 0.375 ;
      RECT  7.995 0.05 8.125 0.375 ;
      RECT  0.325 0.05 0.455 0.385 ;
      RECT  0.845 0.05 0.975 0.385 ;
      RECT  1.37 0.05 1.49 0.59 ;
      RECT  8.59 0.05 8.71 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.63 0.205 4.88 0.345 ;
      RECT  4.71 0.345 4.88 0.45 ;
      RECT  4.71 0.45 6.11 0.51 ;
      RECT  4.71 0.51 6.945 0.62 ;
      RECT  5.94 0.62 6.945 0.69 ;
      RECT  5.94 0.69 6.11 0.99 ;
      RECT  5.515 0.99 6.11 1.02 ;
      RECT  3.59 1.02 6.11 1.16 ;
    END
    ANTENNADIFFAREA 1.426 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.97 0.205 7.22 0.345 ;
      RECT  7.05 0.345 7.22 0.465 ;
      RECT  7.05 0.465 8.455 0.585 ;
      RECT  7.05 0.585 7.22 0.98 ;
      RECT  6.2 0.98 7.22 1.03 ;
      RECT  6.2 1.03 8.455 1.15 ;
      RECT  6.2 1.15 6.37 1.25 ;
      RECT  6.74 1.15 6.86 1.39 ;
      RECT  3.28 1.25 6.37 1.375 ;
      RECT  1.64 0.32 1.76 0.45 ;
      RECT  1.64 0.45 2.65 0.54 ;
      RECT  2.16 0.29 2.28 0.45 ;
      RECT  2.55 0.54 2.65 0.71 ;
      RECT  2.55 0.71 3.24 0.88 ;
      RECT  2.55 0.88 2.65 1.0 ;
      RECT  2.395 1.0 2.65 1.115 ;
      RECT  2.86 0.45 4.62 0.57 ;
      RECT  3.33 0.57 4.62 0.58 ;
      RECT  3.33 0.58 3.5 0.99 ;
      RECT  2.965 0.99 3.5 1.16 ;
      RECT  2.965 1.16 3.135 1.205 ;
      RECT  0.07 0.36 0.19 0.485 ;
      RECT  0.07 0.485 1.28 0.605 ;
      RECT  1.16 0.605 1.28 1.005 ;
      RECT  1.16 1.005 2.045 1.015 ;
      RECT  0.34 1.015 2.045 1.135 ;
      RECT  0.34 1.135 0.45 1.19 ;
      RECT  1.875 1.135 2.045 1.205 ;
      RECT  1.875 1.205 3.135 1.375 ;
      RECT  2.965 1.375 3.135 1.465 ;
      RECT  2.965 1.465 6.13 1.585 ;
  END
END SEN_MUXI2_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_D_1
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_D_1
  CLASS CORE ;
  FOREIGN SEN_MUXI2_D_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.5 1.65 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.71 0.45 0.92 ;
      RECT  0.35 0.92 0.45 1.41 ;
      RECT  0.35 1.41 0.89 1.5 ;
      RECT  0.78 1.5 0.89 1.63 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.108 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.59 0.48 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.615 1.43 1.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.355 0.05 0.485 0.37 ;
      RECT  1.62 0.05 1.74 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.93 0.505 1.055 0.69 ;
      RECT  0.965 0.69 1.055 1.015 ;
      RECT  0.95 1.015 1.055 1.1 ;
      RECT  0.95 1.1 1.285 1.29 ;
      RECT  1.15 1.29 1.285 1.515 ;
    END
    ANTENNADIFFAREA 0.236 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.74 0.29 1.37 0.38 ;
      RECT  0.74 0.38 0.835 0.51 ;
      RECT  1.275 0.38 1.37 0.94 ;
      RECT  0.07 0.32 0.175 0.51 ;
      RECT  0.07 0.51 0.835 0.6 ;
      RECT  0.74 0.6 0.835 0.77 ;
      RECT  0.07 0.6 0.17 1.44 ;
      RECT  0.74 0.77 0.875 0.94 ;
  END
END SEN_MUXI2_D_1
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_D_2
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_D_2
  CLASS CORE ;
  FOREIGN SEN_MUXI2_D_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.11 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.29 0.71 3.65 0.89 ;
      RECT  3.55 0.89 3.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.63 2.64 0.735 ;
      RECT  2.35 0.735 2.45 1.3 ;
      RECT  0.11 0.52 0.21 1.3 ;
      LAYER M2 ;
      RECT  0.07 1.15 2.49 1.25 ;
      LAYER V1 ;
      RECT  2.35 1.15 2.45 1.25 ;
      RECT  0.11 1.15 0.21 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.216 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.2 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.59 1.23 0.71 1.75 ;
      RECT  1.105 1.435 1.235 1.75 ;
      RECT  3.35 1.445 3.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  1.14 0.05 1.31 0.2 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  3.35 0.05 3.48 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.815 0.355 2.92 0.415 ;
      RECT  1.75 0.415 2.92 0.52 ;
      RECT  2.815 0.52 2.92 0.525 ;
      RECT  1.75 0.52 2.05 0.69 ;
      RECT  2.815 0.525 2.915 1.42 ;
      RECT  1.75 0.69 1.875 1.27 ;
      RECT  1.75 1.27 2.255 1.275 ;
      RECT  1.59 1.275 2.255 1.38 ;
      RECT  2.135 1.38 2.255 1.505 ;
    END
    ANTENNADIFFAREA 0.486 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.53 0.15 3.215 0.24 ;
      RECT  2.53 0.24 2.7 0.315 ;
      RECT  3.095 0.24 3.215 0.5 ;
      RECT  3.095 0.5 3.735 0.59 ;
      RECT  3.615 0.37 3.735 0.5 ;
      RECT  0.85 0.17 0.97 0.3 ;
      RECT  0.85 0.3 2.19 0.305 ;
      RECT  1.51 0.215 2.19 0.3 ;
      RECT  0.85 0.305 1.65 0.39 ;
      RECT  0.325 0.32 0.45 0.5 ;
      RECT  0.325 0.5 1.615 0.59 ;
      RECT  1.5 0.59 1.615 0.91 ;
      RECT  0.325 0.59 0.45 1.46 ;
      RECT  3.065 1.21 3.735 1.3 ;
      RECT  3.615 1.3 3.735 1.43 ;
      RECT  3.065 1.3 3.185 1.53 ;
      RECT  2.54 1.41 2.66 1.53 ;
      RECT  2.54 1.53 3.185 1.62 ;
      RECT  0.825 1.21 1.475 1.32 ;
      RECT  1.355 1.32 1.475 1.47 ;
      RECT  1.355 1.47 2.02 1.585 ;
  END
END SEN_MUXI2_D_2
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_D_4
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_D_4
  CLASS CORE ;
  FOREIGN SEN_MUXI2_D_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.71 5.85 0.89 ;
      RECT  5.75 0.89 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.94 2.85 1.07 ;
      RECT  2.15 1.07 2.25 1.21 ;
      RECT  0.315 0.71 0.86 0.89 ;
      RECT  0.74 0.89 0.86 1.01 ;
      RECT  0.74 1.01 1.05 1.1 ;
      RECT  0.95 1.1 1.05 1.21 ;
      RECT  0.95 1.21 2.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.432 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.41 0.455 1.75 ;
      RECT  0.0 1.75 6.2 1.85 ;
      RECT  0.845 1.415 0.975 1.75 ;
      RECT  1.4 1.6 1.61 1.75 ;
      RECT  2.065 1.6 2.275 1.75 ;
      RECT  5.225 1.445 5.355 1.75 ;
      RECT  5.745 1.445 5.875 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      RECT  1.4 0.05 1.61 0.2 ;
      RECT  2.05 0.05 2.18 0.38 ;
      RECT  5.225 0.05 5.355 0.38 ;
      RECT  5.745 0.05 5.875 0.38 ;
      RECT  0.325 0.05 0.455 0.39 ;
      RECT  0.845 0.05 0.975 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.14 0.415 4.855 0.52 ;
      RECT  4.75 0.52 4.855 1.21 ;
      RECT  3.655 0.33 3.775 0.47 ;
      RECT  2.56 0.47 3.775 0.57 ;
      RECT  3.15 0.57 3.25 1.21 ;
      RECT  2.58 1.21 4.855 1.33 ;
    END
    ANTENNADIFFAREA 0.883 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.34 0.21 3.565 0.31 ;
      RECT  2.34 0.31 2.46 0.47 ;
      RECT  1.085 0.29 1.9 0.39 ;
      RECT  1.78 0.39 1.9 0.47 ;
      RECT  1.78 0.47 2.46 0.59 ;
      RECT  3.87 0.205 5.09 0.31 ;
      RECT  4.97 0.31 5.09 0.47 ;
      RECT  4.97 0.47 6.13 0.59 ;
      RECT  6.01 0.37 6.13 0.47 ;
      RECT  0.07 0.41 0.19 0.48 ;
      RECT  0.07 0.48 1.66 0.59 ;
      RECT  1.54 0.59 1.66 0.74 ;
      RECT  0.07 0.59 0.185 1.21 ;
      RECT  1.54 0.74 3.015 0.85 ;
      RECT  2.415 0.71 3.015 0.74 ;
      RECT  0.07 1.21 0.76 1.31 ;
      RECT  3.95 0.5 4.05 0.695 ;
      RECT  3.95 0.695 4.47 0.9 ;
      RECT  3.34 0.9 4.05 1.1 ;
      RECT  4.97 1.21 6.13 1.33 ;
      RECT  6.01 1.33 6.13 1.43 ;
      RECT  4.97 1.33 5.09 1.465 ;
      RECT  3.88 1.465 5.09 1.57 ;
      RECT  1.065 1.39 2.495 1.475 ;
      RECT  1.065 1.475 3.58 1.51 ;
      RECT  2.365 1.51 3.58 1.59 ;
  END
END SEN_MUXI2_D_4
#-----------------------------------------------------------------------
#      Cell        : SEN_MUXI2_8
#      Description : "2-1 multiplexer with inverted output"
#      Equation    : X=!((S&D1)|(!S&D0))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_MUXI2_8
  CLASS CORE ;
  FOREIGN SEN_MUXI2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN D0
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 2.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END D0
  PIN D1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.95 0.51 10.05 0.71 ;
      RECT  8.55 0.71 10.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END D1
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.875 0.71 8.05 0.89 ;
      RECT  7.95 0.89 8.05 1.095 ;
      RECT  0.55 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
      LAYER M2 ;
      RECT  0.91 0.95 8.09 1.05 ;
      LAYER V1 ;
      RECT  7.95 0.95 8.05 1.05 ;
      RECT  0.95 0.95 1.05 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 10.2 1.85 ;
      RECT  0.6 1.45 0.73 1.75 ;
      RECT  1.12 1.45 1.25 1.75 ;
      RECT  1.64 1.455 1.77 1.75 ;
      RECT  2.16 1.455 2.29 1.75 ;
      RECT  2.66 1.48 2.83 1.75 ;
      RECT  3.18 1.475 3.35 1.75 ;
      RECT  7.925 1.455 8.055 1.75 ;
      RECT  8.445 1.455 8.575 1.75 ;
      RECT  8.965 1.455 9.095 1.75 ;
      RECT  9.485 1.455 9.615 1.75 ;
      RECT  10.01 1.21 10.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      RECT  0.6 0.05 0.73 0.345 ;
      RECT  1.12 0.05 1.25 0.36 ;
      RECT  1.64 0.05 1.77 0.36 ;
      RECT  2.16 0.05 2.29 0.36 ;
      RECT  2.68 0.05 2.81 0.36 ;
      RECT  3.2 0.05 3.325 0.36 ;
      RECT  7.915 0.05 8.045 0.36 ;
      RECT  8.445 0.05 8.575 0.36 ;
      RECT  8.965 0.05 9.095 0.36 ;
      RECT  9.485 0.05 9.615 0.36 ;
      RECT  10.005 0.05 10.135 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.43 0.205 7.76 0.345 ;
      RECT  5.49 0.345 5.66 0.985 ;
      RECT  3.43 0.985 7.76 1.105 ;
      RECT  3.43 1.105 7.24 1.125 ;
    END
    ANTENNADIFFAREA 1.87 ;
  END X
  OBS
      LAYER M1 ;
      RECT  9.75 0.36 9.855 0.45 ;
      RECT  5.77 0.45 9.855 0.58 ;
      RECT  7.325 0.58 8.335 0.62 ;
      RECT  1.36 0.45 5.38 0.58 ;
      RECT  2.92 0.58 3.865 0.62 ;
      RECT  5.29 0.58 5.38 0.62 ;
      RECT  3.09 0.785 5.39 0.895 ;
      RECT  3.09 0.895 3.19 1.025 ;
      RECT  1.22 1.025 3.19 1.125 ;
      RECT  1.22 1.125 1.31 1.24 ;
      RECT  0.32 0.44 1.01 0.56 ;
      RECT  0.32 0.56 0.42 1.24 ;
      RECT  0.32 1.24 1.31 1.36 ;
      RECT  7.625 1.195 8.85 1.235 ;
      RECT  7.625 1.235 9.895 1.365 ;
      RECT  7.625 1.365 7.795 1.49 ;
      RECT  3.66 1.49 7.795 1.62 ;
      RECT  5.245 1.62 7.795 1.66 ;
      RECT  1.4 1.215 7.5 1.345 ;
      RECT  2.83 1.345 7.5 1.385 ;
      RECT  1.4 1.345 1.49 1.45 ;
  END
END SEN_MUXI2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_0P5
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_0P5
  CLASS CORE ;
  FOREIGN SEN_ND2_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.5 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.615 1.41 0.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.065 0.05 0.185 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.6 0.17 0.72 0.3 ;
      RECT  0.35 0.3 0.72 0.39 ;
      RECT  0.35 0.39 0.45 1.52 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
END SEN_ND2_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_1
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_1
  CLASS CORE ;
  FOREIGN SEN_ND2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.5 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.615 1.21 0.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.065 0.05 0.185 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.6 0.17 0.72 0.3 ;
      RECT  0.35 0.3 0.72 0.39 ;
      RECT  0.35 0.39 0.45 1.3 ;
    END
    ANTENNADIFFAREA 0.197 ;
  END X
END SEN_ND2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_12
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_12
  CLASS CORE ;
  FOREIGN SEN_ND2_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.65 0.8 ;
      RECT  0.15 0.8 2.2 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.545 0.71 6.45 0.77 ;
      RECT  3.91 0.77 6.45 0.89 ;
      RECT  6.35 0.89 6.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.115 1.41 0.235 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.64 1.41 0.76 1.75 ;
      RECT  1.16 1.41 1.28 1.75 ;
      RECT  1.68 1.41 1.8 1.75 ;
      RECT  2.2 1.415 2.32 1.75 ;
      RECT  2.72 1.41 2.84 1.75 ;
      RECT  3.255 1.42 3.375 1.75 ;
      RECT  3.79 1.42 3.91 1.75 ;
      RECT  4.31 1.42 4.43 1.75 ;
      RECT  4.82 1.405 4.955 1.75 ;
      RECT  5.35 1.415 5.47 1.75 ;
      RECT  5.87 1.42 5.99 1.75 ;
      RECT  6.395 1.415 6.515 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  3.505 0.05 3.675 0.32 ;
      RECT  4.025 0.05 4.195 0.32 ;
      RECT  4.545 0.05 4.715 0.32 ;
      RECT  5.09 0.05 5.21 0.355 ;
      RECT  5.61 0.05 5.73 0.355 ;
      RECT  6.125 0.05 6.255 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.335 0.42 2.085 0.51 ;
      RECT  0.335 0.51 3.095 0.55 ;
      RECT  1.75 0.55 3.095 0.69 ;
      RECT  2.33 0.69 3.05 0.73 ;
      RECT  2.75 0.73 3.05 1.04 ;
      RECT  2.75 1.04 4.435 1.07 ;
      RECT  2.33 1.07 4.435 1.11 ;
      RECT  0.35 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 2.016 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.655 0.16 3.415 0.2 ;
      RECT  0.12 0.2 3.415 0.33 ;
      RECT  2.195 0.33 3.415 0.39 ;
      RECT  0.12 0.33 0.24 0.42 ;
      RECT  3.185 0.39 3.415 0.41 ;
      RECT  3.185 0.41 4.98 0.45 ;
      RECT  3.185 0.45 6.51 0.58 ;
      RECT  6.39 0.36 6.51 0.45 ;
      RECT  3.185 0.58 4.47 0.64 ;
  END
END SEN_ND2_12
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_16
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_16
  CLASS CORE ;
  FOREIGN SEN_ND2_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 2.285 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.065 0.71 8.45 0.785 ;
      RECT  5.07 0.785 8.45 0.89 ;
      RECT  8.35 0.89 8.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.585 1.41 0.705 1.75 ;
      RECT  1.105 1.41 1.225 1.75 ;
      RECT  1.625 1.41 1.745 1.75 ;
      RECT  2.155 1.415 2.285 1.75 ;
      RECT  2.655 1.48 2.825 1.75 ;
      RECT  3.175 1.48 3.345 1.75 ;
      RECT  3.695 1.48 3.865 1.75 ;
      RECT  4.215 1.48 4.385 1.75 ;
      RECT  4.735 1.48 4.905 1.75 ;
      RECT  5.255 1.48 5.425 1.75 ;
      RECT  5.775 1.46 5.945 1.75 ;
      RECT  6.31 1.415 6.445 1.75 ;
      RECT  6.83 1.415 6.965 1.75 ;
      RECT  7.35 1.415 7.485 1.75 ;
      RECT  7.87 1.415 8.005 1.75 ;
      RECT  8.4 1.21 8.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  4.475 0.05 4.645 0.32 ;
      RECT  4.995 0.05 5.165 0.32 ;
      RECT  5.515 0.05 5.685 0.32 ;
      RECT  6.035 0.05 6.205 0.32 ;
      RECT  6.555 0.05 6.725 0.32 ;
      RECT  7.075 0.05 7.245 0.32 ;
      RECT  7.595 0.05 7.765 0.32 ;
      RECT  8.115 0.05 8.285 0.32 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.3 0.445 2.565 0.51 ;
      RECT  0.3 0.51 3.13 0.575 ;
      RECT  1.855 0.575 3.6 0.615 ;
      RECT  2.38 0.615 3.6 0.62 ;
      RECT  2.38 0.62 4.11 0.72 ;
      RECT  3.94 0.56 4.11 0.62 ;
      RECT  2.38 0.72 3.66 0.74 ;
      RECT  2.94 0.74 3.66 0.89 ;
      RECT  3.34 0.89 3.66 1.07 ;
      RECT  3.34 1.07 4.665 1.1 ;
      RECT  3.34 1.1 5.26 1.11 ;
      RECT  0.34 1.11 8.26 1.29 ;
      RECT  2.395 1.29 6.205 1.33 ;
      RECT  2.395 1.33 5.695 1.36 ;
      RECT  2.395 1.36 5.26 1.39 ;
    END
    ANTENNADIFFAREA 2.696 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.75 0.31 4.88 0.41 ;
      RECT  4.75 0.41 8.52 0.49 ;
      RECT  8.4 0.32 8.52 0.41 ;
      RECT  1.595 0.16 3.89 0.2 ;
      RECT  0.065 0.2 3.89 0.26 ;
      RECT  0.065 0.26 4.385 0.32 ;
      RECT  2.13 0.32 4.385 0.355 ;
      RECT  0.065 0.32 0.19 0.42 ;
      RECT  2.645 0.355 4.385 0.4 ;
      RECT  3.2 0.4 4.385 0.45 ;
      RECT  4.2 0.45 4.385 0.49 ;
      RECT  4.2 0.49 8.52 0.54 ;
      RECT  4.2 0.54 6.975 0.58 ;
      RECT  4.2 0.58 6.46 0.605 ;
      RECT  4.2 0.605 5.94 0.645 ;
      RECT  4.2 0.645 5.325 0.68 ;
      LAYER M2 ;
      RECT  3.21 0.35 4.91 0.45 ;
      LAYER V1 ;
      RECT  3.255 0.35 3.355 0.45 ;
      RECT  3.75 0.35 3.85 0.45 ;
      RECT  4.24 0.35 4.34 0.45 ;
      RECT  4.77 0.35 4.87 0.45 ;
  END
END SEN_ND2_16
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_2
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_2
  CLASS CORE ;
  FOREIGN SEN_ND2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.64 1.41 0.76 1.75 ;
      RECT  1.205 1.41 1.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.94 0.05 1.06 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.42 0.45 0.475 ;
      RECT  0.35 0.475 0.65 0.59 ;
      RECT  0.55 0.59 0.65 1.11 ;
      RECT  0.35 1.11 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.2 0.85 0.32 ;
      RECT  0.08 0.32 0.2 0.39 ;
      RECT  0.75 0.32 0.85 0.5 ;
      RECT  0.75 0.5 1.32 0.59 ;
      RECT  1.2 0.37 1.32 0.5 ;
  END
END SEN_ND2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_3
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_3
  CLASS CORE ;
  FOREIGN SEN_ND2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.5 1.65 0.71 ;
      RECT  1.15 0.71 1.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.175 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.565 1.42 0.69 1.75 ;
      RECT  1.095 1.42 1.22 1.75 ;
      RECT  1.62 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.1 0.05 1.22 0.39 ;
      RECT  1.62 0.05 1.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.055 0.19 0.175 0.435 ;
      RECT  0.055 0.435 0.83 0.555 ;
      RECT  0.74 0.555 0.83 0.63 ;
      RECT  0.74 0.63 0.85 1.21 ;
      RECT  0.29 1.21 1.51 1.33 ;
    END
    ANTENNADIFFAREA 0.529 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.355 0.21 1.48 0.385 ;
      RECT  1.355 0.385 1.45 0.48 ;
      RECT  0.29 0.225 1.01 0.345 ;
      RECT  0.92 0.345 1.01 0.48 ;
      RECT  0.92 0.48 1.45 0.57 ;
  END
END SEN_ND2_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_4
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_4
  CLASS CORE ;
  FOREIGN SEN_ND2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.7 2.25 0.9 ;
      RECT  2.15 0.9 2.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.585 1.41 0.705 1.75 ;
      RECT  1.105 1.41 1.225 1.75 ;
      RECT  1.625 1.41 1.745 1.75 ;
      RECT  2.165 1.41 2.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.36 0.05 1.485 0.375 ;
      RECT  1.885 0.05 2.005 0.375 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.3 0.44 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.11 ;
      RECT  0.34 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.215 1.25 0.335 ;
      RECT  0.065 0.335 0.18 0.44 ;
      RECT  1.16 0.335 1.25 0.465 ;
      RECT  1.16 0.465 2.32 0.585 ;
  END
END SEN_ND2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_6
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_6
  CLASS CORE ;
  FOREIGN SEN_ND2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.41 0.2 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.6 1.41 0.72 1.75 ;
      RECT  1.12 1.41 1.24 1.75 ;
      RECT  1.64 1.41 1.76 1.75 ;
      RECT  2.16 1.41 2.28 1.75 ;
      RECT  2.68 1.41 2.8 1.75 ;
      RECT  3.2 1.41 3.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  1.895 0.05 2.025 0.375 ;
      RECT  2.415 0.05 2.545 0.375 ;
      RECT  2.935 0.05 3.065 0.375 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.445 1.5 0.575 ;
      RECT  0.34 0.575 0.46 0.615 ;
      RECT  1.35 0.575 1.5 1.11 ;
      RECT  0.35 1.11 3.05 1.29 ;
    END
    ANTENNADIFFAREA 1.008 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.21 1.765 0.33 ;
      RECT  0.075 0.33 0.205 0.39 ;
      RECT  1.635 0.33 1.765 0.47 ;
      RECT  1.635 0.47 3.32 0.59 ;
      RECT  3.2 0.37 3.32 0.47 ;
  END
END SEN_ND2_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_8
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_8
  CLASS CORE ;
  FOREIGN SEN_ND2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.585 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.7 4.25 0.9 ;
      RECT  4.15 0.9 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.175 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.575 1.41 0.695 1.75 ;
      RECT  1.095 1.41 1.215 1.75 ;
      RECT  1.615 1.41 1.74 1.75 ;
      RECT  2.13 1.41 2.25 1.75 ;
      RECT  2.655 1.41 2.775 1.75 ;
      RECT  3.175 1.41 3.295 1.75 ;
      RECT  3.695 1.41 3.815 1.75 ;
      RECT  4.215 1.41 4.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  2.37 0.05 2.54 0.325 ;
      RECT  2.91 0.05 3.04 0.365 ;
      RECT  3.43 0.05 3.56 0.37 ;
      RECT  3.95 0.05 4.08 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.29 0.42 1.995 0.56 ;
      RECT  1.68 0.56 1.995 0.6 ;
      RECT  1.68 0.6 1.85 1.11 ;
      RECT  0.35 1.11 4.06 1.18 ;
      RECT  0.245 1.18 4.06 1.29 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.59 0.18 2.27 0.2 ;
      RECT  0.065 0.2 2.27 0.33 ;
      RECT  0.065 0.33 0.175 0.43 ;
      RECT  2.12 0.33 2.27 0.435 ;
      RECT  2.12 0.435 2.805 0.465 ;
      RECT  2.12 0.465 4.335 0.585 ;
      RECT  4.215 0.36 4.335 0.465 ;
  END
END SEN_ND2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_12
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_12
  CLASS CORE ;
  FOREIGN SEN_ND2_S_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.51 6.05 0.98 ;
      RECT  4.75 0.51 4.85 0.98 ;
      RECT  3.75 0.51 3.85 0.98 ;
      RECT  2.75 0.51 2.85 0.945 ;
      RECT  1.55 0.51 1.65 0.98 ;
      RECT  0.55 0.51 0.65 0.98 ;
      LAYER M2 ;
      RECT  0.51 0.55 6.09 0.65 ;
      LAYER V1 ;
      RECT  5.95 0.55 6.05 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5766 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.14 6.25 0.23 ;
      RECT  5.55 0.23 5.65 0.71 ;
      RECT  6.15 0.23 6.25 0.71 ;
      RECT  4.545 0.14 5.25 0.23 ;
      RECT  4.545 0.23 4.65 0.71 ;
      RECT  5.15 0.23 5.25 0.71 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.95 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.91 ;
      RECT  0.94 0.71 1.45 0.91 ;
      RECT  1.95 0.71 2.45 0.91 ;
      RECT  2.95 0.71 3.47 0.91 ;
      RECT  3.95 0.71 4.65 0.91 ;
      RECT  5.15 0.71 5.65 0.91 ;
      RECT  6.15 0.71 6.45 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5766 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.075 1.415 1.205 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.62 1.415 1.75 1.75 ;
      RECT  2.14 1.415 2.27 1.75 ;
      RECT  2.66 1.415 2.79 1.75 ;
      RECT  3.18 1.415 3.31 1.75 ;
      RECT  3.7 1.415 3.83 1.75 ;
      RECT  4.25 1.415 4.38 1.75 ;
      RECT  4.825 1.415 4.955 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  3.185 0.05 3.29 0.585 ;
      RECT  4.255 0.05 4.375 0.585 ;
      RECT  5.34 0.05 5.46 0.585 ;
      RECT  6.415 0.05 6.535 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.32 6.015 0.42 ;
      RECT  5.75 0.42 5.85 1.11 ;
      RECT  4.78 0.32 5.05 0.42 ;
      RECT  4.95 0.42 5.05 1.11 ;
      RECT  3.56 0.32 3.85 0.42 ;
      RECT  3.56 0.42 3.66 1.035 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.035 ;
      RECT  2.55 1.035 3.66 1.11 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.75 1.11 5.85 1.29 ;
    END
    ANTENNADIFFAREA 1.346 ;
  END X
END SEN_ND2_S_12
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_16
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_16
  CLASS CORE ;
  FOREIGN SEN_ND2_S_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.51 8.05 0.96 ;
      RECT  6.75 0.51 6.85 0.96 ;
      RECT  5.75 0.51 5.85 0.95 ;
      RECT  4.75 0.51 4.85 0.96 ;
      RECT  3.75 0.51 3.85 0.96 ;
      RECT  2.75 0.51 2.85 0.95 ;
      RECT  1.55 0.51 1.65 0.96 ;
      RECT  0.55 0.51 0.65 0.96 ;
      LAYER M2 ;
      RECT  0.51 0.55 8.09 0.65 ;
      LAYER V1 ;
      RECT  7.95 0.55 8.05 0.65 ;
      RECT  6.75 0.55 6.85 0.65 ;
      RECT  5.75 0.55 5.85 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7686 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.57 0.14 8.25 0.23 ;
      RECT  7.57 0.23 7.66 0.71 ;
      RECT  8.15 0.23 8.25 0.71 ;
      RECT  6.55 0.14 7.25 0.23 ;
      RECT  6.55 0.23 6.65 0.71 ;
      RECT  7.15 0.23 7.25 0.71 ;
      RECT  5.55 0.14 6.25 0.23 ;
      RECT  5.55 0.23 5.65 0.71 ;
      RECT  6.15 0.23 6.25 0.71 ;
      RECT  4.455 0.14 5.21 0.23 ;
      RECT  4.455 0.23 4.56 0.71 ;
      RECT  5.12 0.23 5.21 0.71 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.945 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  3.945 0.71 4.56 0.895 ;
      RECT  5.12 0.71 5.65 0.895 ;
      RECT  6.15 0.71 6.65 0.89 ;
      RECT  7.15 0.71 7.66 0.89 ;
      RECT  8.15 0.71 8.47 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7686 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.595 1.41 1.725 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.18 1.41 3.31 1.75 ;
      RECT  3.68 1.48 3.85 1.75 ;
      RECT  4.2 1.48 4.37 1.75 ;
      RECT  4.72 1.48 4.89 1.75 ;
      RECT  5.28 1.41 5.41 1.75 ;
      RECT  5.8 1.41 5.93 1.75 ;
      RECT  6.345 1.415 6.475 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  3.185 0.05 3.29 0.585 ;
      RECT  4.225 0.05 4.345 0.585 ;
      RECT  5.3 0.05 5.405 0.585 ;
      RECT  6.34 0.05 6.445 0.585 ;
      RECT  7.365 0.05 7.48 0.585 ;
      RECT  8.405 0.05 8.525 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.32 8.03 0.42 ;
      RECT  7.75 0.42 7.85 1.11 ;
      RECT  6.8 0.32 7.05 0.42 ;
      RECT  6.95 0.42 7.05 1.06 ;
      RECT  5.78 0.32 6.05 0.42 ;
      RECT  5.95 0.42 6.05 1.04 ;
      RECT  4.72 0.32 5.03 0.42 ;
      RECT  4.94 0.42 5.03 1.04 ;
      RECT  4.94 1.04 6.05 1.06 ;
      RECT  4.94 1.06 7.05 1.075 ;
      RECT  3.56 0.32 3.85 0.42 ;
      RECT  3.56 0.42 3.65 1.04 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.04 ;
      RECT  2.55 1.04 3.65 1.06 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.06 ;
      RECT  1.75 1.06 3.65 1.075 ;
      RECT  1.75 1.075 7.05 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.75 1.11 7.85 1.29 ;
      RECT  3.4 1.29 5.19 1.39 ;
    END
    ANTENNADIFFAREA 1.806 ;
  END X
END SEN_ND2_S_16
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_6
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_6
  CLASS CORE ;
  FOREIGN SEN_ND2_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 0.96 ;
      RECT  1.55 0.51 1.65 1.02 ;
      RECT  0.55 0.51 0.65 0.96 ;
      LAYER M2 ;
      RECT  0.51 0.55 2.89 0.65 ;
      LAYER V1 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.288 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.288 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.54 1.21 0.66 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.74 1.21 2.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  3.185 0.05 3.305 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.11 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.75 1.11 2.65 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
END SEN_ND2_S_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_8
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_8
  CLASS CORE ;
  FOREIGN SEN_ND2_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.51 3.85 0.96 ;
      RECT  2.75 0.51 2.85 0.98 ;
      RECT  1.55 0.51 1.65 1.0 ;
      RECT  0.55 0.51 0.65 0.98 ;
      LAYER M2 ;
      RECT  0.51 0.55 3.89 0.65 ;
      LAYER V1 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3834 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.95 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  3.95 0.71 4.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3834 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.555 1.41 0.685 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.205 1.41 3.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  4.225 0.05 4.345 0.385 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  3.185 0.05 3.29 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.32 3.85 0.42 ;
      RECT  3.56 0.42 3.66 1.11 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.11 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.75 1.11 3.66 1.29 ;
    END
    ANTENNADIFFAREA 0.894 ;
  END X
END SEN_ND2_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_12
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_12
  CLASS CORE ;
  FOREIGN SEN_ND2_G_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.51 6.05 0.96 ;
      RECT  4.75 0.51 4.85 0.96 ;
      RECT  3.75 0.51 3.85 0.96 ;
      RECT  2.75 0.51 2.85 0.93 ;
      RECT  1.55 0.51 1.65 0.96 ;
      RECT  0.55 0.51 0.65 0.96 ;
      LAYER M2 ;
      RECT  0.51 0.55 6.09 0.65 ;
      LAYER V1 ;
      RECT  5.95 0.55 6.05 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.14 6.25 0.23 ;
      RECT  5.55 0.23 5.65 0.71 ;
      RECT  6.15 0.23 6.25 0.71 ;
      RECT  4.545 0.14 5.25 0.23 ;
      RECT  4.545 0.23 4.65 0.71 ;
      RECT  5.15 0.23 5.25 0.71 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.95 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  3.95 0.71 4.65 0.895 ;
      RECT  5.15 0.71 5.65 0.895 ;
      RECT  6.15 0.71 6.45 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.18 1.41 3.31 1.75 ;
      RECT  3.7 1.41 3.83 1.75 ;
      RECT  4.25 1.41 4.38 1.75 ;
      RECT  4.8 1.41 4.93 1.75 ;
      RECT  5.335 1.41 5.465 1.75 ;
      RECT  5.865 1.41 5.995 1.75 ;
      RECT  6.41 1.21 6.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  3.185 0.05 3.29 0.585 ;
      RECT  4.255 0.05 4.375 0.585 ;
      RECT  5.34 0.05 5.46 0.585 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.41 0.05 6.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.32 6.015 0.42 ;
      RECT  5.75 0.42 5.85 1.11 ;
      RECT  4.78 0.32 5.05 0.42 ;
      RECT  4.95 0.42 5.05 1.11 ;
      RECT  3.56 0.32 3.85 0.42 ;
      RECT  3.56 0.42 3.66 1.035 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.035 ;
      RECT  2.55 1.035 3.66 1.11 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.3 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 2.016 ;
  END X
END SEN_ND2_G_12
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_16
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_16
  CLASS CORE ;
  FOREIGN SEN_ND2_G_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.51 8.05 0.96 ;
      RECT  6.75 0.51 6.85 0.96 ;
      RECT  5.75 0.51 5.85 0.93 ;
      RECT  4.75 0.51 4.85 0.96 ;
      RECT  3.75 0.51 3.85 0.96 ;
      RECT  2.75 0.51 2.85 0.93 ;
      RECT  1.55 0.51 1.65 0.96 ;
      RECT  0.55 0.51 0.65 0.96 ;
      LAYER M2 ;
      RECT  0.51 0.55 8.09 0.65 ;
      LAYER V1 ;
      RECT  7.95 0.55 8.05 0.65 ;
      RECT  6.75 0.55 6.85 0.65 ;
      RECT  5.75 0.55 5.85 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.57 0.14 8.25 0.23 ;
      RECT  7.57 0.23 7.66 0.71 ;
      RECT  8.15 0.23 8.25 0.71 ;
      RECT  6.55 0.14 7.25 0.23 ;
      RECT  6.55 0.23 6.65 0.71 ;
      RECT  7.15 0.23 7.25 0.71 ;
      RECT  5.55 0.14 6.25 0.23 ;
      RECT  5.55 0.23 5.65 0.71 ;
      RECT  6.15 0.23 6.25 0.71 ;
      RECT  4.455 0.14 5.21 0.23 ;
      RECT  4.455 0.23 4.56 0.71 ;
      RECT  5.12 0.23 5.21 0.71 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.945 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  3.945 0.71 4.56 0.895 ;
      RECT  5.12 0.71 5.65 0.895 ;
      RECT  6.15 0.71 6.65 0.89 ;
      RECT  7.15 0.71 7.66 0.89 ;
      RECT  8.15 0.71 8.47 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.18 1.41 3.31 1.75 ;
      RECT  3.68 1.48 3.85 1.75 ;
      RECT  4.2 1.48 4.37 1.75 ;
      RECT  4.72 1.48 4.89 1.75 ;
      RECT  5.28 1.41 5.41 1.75 ;
      RECT  5.8 1.41 5.93 1.75 ;
      RECT  6.32 1.41 6.45 1.75 ;
      RECT  6.84 1.41 6.97 1.75 ;
      RECT  7.36 1.41 7.49 1.75 ;
      RECT  7.88 1.41 8.01 1.75 ;
      RECT  8.405 1.21 8.525 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  3.185 0.05 3.29 0.585 ;
      RECT  4.225 0.05 4.345 0.585 ;
      RECT  5.3 0.05 5.405 0.585 ;
      RECT  6.34 0.05 6.445 0.585 ;
      RECT  7.365 0.05 7.48 0.585 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  8.405 0.05 8.525 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.32 8.03 0.42 ;
      RECT  7.75 0.42 7.85 1.11 ;
      RECT  6.8 0.32 7.05 0.42 ;
      RECT  6.95 0.42 7.05 1.06 ;
      RECT  5.78 0.32 6.05 0.42 ;
      RECT  5.95 0.42 6.05 1.04 ;
      RECT  4.72 0.32 5.03 0.42 ;
      RECT  4.94 0.42 5.03 1.04 ;
      RECT  4.94 1.04 6.05 1.06 ;
      RECT  4.94 1.06 7.05 1.075 ;
      RECT  3.56 0.32 3.85 0.42 ;
      RECT  3.56 0.42 3.65 1.04 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.04 ;
      RECT  2.55 1.04 3.65 1.06 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.06 ;
      RECT  1.75 1.06 3.65 1.075 ;
      RECT  1.75 1.075 7.05 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.3 1.11 8.29 1.29 ;
      RECT  3.4 1.29 5.19 1.39 ;
    END
    ANTENNADIFFAREA 2.7 ;
  END X
END SEN_ND2_G_16
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_24
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_24
  CLASS CORE ;
  FOREIGN SEN_ND2_G_24 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.15 0.51 12.25 0.96 ;
      RECT  10.95 0.51 11.05 0.96 ;
      RECT  9.95 0.51 10.05 0.95 ;
      RECT  8.95 0.51 9.05 0.95 ;
      RECT  7.95 0.51 8.05 0.95 ;
      RECT  6.94 0.51 7.06 0.885 ;
      RECT  5.74 0.51 5.86 0.885 ;
      RECT  4.75 0.51 4.85 0.93 ;
      RECT  3.75 0.51 3.85 0.93 ;
      RECT  2.75 0.51 2.85 0.95 ;
      RECT  1.55 0.51 1.65 0.96 ;
      RECT  0.55 0.51 0.65 0.96 ;
      LAYER M2 ;
      RECT  0.51 0.55 12.29 0.65 ;
      LAYER V1 ;
      RECT  12.15 0.55 12.25 0.65 ;
      RECT  10.95 0.55 11.05 0.65 ;
      RECT  9.95 0.55 10.05 0.65 ;
      RECT  8.95 0.55 9.05 0.65 ;
      RECT  7.95 0.55 8.05 0.65 ;
      RECT  6.95 0.55 7.05 0.65 ;
      RECT  5.75 0.55 5.85 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5552 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.75 0.14 12.45 0.23 ;
      RECT  11.75 0.23 11.85 0.71 ;
      RECT  12.35 0.23 12.45 0.71 ;
      RECT  10.75 0.14 11.45 0.23 ;
      RECT  10.75 0.23 10.85 0.71 ;
      RECT  11.35 0.23 11.45 0.71 ;
      RECT  9.75 0.14 10.415 0.23 ;
      RECT  9.75 0.23 9.85 0.71 ;
      RECT  10.325 0.23 10.415 0.71 ;
      RECT  8.55 0.14 9.325 0.23 ;
      RECT  8.55 0.23 8.65 0.71 ;
      RECT  9.235 0.23 9.325 0.71 ;
      RECT  7.57 0.14 8.25 0.23 ;
      RECT  7.57 0.23 7.66 0.71 ;
      RECT  8.15 0.23 8.25 0.71 ;
      RECT  6.55 0.14 7.25 0.23 ;
      RECT  6.55 0.23 6.65 0.71 ;
      RECT  7.15 0.23 7.25 0.71 ;
      RECT  5.55 0.14 6.25 0.23 ;
      RECT  5.55 0.23 5.65 0.71 ;
      RECT  6.15 0.23 6.25 0.71 ;
      RECT  4.455 0.14 5.21 0.23 ;
      RECT  4.455 0.23 4.56 0.71 ;
      RECT  5.12 0.23 5.21 0.71 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.945 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  3.945 0.71 4.56 0.895 ;
      RECT  5.12 0.71 5.65 0.865 ;
      RECT  6.15 0.71 6.65 0.865 ;
      RECT  7.15 0.71 7.66 0.865 ;
      RECT  8.15 0.71 8.65 0.89 ;
      RECT  9.235 0.71 9.85 0.89 ;
      RECT  10.325 0.71 10.85 0.89 ;
      RECT  11.35 0.71 11.85 0.89 ;
      RECT  12.35 0.71 12.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5552 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.18 1.41 3.31 1.75 ;
      RECT  3.7 1.435 3.83 1.75 ;
      RECT  4.22 1.435 4.35 1.75 ;
      RECT  4.74 1.435 4.87 1.75 ;
      RECT  5.28 1.435 5.41 1.75 ;
      RECT  5.8 1.435 5.93 1.75 ;
      RECT  6.32 1.435 6.45 1.75 ;
      RECT  6.84 1.435 6.97 1.75 ;
      RECT  7.36 1.435 7.49 1.75 ;
      RECT  7.88 1.44 8.01 1.75 ;
      RECT  8.4 1.44 8.53 1.75 ;
      RECT  8.92 1.44 9.05 1.75 ;
      RECT  9.45 1.41 9.58 1.75 ;
      RECT  9.98 1.41 10.11 1.75 ;
      RECT  10.5 1.41 10.63 1.75 ;
      RECT  11.02 1.41 11.15 1.75 ;
      RECT  11.54 1.41 11.67 1.75 ;
      RECT  12.06 1.41 12.19 1.75 ;
      RECT  12.6 1.21 12.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  3.185 0.05 3.29 0.585 ;
      RECT  4.225 0.05 4.345 0.585 ;
      RECT  5.3 0.05 5.405 0.585 ;
      RECT  6.34 0.05 6.445 0.585 ;
      RECT  7.365 0.05 7.48 0.585 ;
      RECT  8.345 0.05 8.46 0.585 ;
      RECT  9.455 0.05 9.575 0.585 ;
      RECT  10.505 0.05 10.625 0.585 ;
      RECT  11.545 0.05 11.66 0.585 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  12.6 0.05 12.72 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  11.95 0.32 12.21 0.42 ;
      RECT  11.95 0.42 12.05 1.11 ;
      RECT  11.0 0.32 11.25 0.42 ;
      RECT  11.15 0.42 11.25 1.11 ;
      RECT  9.96 0.32 10.235 0.42 ;
      RECT  10.145 0.42 10.235 1.045 ;
      RECT  8.75 0.32 9.07 0.42 ;
      RECT  8.75 0.42 8.85 1.045 ;
      RECT  7.75 0.32 8.03 0.42 ;
      RECT  7.75 0.42 7.85 0.975 ;
      RECT  6.75 0.32 6.99 0.42 ;
      RECT  6.75 0.42 6.85 0.975 ;
      RECT  5.78 0.32 6.05 0.42 ;
      RECT  5.95 0.42 6.05 0.975 ;
      RECT  4.72 0.32 5.03 0.42 ;
      RECT  4.94 0.42 5.03 0.975 ;
      RECT  4.94 0.975 7.85 1.04 ;
      RECT  3.56 0.32 3.85 0.42 ;
      RECT  3.56 0.42 3.65 1.04 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.04 ;
      RECT  2.55 1.04 7.85 1.045 ;
      RECT  2.55 1.045 10.235 1.06 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.06 ;
      RECT  1.75 1.06 10.235 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.3 1.11 12.45 1.29 ;
      RECT  3.38 1.29 9.38 1.345 ;
      RECT  7.8 1.345 9.38 1.35 ;
    END
    ANTENNADIFFAREA 4.044 ;
  END X
END SEN_ND2_G_24
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_6
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_6
  CLASS CORE ;
  FOREIGN SEN_ND2_G_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 0.96 ;
      RECT  1.55 0.51 1.65 0.96 ;
      RECT  0.55 0.51 0.65 0.96 ;
      LAYER M2 ;
      RECT  0.51 0.55 2.89 0.65 ;
      LAYER V1 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.2 1.21 3.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.2 0.05 3.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.11 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.3 1.11 3.05 1.29 ;
    END
    ANTENNADIFFAREA 1.008 ;
  END X
END SEN_ND2_G_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_8
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_8
  CLASS CORE ;
  FOREIGN SEN_ND2_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.51 3.85 0.96 ;
      RECT  2.75 0.51 2.85 0.96 ;
      RECT  1.55 0.51 1.65 0.96 ;
      RECT  0.55 0.51 0.65 0.96 ;
      LAYER M2 ;
      RECT  0.51 0.55 3.89 0.65 ;
      LAYER V1 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.95 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  3.95 0.71 4.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.14 1.41 2.27 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.18 1.41 3.31 1.75 ;
      RECT  3.7 1.41 3.83 1.75 ;
      RECT  4.22 1.41 4.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  4.22 0.05 4.345 0.39 ;
      RECT  1.12 0.05 1.225 0.585 ;
      RECT  2.145 0.05 2.26 0.585 ;
      RECT  3.185 0.05 3.29 0.585 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.32 3.85 0.42 ;
      RECT  3.56 0.42 3.66 1.11 ;
      RECT  2.55 0.32 2.81 0.42 ;
      RECT  2.55 0.42 2.65 1.11 ;
      RECT  1.6 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.56 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.3 1.11 4.085 1.29 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
END SEN_ND2_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_0P65
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_0P65
  CLASS CORE ;
  FOREIGN SEN_ND2_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0402 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0402 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.18 0.2 0.27 ;
      RECT  0.08 0.27 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.122 ;
  END X
END SEN_ND2_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_0P8
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_0P8
  CLASS CORE ;
  FOREIGN SEN_ND2_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0495 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0495 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.17 0.2 0.27 ;
      RECT  0.08 0.27 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.15 ;
  END X
END SEN_ND2_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_1P5
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_1P5
  CLASS CORE ;
  FOREIGN SEN_ND2_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0918 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0918 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.635 1.41 0.765 1.75 ;
      RECT  1.2 1.21 1.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.925 0.05 1.055 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.435 0.65 0.555 ;
      RECT  0.55 0.555 0.65 1.11 ;
      RECT  0.35 1.11 1.05 1.29 ;
      RECT  0.35 1.29 0.45 1.49 ;
      RECT  0.95 1.29 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.274 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.21 0.83 0.33 ;
      RECT  0.08 0.33 0.2 0.39 ;
      RECT  0.74 0.33 0.83 0.495 ;
      RECT  0.74 0.495 1.32 0.585 ;
      RECT  1.2 0.33 1.32 0.495 ;
  END
END SEN_ND2_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_0P5
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_0P5
  CLASS CORE ;
  FOREIGN SEN_ND2_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0258 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0258 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.17 0.2 0.27 ;
      RECT  0.08 0.27 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.61 ;
    END
    ANTENNADIFFAREA 0.076 ;
  END X
END SEN_ND2_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_0P65
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_0P65
  CLASS CORE ;
  FOREIGN SEN_ND2_S_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.17 0.2 0.27 ;
      RECT  0.08 0.27 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.61 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END X
END SEN_ND2_S_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_0P8
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_0P8
  CLASS CORE ;
  FOREIGN SEN_ND2_S_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0384 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0384 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.17 0.2 0.27 ;
      RECT  0.08 0.27 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.58 ;
    END
    ANTENNADIFFAREA 0.112 ;
  END X
END SEN_ND2_S_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_1
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_1
  CLASS CORE ;
  FOREIGN SEN_ND2_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.17 0.2 0.27 ;
      RECT  0.08 0.27 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.51 ;
    END
    ANTENNADIFFAREA 0.141 ;
  END X
END SEN_ND2_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_1P5
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_1P5
  CLASS CORE ;
  FOREIGN SEN_ND2_S_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0714 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0714 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.415 0.48 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.94 1.415 1.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.92 0.05 1.045 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.435 0.65 0.555 ;
      RECT  0.55 0.555 0.65 1.11 ;
      RECT  0.55 1.11 0.785 1.29 ;
    END
    ANTENNADIFFAREA 0.192 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.21 0.83 0.33 ;
      RECT  0.08 0.33 0.2 0.39 ;
      RECT  0.74 0.33 0.83 0.435 ;
      RECT  0.74 0.435 1.325 0.555 ;
  END
END SEN_ND2_S_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_2
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_2
  CLASS CORE ;
  FOREIGN SEN_ND2_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.635 1.41 0.765 1.75 ;
      RECT  1.195 1.41 1.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.925 0.05 1.055 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.44 0.65 0.56 ;
      RECT  0.55 0.56 0.65 1.11 ;
      RECT  0.35 1.11 1.05 1.29 ;
      RECT  0.35 1.29 0.45 1.51 ;
      RECT  0.95 1.29 1.05 1.51 ;
    END
    ANTENNADIFFAREA 0.262 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.21 0.83 0.33 ;
      RECT  0.08 0.33 0.2 0.39 ;
      RECT  0.74 0.33 0.83 0.48 ;
      RECT  0.74 0.48 1.32 0.59 ;
      RECT  1.2 0.37 1.32 0.48 ;
  END
END SEN_ND2_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_3
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_3
  CLASS CORE ;
  FOREIGN SEN_ND2_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.144 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.144 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.28 1.21 0.4 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.4 1.21 1.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.12 0.05 1.23 0.39 ;
      RECT  1.62 0.05 1.745 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.37 0.185 0.47 ;
      RECT  0.065 0.47 0.85 0.59 ;
      RECT  0.75 0.59 0.85 1.11 ;
      RECT  0.55 1.11 1.25 1.29 ;
    END
    ANTENNADIFFAREA 0.365 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.3 0.23 1.03 0.35 ;
      RECT  0.94 0.35 1.03 0.48 ;
      RECT  0.94 0.48 1.54 0.6 ;
  END
END SEN_ND2_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_S_4
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_S_4
  CLASS CORE ;
  FOREIGN SEN_ND2_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  1.35 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.28 1.21 0.4 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.85 1.43 0.98 1.75 ;
      RECT  1.37 1.43 1.5 1.75 ;
      RECT  2.0 1.21 2.12 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.37 0.05 1.5 0.39 ;
      RECT  1.89 0.05 2.02 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.29 0.44 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.22 ;
      RECT  0.54 1.22 1.78 1.34 ;
    END
    ANTENNADIFFAREA 0.45 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.23 1.26 0.35 ;
      RECT  0.075 0.35 0.195 0.45 ;
      RECT  1.16 0.35 1.26 0.49 ;
      RECT  1.16 0.49 2.3 0.61 ;
  END
END SEN_ND2_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_0P5
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_0P5
  CLASS CORE ;
  FOREIGN SEN_ND2_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0453 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.595 1.41 0.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.17 0.2 0.27 ;
      RECT  0.08 0.27 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.56 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END X
END SEN_ND2_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_1
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_1
  CLASS CORE ;
  FOREIGN SEN_ND2_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0906 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.635 1.41 0.765 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.72 0.05 0.85 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.095 0.3 0.25 0.44 ;
      RECT  0.095 0.44 0.45 0.56 ;
      RECT  0.35 0.56 0.45 1.3 ;
    END
    ANTENNADIFFAREA 0.187 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.36 0.225 0.63 0.345 ;
      RECT  0.54 0.345 0.63 0.48 ;
      RECT  0.54 0.48 1.13 0.59 ;
      RECT  1.01 0.37 1.13 0.48 ;
  END
END SEN_ND2_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_16
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_16
  CLASS CORE ;
  FOREIGN SEN_ND2_T_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 2.25 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9873 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.75 0.71 8.85 0.91 ;
      RECT  6.15 0.91 8.85 1.055 ;
      RECT  7.355 1.055 8.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.4481 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 10.6 1.85 ;
      RECT  0.6 1.415 0.72 1.75 ;
      RECT  1.12 1.415 1.24 1.75 ;
      RECT  1.64 1.415 1.76 1.75 ;
      RECT  2.16 1.415 2.28 1.75 ;
      RECT  2.68 1.415 2.8 1.75 ;
      RECT  3.2 1.415 3.32 1.75 ;
      RECT  3.73 1.415 3.85 1.75 ;
      RECT  4.61 1.415 4.73 1.75 ;
      RECT  5.13 1.415 5.25 1.75 ;
      RECT  5.625 1.475 5.795 1.75 ;
      RECT  6.145 1.475 6.315 1.75 ;
      RECT  6.68 1.475 6.85 1.75 ;
      RECT  7.22 1.475 7.39 1.75 ;
      RECT  7.765 1.455 7.885 1.75 ;
      RECT  8.285 1.43 8.405 1.75 ;
      RECT  8.805 1.415 8.925 1.75 ;
      RECT  9.325 1.415 9.445 1.75 ;
      RECT  9.845 1.39 9.965 1.75 ;
      RECT  10.385 1.21 10.505 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.6 0.05 ;
      RECT  4.63 0.05 4.75 0.385 ;
      RECT  5.165 0.05 5.285 0.385 ;
      RECT  5.685 0.05 5.805 0.385 ;
      RECT  6.205 0.05 6.325 0.385 ;
      RECT  6.725 0.05 6.845 0.385 ;
      RECT  7.245 0.05 7.365 0.385 ;
      RECT  7.765 0.05 7.885 0.385 ;
      RECT  8.285 0.05 8.405 0.385 ;
      RECT  8.805 0.05 8.925 0.385 ;
      RECT  9.325 0.05 9.445 0.385 ;
      RECT  9.845 0.05 9.965 0.385 ;
      RECT  10.385 0.05 10.505 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.29 0.46 2.65 0.555 ;
      RECT  0.29 0.555 4.125 0.62 ;
      RECT  2.34 0.62 4.125 0.675 ;
      RECT  2.34 0.675 2.66 1.005 ;
      RECT  2.34 1.005 6.06 1.11 ;
      RECT  0.34 1.11 6.06 1.165 ;
      RECT  0.34 1.165 7.305 1.205 ;
      RECT  0.34 1.205 10.25 1.295 ;
      RECT  0.34 1.295 9.185 1.315 ;
      RECT  9.55 1.295 9.705 1.49 ;
      RECT  10.105 1.295 10.25 1.49 ;
      RECT  0.34 1.315 8.665 1.325 ;
      RECT  9.065 1.315 9.185 1.495 ;
      RECT  5.35 1.325 8.665 1.34 ;
      RECT  4.14 1.325 4.26 1.49 ;
      RECT  4.87 1.325 4.99 1.49 ;
      RECT  5.35 1.34 8.145 1.365 ;
      RECT  8.545 1.34 8.665 1.49 ;
      RECT  5.35 1.365 7.65 1.38 ;
      RECT  8.025 1.365 8.145 1.49 ;
      RECT  6.95 1.38 7.65 1.385 ;
      RECT  5.35 1.38 5.51 1.49 ;
      RECT  6.95 1.385 7.105 1.49 ;
      RECT  7.505 1.385 7.65 1.49 ;
    END
    ANTENNADIFFAREA 2.643 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.55 0.16 4.535 0.19 ;
      RECT  0.08 0.19 4.535 0.37 ;
      RECT  0.08 0.37 0.2 0.395 ;
      RECT  2.74 0.37 4.535 0.445 ;
      RECT  4.215 0.445 4.535 0.475 ;
      RECT  4.215 0.475 10.275 0.61 ;
      RECT  4.215 0.61 7.71 0.69 ;
      RECT  4.215 0.69 6.2 0.77 ;
  END
END SEN_ND2_T_16
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_1P5
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_1P5
  CLASS CORE ;
  FOREIGN SEN_ND2_T_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0918 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1356 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.6 1.4 0.72 1.75 ;
      RECT  1.18 1.21 1.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.87 0.05 0.99 0.39 ;
      RECT  1.415 0.05 1.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.39 0.45 1.11 ;
      RECT  0.35 1.11 1.05 1.31 ;
      RECT  0.35 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.244 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.17 0.72 0.28 ;
      RECT  0.08 0.28 0.2 0.39 ;
      RECT  0.6 0.28 0.72 0.48 ;
      RECT  0.6 0.48 1.31 0.6 ;
  END
END SEN_ND2_T_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_2
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_2
  CLASS CORE ;
  FOREIGN SEN_ND2_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.915 ;
      RECT  1.35 0.915 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1812 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.58 1.39 0.71 1.75 ;
      RECT  1.14 1.21 1.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.325 0.415 0.45 0.61 ;
      RECT  0.35 0.61 0.45 1.11 ;
      RECT  0.35 1.11 1.05 1.29 ;
      RECT  0.35 1.29 0.45 1.34 ;
      RECT  0.325 1.34 0.45 1.535 ;
    END
    ANTENNADIFFAREA 0.316 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.21 0.705 0.305 ;
      RECT  0.065 0.305 0.185 0.425 ;
      RECT  0.585 0.305 0.705 0.48 ;
      RECT  0.585 0.48 1.745 0.6 ;
      RECT  1.625 0.6 1.745 0.69 ;
  END
END SEN_ND2_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_3
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_3
  CLASS CORE ;
  FOREIGN SEN_ND2_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1854 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 0.91 ;
      RECT  1.15 0.91 1.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2718 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  1.13 1.415 1.25 1.75 ;
      RECT  1.67 1.415 1.79 1.75 ;
      RECT  2.19 1.23 2.31 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.14 0.05 1.26 0.385 ;
      RECT  1.67 0.05 1.79 0.385 ;
      RECT  2.21 0.05 2.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.365 0.185 0.44 ;
      RECT  0.065 0.44 0.85 0.56 ;
      RECT  0.75 0.56 0.85 1.21 ;
      RECT  0.275 1.21 2.05 1.325 ;
      RECT  1.41 1.325 1.53 1.51 ;
      RECT  1.93 1.325 2.05 1.515 ;
    END
    ANTENNADIFFAREA 0.524 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 0.23 1.04 0.35 ;
      RECT  0.95 0.35 1.04 0.48 ;
      RECT  0.95 0.48 2.1 0.6 ;
  END
END SEN_ND2_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_4
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_4
  CLASS CORE ;
  FOREIGN SEN_ND2_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.45 0.91 ;
      RECT  1.75 0.91 2.45 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3624 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  0.595 1.415 0.715 1.75 ;
      RECT  1.135 1.445 1.255 1.75 ;
      RECT  1.725 1.445 1.845 1.75 ;
      RECT  2.245 1.445 2.365 1.75 ;
      RECT  2.795 1.23 2.915 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  1.44 0.05 1.56 0.385 ;
      RECT  1.985 0.05 2.105 0.385 ;
      RECT  2.52 0.05 2.64 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.285 0.495 1.05 0.615 ;
      RECT  0.95 0.615 1.05 1.11 ;
      RECT  0.34 1.11 1.05 1.235 ;
      RECT  0.34 1.235 2.675 1.29 ;
      RECT  0.95 1.29 2.675 1.355 ;
    END
    ANTENNADIFFAREA 0.66 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.19 0.195 0.285 ;
      RECT  0.075 0.285 1.26 0.405 ;
      RECT  1.15 0.405 1.26 0.49 ;
      RECT  1.15 0.49 2.915 0.61 ;
      RECT  2.795 0.375 2.915 0.49 ;
  END
END SEN_ND2_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_5
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_5
  CLASS CORE ;
  FOREIGN SEN_ND2_T_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.05 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.309 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.25 0.9 ;
      RECT  2.15 0.9 3.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.453 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.615 1.39 0.735 1.75 ;
      RECT  1.135 1.415 1.265 1.75 ;
      RECT  1.725 1.405 1.845 1.75 ;
      RECT  2.265 1.405 2.385 1.75 ;
      RECT  2.785 1.405 2.905 1.75 ;
      RECT  3.32 1.405 3.44 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  1.725 0.05 1.845 0.385 ;
      RECT  2.265 0.05 2.385 0.385 ;
      RECT  2.785 0.05 2.905 0.385 ;
      RECT  3.325 0.05 3.445 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.045 0.47 1.255 0.59 ;
      RECT  1.14 0.59 1.255 1.11 ;
      RECT  0.35 1.11 2.05 1.225 ;
      RECT  0.35 1.225 3.72 1.29 ;
      RECT  1.95 1.29 3.72 1.315 ;
      RECT  1.42 1.29 1.54 1.49 ;
      RECT  1.95 1.315 2.125 1.49 ;
      RECT  2.525 1.315 2.65 1.49 ;
      RECT  3.045 1.315 3.165 1.49 ;
      RECT  3.55 1.315 3.72 1.49 ;
    END
    ANTENNADIFFAREA 0.859 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.305 0.23 1.54 0.35 ;
      RECT  1.42 0.35 1.54 0.475 ;
      RECT  1.42 0.475 3.72 0.59 ;
      RECT  3.6 0.36 3.72 0.475 ;
  END
END SEN_ND2_T_5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_6
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_6
  CLASS CORE ;
  FOREIGN SEN_ND2_T_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 1.34 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3708 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 3.65 0.9 ;
      RECT  2.55 0.9 3.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5436 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.365 1.39 0.485 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.885 1.39 1.005 1.75 ;
      RECT  1.405 1.39 1.525 1.75 ;
      RECT  1.995 1.405 2.115 1.75 ;
      RECT  2.56 1.405 2.68 1.75 ;
      RECT  3.125 1.405 3.245 1.75 ;
      RECT  3.67 1.405 3.79 1.75 ;
      RECT  4.2 1.23 4.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  1.995 0.05 2.115 0.385 ;
      RECT  2.555 0.05 2.675 0.385 ;
      RECT  3.125 0.05 3.245 0.385 ;
      RECT  3.67 0.05 3.79 0.385 ;
      RECT  4.21 0.05 4.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.44 1.65 0.57 ;
      RECT  1.52 0.57 1.65 1.11 ;
      RECT  0.105 1.11 2.45 1.225 ;
      RECT  0.105 1.225 4.05 1.29 ;
      RECT  2.275 1.29 4.05 1.315 ;
      RECT  1.695 1.29 1.85 1.49 ;
      RECT  2.275 1.315 2.395 1.49 ;
      RECT  2.84 1.315 2.96 1.49 ;
      RECT  3.41 1.315 3.53 1.49 ;
      RECT  3.93 1.315 4.05 1.49 ;
    END
    ANTENNADIFFAREA 1.002 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.22 1.88 0.35 ;
      RECT  1.75 0.35 1.88 0.475 ;
      RECT  1.75 0.475 4.1 0.61 ;
  END
END SEN_ND2_T_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_T_8
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_T_8
  CLASS CORE ;
  FOREIGN SEN_ND2_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.685 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 0.9 ;
      RECT  3.35 0.9 4.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7248 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.61 1.39 0.73 1.75 ;
      RECT  1.13 1.39 1.25 1.75 ;
      RECT  1.66 1.39 1.78 1.75 ;
      RECT  2.2 1.39 2.32 1.75 ;
      RECT  2.735 1.415 2.855 1.75 ;
      RECT  3.255 1.415 3.375 1.75 ;
      RECT  3.775 1.415 3.895 1.75 ;
      RECT  4.31 1.415 4.43 1.75 ;
      RECT  4.85 1.415 4.97 1.75 ;
      RECT  5.39 1.21 5.51 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  2.475 0.05 2.595 0.38 ;
      RECT  2.995 0.05 3.115 0.38 ;
      RECT  3.515 0.05 3.635 0.38 ;
      RECT  4.055 0.05 4.175 0.38 ;
      RECT  4.59 0.05 4.71 0.38 ;
      RECT  5.11 0.05 5.23 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.3 0.46 2.06 0.6 ;
      RECT  1.89 0.6 2.06 1.11 ;
      RECT  0.35 1.11 3.25 1.21 ;
      RECT  0.35 1.21 5.25 1.29 ;
      RECT  2.95 1.29 5.25 1.325 ;
      RECT  2.475 1.29 2.595 1.49 ;
      RECT  2.95 1.325 3.115 1.49 ;
      RECT  3.515 1.325 3.65 1.49 ;
      RECT  4.035 1.325 4.155 1.49 ;
      RECT  4.55 1.325 4.71 1.49 ;
      RECT  5.11 1.325 5.25 1.49 ;
    END
    ANTENNADIFFAREA 1.264 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.09 0.22 2.345 0.36 ;
      RECT  0.09 0.36 0.21 0.445 ;
      RECT  2.175 0.36 2.345 0.47 ;
      RECT  2.175 0.47 5.54 0.62 ;
  END
END SEN_ND2_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_0P65
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_0P65
  CLASS CORE ;
  FOREIGN SEN_ND2_G_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.64 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0423 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0423 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.615 1.21 0.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.61 0.05 0.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.31 0.45 0.49 ;
      RECT  0.35 0.49 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.128 ;
  END X
END SEN_ND2_G_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_1
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_1
  CLASS CORE ;
  FOREIGN SEN_ND2_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.615 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      RECT  0.605 1.41 0.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.61 0.05 0.73 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.31 0.45 0.49 ;
      RECT  0.35 0.49 0.45 1.29 ;
    END
    ANTENNADIFFAREA 0.197 ;
  END X
END SEN_ND2_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_2
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_2
  CLASS CORE ;
  FOREIGN SEN_ND2_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.64 1.39 0.76 1.75 ;
      RECT  1.2 1.21 1.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.92 0.05 1.045 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.465 0.65 0.585 ;
      RECT  0.55 0.585 0.65 1.11 ;
      RECT  0.34 1.11 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.392 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.18 0.2 0.255 ;
      RECT  0.08 0.255 0.83 0.375 ;
      RECT  0.74 0.375 0.83 0.48 ;
      RECT  0.74 0.48 1.3 0.59 ;
      RECT  1.18 0.37 1.3 0.48 ;
  END
END SEN_ND2_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_3
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_3
  CLASS CORE ;
  FOREIGN SEN_ND2_G_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  1.105 1.415 1.225 1.75 ;
      RECT  1.615 1.41 1.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.12 0.05 1.225 0.385 ;
      RECT  1.615 0.05 1.745 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.34 0.185 0.44 ;
      RECT  0.065 0.44 0.85 0.56 ;
      RECT  0.75 0.56 0.85 1.21 ;
      RECT  0.275 1.21 1.535 1.325 ;
    END
    ANTENNADIFFAREA 0.533 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 0.23 1.03 0.35 ;
      RECT  0.94 0.35 1.03 0.48 ;
      RECT  0.94 0.48 1.535 0.6 ;
  END
END SEN_ND2_G_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2_G_4
#      Description : "2-Input NAND"
#      Equation    : X=!(A1&A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2_G_4
  CLASS CORE ;
  FOREIGN SEN_ND2_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.595 1.39 0.715 1.75 ;
      RECT  1.115 1.39 1.235 1.75 ;
      RECT  1.635 1.39 1.755 1.75 ;
      RECT  2.175 1.21 2.295 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.375 0.05 1.495 0.4 ;
      RECT  1.895 0.05 2.015 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.285 0.44 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.11 ;
      RECT  0.34 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.23 1.26 0.35 ;
      RECT  0.075 0.35 0.195 0.455 ;
      RECT  1.16 0.35 1.26 0.49 ;
      RECT  1.16 0.49 2.325 0.61 ;
  END
END SEN_ND2_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_1
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_1
  CLASS CORE ;
  FOREIGN SEN_ND2B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.67 0.255 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0516 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.525 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.41 0.49 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.935 1.22 1.055 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.37 0.05 0.5 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.31 1.06 1.035 ;
      RECT  0.74 1.035 1.06 1.125 ;
      RECT  0.74 1.125 0.83 1.41 ;
      RECT  0.62 1.41 0.83 1.53 ;
    END
    ANTENNADIFFAREA 0.209 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.34 0.185 0.47 ;
      RECT  0.065 0.47 0.85 0.56 ;
      RECT  0.745 0.56 0.85 0.925 ;
      RECT  0.345 0.56 0.435 1.21 ;
      RECT  0.065 1.21 0.435 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
  END
END SEN_ND2B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_2
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_2
  CLASS CORE ;
  FOREIGN SEN_ND2B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1032 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.585 1.21 0.705 1.75 ;
      RECT  1.205 1.41 1.335 1.75 ;
      RECT  1.81 1.21 1.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.58 0.05 0.705 0.36 ;
      RECT  1.545 0.05 1.675 0.36 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.005 0.57 1.205 0.68 ;
      RECT  1.115 0.68 1.205 0.69 ;
      RECT  1.115 0.69 1.25 1.11 ;
      RECT  0.845 1.11 1.66 1.29 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.795 0.34 1.41 0.43 ;
      RECT  1.29 0.43 1.41 0.45 ;
      RECT  0.77 0.43 0.89 0.635 ;
      RECT  1.29 0.45 1.93 0.54 ;
      RECT  1.81 0.32 1.93 0.45 ;
      RECT  0.34 0.36 0.445 0.78 ;
      RECT  0.34 0.78 1.0 0.9 ;
      RECT  0.34 0.9 0.445 1.36 ;
  END
END SEN_ND2B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_3
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_3
  CLASS CORE ;
  FOREIGN SEN_ND2B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.45 0.925 ;
      RECT  0.15 0.925 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1548 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.8 1.45 1.09 ;
      RECT  0.75 1.09 0.85 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.36 1.44 1.49 1.75 ;
      RECT  1.88 1.44 2.01 1.75 ;
      RECT  2.405 1.21 2.525 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.34 0.05 1.51 0.32 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  0.84 0.05 0.97 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.86 0.51 2.53 0.69 ;
      RECT  2.15 0.69 2.265 1.23 ;
      RECT  1.075 1.23 2.265 1.35 ;
    END
    ANTENNADIFFAREA 0.535 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.625 0.23 2.32 0.35 ;
      RECT  1.625 0.35 1.745 0.41 ;
      RECT  1.08 0.41 1.745 0.51 ;
      RECT  0.065 0.36 0.185 0.47 ;
      RECT  0.065 0.47 0.97 0.59 ;
      RECT  0.88 0.59 0.97 0.6 ;
      RECT  0.54 0.59 0.63 1.21 ;
      RECT  0.88 0.6 1.65 0.69 ;
      RECT  1.55 0.69 1.65 0.785 ;
      RECT  1.55 0.785 2.04 0.895 ;
      RECT  0.065 1.21 0.63 1.3 ;
      RECT  0.54 1.3 0.63 1.38 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.54 1.38 0.705 1.55 ;
  END
END SEN_ND2B_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_4
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_4
  CLASS CORE ;
  FOREIGN SEN_ND2B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.9 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2064 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.245 1.21 1.365 1.75 ;
      RECT  1.85 1.41 1.98 1.75 ;
      RECT  2.37 1.41 2.5 1.75 ;
      RECT  2.89 1.41 3.02 1.75 ;
      RECT  3.415 1.21 3.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.1 0.05 1.23 0.39 ;
      RECT  2.63 0.05 2.76 0.39 ;
      RECT  3.15 0.05 3.28 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 2.26 0.69 ;
      RECT  2.14 0.69 2.26 1.11 ;
      RECT  1.55 1.11 3.26 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.335 0.2 2.495 0.32 ;
      RECT  1.335 0.32 1.455 0.395 ;
      RECT  2.375 0.32 2.495 0.48 ;
      RECT  2.375 0.48 3.535 0.6 ;
      RECT  3.415 0.38 3.535 0.48 ;
      RECT  0.3 0.48 1.12 0.58 ;
      RECT  1.0 0.58 1.12 0.785 ;
      RECT  1.0 0.785 2.04 0.895 ;
      RECT  1.0 0.895 1.12 1.21 ;
      RECT  0.3 1.21 1.12 1.32 ;
  END
END SEN_ND2B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_6
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_6
  CLASS CORE ;
  FOREIGN SEN_ND2B_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.11 0.9 ;
      RECT  0.35 0.9 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3105 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.65 0.89 ;
      RECT  4.55 0.89 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  1.49 1.11 1.61 1.75 ;
      RECT  2.13 1.41 2.26 1.75 ;
      RECT  2.65 1.41 2.78 1.75 ;
      RECT  3.17 1.41 3.3 1.75 ;
      RECT  3.69 1.41 3.82 1.75 ;
      RECT  4.21 1.41 4.34 1.75 ;
      RECT  4.755 1.21 4.875 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      RECT  3.43 0.05 3.56 0.39 ;
      RECT  3.95 0.05 4.08 0.39 ;
      RECT  4.47 0.05 4.6 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.835 0.51 3.06 0.69 ;
      RECT  2.93 0.69 3.06 1.11 ;
      RECT  1.75 1.11 4.45 1.18 ;
      RECT  1.75 1.18 4.62 1.29 ;
    END
    ANTENNADIFFAREA 1.008 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.615 0.24 3.295 0.36 ;
      RECT  1.615 0.36 1.735 0.46 ;
      RECT  3.175 0.36 3.295 0.48 ;
      RECT  3.175 0.48 4.855 0.59 ;
      RECT  4.735 0.37 4.855 0.48 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 1.325 0.59 ;
      RECT  1.2 0.59 1.325 0.78 ;
      RECT  1.2 0.78 2.82 0.9 ;
      RECT  1.2 0.9 1.325 1.21 ;
      RECT  0.065 1.21 1.325 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
  END
END SEN_ND2B_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1DG_8
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1DG_8
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.51 3.85 0.93 ;
      RECT  2.75 0.51 2.85 0.93 ;
      RECT  1.55 0.51 1.65 0.93 ;
      RECT  0.55 0.51 0.65 0.93 ;
      LAYER M2 ;
      RECT  0.51 0.55 3.89 0.65 ;
      LAYER V1 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.39 1.225 1.75 ;
      RECT  1.625 1.39 1.745 1.75 ;
      RECT  2.145 1.39 2.265 1.75 ;
      RECT  2.665 1.39 2.785 1.75 ;
      RECT  3.185 1.39 3.305 1.75 ;
      RECT  3.705 1.39 3.825 1.75 ;
      RECT  4.255 1.19 4.375 1.75 ;
      RECT  4.81 1.21 4.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  4.805 0.05 4.94 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.12 0.05 1.225 0.61 ;
      RECT  2.145 0.05 2.26 0.61 ;
      RECT  3.185 0.05 3.29 0.61 ;
      RECT  4.25 0.05 4.37 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.32 3.86 0.42 ;
      RECT  3.56 0.42 3.66 1.11 ;
      RECT  2.55 0.32 2.835 0.42 ;
      RECT  2.55 0.42 2.65 1.11 ;
      RECT  1.575 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.54 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.325 1.11 4.085 1.29 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.95 0.23 4.05 0.775 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  3.95 0.775 4.66 0.895 ;
      RECT  4.54 0.45 4.66 0.775 ;
      RECT  4.54 0.895 4.66 1.32 ;
  END
END SEN_ND2B_V1DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1_16
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1_16
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.15 0.71 10.05 0.915 ;
      RECT  9.15 0.915 9.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4944 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.51 8.05 0.955 ;
      RECT  6.75 0.51 6.85 0.955 ;
      RECT  5.75 0.51 5.85 0.95 ;
      RECT  4.75 0.51 4.85 0.955 ;
      RECT  3.75 0.51 3.85 0.955 ;
      RECT  2.75 0.51 2.85 0.95 ;
      RECT  1.55 0.51 1.65 0.955 ;
      RECT  0.55 0.51 0.65 0.955 ;
      LAYER M2 ;
      RECT  0.51 0.55 8.09 0.65 ;
      LAYER V1 ;
      RECT  7.95 0.55 8.05 0.65 ;
      RECT  6.75 0.55 6.85 0.65 ;
      RECT  5.75 0.55 5.85 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9888 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 10.8 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.39 1.225 1.75 ;
      RECT  1.625 1.39 1.745 1.75 ;
      RECT  2.145 1.39 2.265 1.75 ;
      RECT  2.665 1.39 2.785 1.75 ;
      RECT  3.185 1.415 3.305 1.75 ;
      RECT  3.68 1.48 3.85 1.75 ;
      RECT  4.2 1.48 4.37 1.75 ;
      RECT  4.72 1.48 4.89 1.75 ;
      RECT  5.275 1.39 5.395 1.75 ;
      RECT  5.805 1.39 5.925 1.75 ;
      RECT  6.325 1.39 6.445 1.75 ;
      RECT  6.845 1.39 6.965 1.75 ;
      RECT  7.365 1.39 7.485 1.75 ;
      RECT  7.885 1.39 8.005 1.75 ;
      RECT  8.42 1.19 8.54 1.75 ;
      RECT  8.96 1.415 9.08 1.75 ;
      RECT  9.48 1.415 9.6 1.75 ;
      RECT  10.0 1.415 10.12 1.75 ;
      RECT  10.54 1.21 10.66 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      RECT  8.96 0.05 9.08 0.385 ;
      RECT  9.48 0.05 9.6 0.385 ;
      RECT  10.0 0.05 10.12 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  10.54 0.05 10.66 0.59 ;
      RECT  1.12 0.05 1.225 0.61 ;
      RECT  2.145 0.05 2.26 0.61 ;
      RECT  3.185 0.05 3.29 0.61 ;
      RECT  4.225 0.05 4.345 0.61 ;
      RECT  5.3 0.05 5.405 0.61 ;
      RECT  6.34 0.05 6.445 0.61 ;
      RECT  7.365 0.05 7.48 0.61 ;
      RECT  8.42 0.05 8.54 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.32 8.03 0.42 ;
      RECT  7.75 0.42 7.85 1.11 ;
      RECT  6.795 0.32 7.05 0.42 ;
      RECT  6.95 0.42 7.05 1.06 ;
      RECT  5.755 0.32 6.05 0.42 ;
      RECT  5.95 0.42 6.05 1.04 ;
      RECT  4.695 0.32 5.03 0.42 ;
      RECT  4.94 0.42 5.03 1.04 ;
      RECT  4.94 1.04 6.05 1.06 ;
      RECT  4.94 1.06 7.05 1.075 ;
      RECT  3.56 0.32 3.85 0.42 ;
      RECT  3.56 0.42 3.65 1.04 ;
      RECT  2.55 0.32 2.835 0.42 ;
      RECT  2.55 0.42 2.65 1.04 ;
      RECT  2.55 1.04 3.65 1.06 ;
      RECT  1.575 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.06 ;
      RECT  1.75 1.06 3.65 1.075 ;
      RECT  1.75 1.075 7.05 1.11 ;
      RECT  0.54 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.3 1.11 8.265 1.29 ;
      RECT  3.395 1.29 5.185 1.39 ;
    END
    ANTENNADIFFAREA 2.528 ;
  END X
  OBS
      LAYER M1 ;
      RECT  8.675 0.475 10.43 0.6 ;
      RECT  8.675 0.6 8.845 0.71 ;
      RECT  7.57 0.14 8.32 0.23 ;
      RECT  7.57 0.23 7.66 0.71 ;
      RECT  8.15 0.23 8.32 0.71 ;
      RECT  6.55 0.14 7.25 0.23 ;
      RECT  6.55 0.23 6.65 0.71 ;
      RECT  7.15 0.23 7.25 0.71 ;
      RECT  5.55 0.14 6.25 0.23 ;
      RECT  5.55 0.23 5.65 0.71 ;
      RECT  6.15 0.23 6.25 0.71 ;
      RECT  4.455 0.14 5.21 0.23 ;
      RECT  4.455 0.23 4.56 0.71 ;
      RECT  5.12 0.23 5.21 0.71 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.945 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.915 ;
      RECT  0.94 0.71 1.45 0.915 ;
      RECT  1.95 0.71 2.45 0.915 ;
      RECT  2.95 0.71 3.47 0.915 ;
      RECT  3.945 0.71 4.56 0.915 ;
      RECT  5.12 0.71 5.65 0.915 ;
      RECT  6.15 0.71 6.65 0.915 ;
      RECT  7.15 0.71 7.66 0.915 ;
      RECT  8.15 0.71 8.845 0.915 ;
      RECT  8.675 0.915 8.845 1.195 ;
      RECT  8.675 1.195 10.43 1.325 ;
      LAYER M2 ;
      RECT  3.91 0.35 8.29 0.45 ;
      LAYER V1 ;
      RECT  3.95 0.35 4.05 0.45 ;
      RECT  5.55 0.35 5.65 0.45 ;
      RECT  6.55 0.35 6.65 0.45 ;
      RECT  7.15 0.35 7.25 0.45 ;
      RECT  8.15 0.35 8.25 0.45 ;
  END
END SEN_ND2B_V1_16
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1_6
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1_6
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 4.05 0.915 ;
      RECT  3.95 0.915 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1854 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 0.955 ;
      RECT  1.55 0.51 1.65 0.955 ;
      RECT  0.55 0.51 0.65 0.955 ;
      LAYER M2 ;
      RECT  0.51 0.55 2.89 0.65 ;
      LAYER V1 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3708 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.39 1.225 1.75 ;
      RECT  1.625 1.39 1.745 1.75 ;
      RECT  2.145 1.39 2.265 1.75 ;
      RECT  2.665 1.39 2.785 1.75 ;
      RECT  3.185 1.405 3.305 1.75 ;
      RECT  3.72 1.415 3.84 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  3.185 0.05 3.305 0.385 ;
      RECT  3.72 0.05 3.84 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.12 0.05 1.225 0.61 ;
      RECT  2.145 0.05 2.26 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.32 2.835 0.42 ;
      RECT  2.55 0.42 2.65 1.11 ;
      RECT  1.575 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.54 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.3 1.11 3.05 1.29 ;
    END
    ANTENNADIFFAREA 0.948 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.0 0.37 4.12 0.475 ;
      RECT  3.35 0.475 4.12 0.595 ;
      RECT  3.35 0.595 3.45 0.81 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.81 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.915 ;
      RECT  0.94 0.71 1.45 0.915 ;
      RECT  1.95 0.71 2.45 0.915 ;
      RECT  2.95 0.81 3.45 0.92 ;
      RECT  3.35 0.92 3.45 1.205 ;
      RECT  3.35 1.205 4.12 1.325 ;
      RECT  4.0 1.325 4.12 1.435 ;
  END
END SEN_ND2B_V1_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1_8
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1_8
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.25 0.915 ;
      RECT  5.15 0.915 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.51 3.85 0.955 ;
      RECT  2.75 0.51 2.85 0.955 ;
      RECT  1.55 0.51 1.65 0.955 ;
      RECT  0.55 0.51 0.65 0.955 ;
      LAYER M2 ;
      RECT  0.51 0.55 3.89 0.65 ;
      LAYER V1 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.39 1.225 1.75 ;
      RECT  1.625 1.39 1.745 1.75 ;
      RECT  2.145 1.39 2.265 1.75 ;
      RECT  2.665 1.39 2.785 1.75 ;
      RECT  3.185 1.39 3.305 1.75 ;
      RECT  3.705 1.39 3.825 1.75 ;
      RECT  4.255 1.19 4.375 1.75 ;
      RECT  4.81 1.415 4.93 1.75 ;
      RECT  5.36 1.21 5.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  4.81 0.05 4.93 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.36 0.05 5.48 0.59 ;
      RECT  1.12 0.05 1.225 0.61 ;
      RECT  2.145 0.05 2.26 0.61 ;
      RECT  3.185 0.05 3.29 0.61 ;
      RECT  4.255 0.05 4.375 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.32 3.86 0.42 ;
      RECT  3.56 0.42 3.66 1.11 ;
      RECT  2.55 0.32 2.835 0.42 ;
      RECT  2.55 0.42 2.65 1.11 ;
      RECT  1.575 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.54 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.3 1.11 4.085 1.29 ;
    END
    ANTENNADIFFAREA 1.264 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.54 0.475 5.25 0.595 ;
      RECT  4.54 0.595 4.66 0.805 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.95 0.23 4.05 0.805 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.915 ;
      RECT  0.94 0.71 1.45 0.915 ;
      RECT  1.95 0.71 2.45 0.915 ;
      RECT  2.95 0.71 3.47 0.915 ;
      RECT  3.95 0.805 4.66 0.925 ;
      RECT  4.54 0.925 4.66 1.205 ;
      RECT  4.54 1.205 5.25 1.325 ;
  END
END SEN_ND2B_V1_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_12
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_12
  CLASS CORE ;
  FOREIGN SEN_ND2B_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.71 7.65 0.915 ;
      RECT  7.55 0.915 7.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3708 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.14 6.25 0.23 ;
      RECT  5.55 0.23 5.65 0.71 ;
      RECT  6.15 0.23 6.25 0.71 ;
      RECT  4.545 0.14 5.25 0.23 ;
      RECT  4.545 0.23 4.65 0.71 ;
      RECT  5.15 0.23 5.25 0.71 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.95 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.915 ;
      RECT  0.94 0.71 1.45 0.915 ;
      RECT  1.95 0.71 2.45 0.915 ;
      RECT  2.95 0.71 3.47 0.915 ;
      RECT  3.95 0.71 4.65 0.915 ;
      RECT  5.15 0.71 5.65 0.915 ;
      RECT  6.15 0.71 6.45 0.915 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7416 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.39 1.225 1.75 ;
      RECT  1.625 1.39 1.745 1.75 ;
      RECT  2.145 1.39 2.265 1.75 ;
      RECT  2.665 1.39 2.785 1.75 ;
      RECT  3.185 1.39 3.305 1.75 ;
      RECT  3.705 1.39 3.825 1.75 ;
      RECT  4.255 1.39 4.375 1.75 ;
      RECT  4.805 1.39 4.925 1.75 ;
      RECT  5.35 1.39 5.47 1.75 ;
      RECT  5.87 1.39 5.99 1.75 ;
      RECT  6.415 1.19 6.535 1.75 ;
      RECT  6.96 1.415 7.08 1.75 ;
      RECT  7.48 1.415 7.6 1.75 ;
      RECT  8.015 1.21 8.135 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  6.96 0.05 7.08 0.385 ;
      RECT  7.48 0.05 7.6 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  8.015 0.05 8.135 0.59 ;
      RECT  1.12 0.05 1.225 0.61 ;
      RECT  2.145 0.05 2.26 0.61 ;
      RECT  3.185 0.05 3.29 0.61 ;
      RECT  4.255 0.05 4.375 0.61 ;
      RECT  5.34 0.05 5.46 0.61 ;
      RECT  6.415 0.05 6.535 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.32 6.04 0.42 ;
      RECT  5.75 0.42 5.85 1.11 ;
      RECT  4.755 0.32 5.05 0.42 ;
      RECT  4.95 0.42 5.05 1.11 ;
      RECT  3.56 0.32 3.86 0.42 ;
      RECT  3.56 0.42 3.66 1.035 ;
      RECT  2.55 0.32 2.835 0.42 ;
      RECT  2.55 0.42 2.65 1.035 ;
      RECT  2.55 1.035 3.66 1.11 ;
      RECT  1.575 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.54 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.325 1.11 6.25 1.29 ;
    END
    ANTENNADIFFAREA 1.896 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.7 0.475 7.91 0.595 ;
      RECT  6.7 0.595 6.85 1.205 ;
      RECT  6.7 1.205 7.91 1.325 ;
      RECT  2.75 0.51 2.85 0.945 ;
      RECT  3.75 0.51 3.85 0.945 ;
      RECT  0.55 0.51 0.65 0.955 ;
      RECT  1.55 0.51 1.65 0.955 ;
      RECT  4.75 0.51 4.85 0.955 ;
      RECT  5.95 0.51 6.05 0.955 ;
      LAYER M2 ;
      RECT  0.51 0.55 6.89 0.65 ;
      LAYER V1 ;
      RECT  0.55 0.55 0.65 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  5.95 0.55 6.05 0.65 ;
      RECT  6.75 0.55 6.85 0.65 ;
  END
END SEN_ND2B_12
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_16
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_16
  CLASS CORE ;
  FOREIGN SEN_ND2B_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.15 0.71 10.05 0.915 ;
      RECT  9.15 0.915 9.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4944 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.57 0.14 8.25 0.23 ;
      RECT  7.57 0.23 7.66 0.71 ;
      RECT  8.15 0.23 8.25 0.71 ;
      RECT  6.55 0.14 7.25 0.23 ;
      RECT  6.55 0.23 6.65 0.71 ;
      RECT  7.15 0.23 7.25 0.71 ;
      RECT  5.55 0.14 6.25 0.23 ;
      RECT  5.55 0.23 5.65 0.71 ;
      RECT  6.15 0.23 6.25 0.71 ;
      RECT  4.455 0.14 5.21 0.23 ;
      RECT  4.455 0.23 4.56 0.71 ;
      RECT  5.12 0.23 5.21 0.71 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.945 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.915 ;
      RECT  0.94 0.71 1.45 0.915 ;
      RECT  1.95 0.71 2.45 0.915 ;
      RECT  2.95 0.71 3.47 0.915 ;
      RECT  3.945 0.71 4.56 0.915 ;
      RECT  5.12 0.71 5.65 0.915 ;
      RECT  6.15 0.71 6.65 0.915 ;
      RECT  7.15 0.71 7.66 0.915 ;
      RECT  8.15 0.71 8.45 0.915 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9888 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 10.8 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.39 1.225 1.75 ;
      RECT  1.625 1.39 1.745 1.75 ;
      RECT  2.145 1.39 2.265 1.75 ;
      RECT  2.665 1.39 2.785 1.75 ;
      RECT  3.185 1.415 3.305 1.75 ;
      RECT  3.68 1.48 3.85 1.75 ;
      RECT  4.2 1.48 4.37 1.75 ;
      RECT  4.72 1.48 4.89 1.75 ;
      RECT  5.285 1.415 5.405 1.75 ;
      RECT  5.805 1.39 5.925 1.75 ;
      RECT  6.325 1.39 6.445 1.75 ;
      RECT  6.845 1.39 6.965 1.75 ;
      RECT  7.365 1.39 7.485 1.75 ;
      RECT  7.885 1.39 8.005 1.75 ;
      RECT  8.44 1.19 8.56 1.75 ;
      RECT  9.0 1.415 9.12 1.75 ;
      RECT  9.52 1.415 9.64 1.75 ;
      RECT  10.04 1.415 10.16 1.75 ;
      RECT  10.58 1.21 10.7 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      RECT  9.0 0.05 9.12 0.385 ;
      RECT  9.52 0.05 9.64 0.385 ;
      RECT  10.04 0.05 10.16 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  10.58 0.05 10.7 0.59 ;
      RECT  1.12 0.05 1.225 0.61 ;
      RECT  2.145 0.05 2.26 0.61 ;
      RECT  3.185 0.05 3.29 0.61 ;
      RECT  4.225 0.05 4.345 0.61 ;
      RECT  5.3 0.05 5.405 0.61 ;
      RECT  6.34 0.05 6.445 0.61 ;
      RECT  8.44 0.05 8.56 0.61 ;
      RECT  7.365 0.05 7.48 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.32 8.055 0.42 ;
      RECT  7.75 0.42 7.85 1.11 ;
      RECT  6.795 0.32 7.05 0.42 ;
      RECT  6.95 0.42 7.05 1.06 ;
      RECT  5.755 0.32 6.05 0.42 ;
      RECT  5.95 0.42 6.05 1.04 ;
      RECT  4.695 0.32 5.03 0.42 ;
      RECT  4.94 0.42 5.03 1.04 ;
      RECT  4.94 1.04 6.05 1.06 ;
      RECT  4.94 1.06 7.05 1.075 ;
      RECT  3.56 0.32 3.855 0.42 ;
      RECT  3.56 0.42 3.65 1.04 ;
      RECT  2.55 0.32 2.835 0.42 ;
      RECT  2.55 0.42 2.65 1.04 ;
      RECT  2.55 1.04 3.65 1.06 ;
      RECT  1.575 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.06 ;
      RECT  1.75 1.06 3.65 1.075 ;
      RECT  1.75 1.075 7.05 1.11 ;
      RECT  0.54 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.325 1.11 8.29 1.29 ;
      RECT  3.395 1.29 5.195 1.39 ;
    END
    ANTENNADIFFAREA 2.538 ;
  END X
  OBS
      LAYER M1 ;
      RECT  8.74 0.475 10.47 0.6 ;
      RECT  8.74 0.6 8.91 1.195 ;
      RECT  8.74 1.195 10.47 1.325 ;
      RECT  2.75 0.51 2.85 0.95 ;
      RECT  5.75 0.51 5.85 0.95 ;
      RECT  0.55 0.51 0.65 0.955 ;
      RECT  3.75 0.51 3.85 0.955 ;
      RECT  4.75 0.51 4.85 0.955 ;
      RECT  6.75 0.51 6.85 0.955 ;
      RECT  7.95 0.51 8.05 0.955 ;
      RECT  1.55 0.51 1.65 0.995 ;
      LAYER M2 ;
      RECT  0.51 0.55 8.89 0.65 ;
      LAYER V1 ;
      RECT  0.55 0.55 0.65 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  5.75 0.55 5.85 0.65 ;
      RECT  6.75 0.55 6.85 0.65 ;
      RECT  7.95 0.55 8.05 0.65 ;
      RECT  8.75 0.55 8.85 0.65 ;
  END
END SEN_ND2B_16
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_8
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_8
  CLASS CORE ;
  FOREIGN SEN_ND2B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.25 0.915 ;
      RECT  5.15 0.915 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.38 0.14 4.05 0.23 ;
      RECT  3.38 0.23 3.47 0.71 ;
      RECT  3.95 0.23 4.05 0.71 ;
      RECT  2.35 0.14 3.05 0.23 ;
      RECT  2.35 0.23 2.45 0.71 ;
      RECT  2.95 0.23 3.05 0.71 ;
      RECT  1.35 0.14 2.05 0.23 ;
      RECT  1.35 0.23 1.45 0.71 ;
      RECT  1.95 0.23 2.05 0.71 ;
      RECT  0.35 0.14 1.03 0.23 ;
      RECT  0.35 0.23 0.45 0.71 ;
      RECT  0.94 0.23 1.03 0.71 ;
      RECT  0.15 0.71 0.45 0.915 ;
      RECT  0.94 0.71 1.45 0.915 ;
      RECT  1.95 0.71 2.45 0.915 ;
      RECT  2.95 0.71 3.47 0.915 ;
      RECT  3.95 0.71 4.25 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.39 1.225 1.75 ;
      RECT  1.625 1.39 1.745 1.75 ;
      RECT  2.145 1.39 2.265 1.75 ;
      RECT  2.665 1.39 2.785 1.75 ;
      RECT  3.185 1.39 3.305 1.75 ;
      RECT  3.705 1.39 3.825 1.75 ;
      RECT  4.25 1.19 4.37 1.75 ;
      RECT  4.81 1.415 4.93 1.75 ;
      RECT  5.36 1.21 5.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  4.81 0.05 4.93 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.36 0.05 5.48 0.59 ;
      RECT  1.12 0.05 1.225 0.61 ;
      RECT  2.145 0.05 2.26 0.61 ;
      RECT  3.185 0.05 3.29 0.61 ;
      RECT  4.25 0.05 4.37 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.32 3.86 0.42 ;
      RECT  3.56 0.42 3.66 1.11 ;
      RECT  2.55 0.32 2.835 0.42 ;
      RECT  2.55 0.42 2.65 1.11 ;
      RECT  1.575 0.32 1.85 0.42 ;
      RECT  1.75 0.42 1.85 1.11 ;
      RECT  0.54 0.32 0.85 0.42 ;
      RECT  0.75 0.42 0.85 1.11 ;
      RECT  0.325 1.11 4.085 1.29 ;
    END
    ANTENNADIFFAREA 1.264 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.54 0.475 5.25 0.595 ;
      RECT  4.54 0.595 4.66 1.205 ;
      RECT  4.54 1.205 5.25 1.325 ;
      RECT  0.55 0.51 0.65 0.955 ;
      RECT  1.55 0.51 1.65 0.955 ;
      RECT  2.75 0.51 2.85 0.955 ;
      RECT  3.75 0.51 3.85 0.955 ;
      LAYER M2 ;
      RECT  0.51 0.55 4.69 0.65 ;
      LAYER V1 ;
      RECT  0.55 0.55 0.65 0.65 ;
      RECT  1.55 0.55 1.65 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  4.55 0.55 4.65 0.65 ;
  END
END SEN_ND2B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1DG_1
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1DG_1
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.63 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.66 1.39 0.79 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.655 0.05 0.785 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.31 0.45 0.49 ;
      RECT  0.35 0.49 0.45 1.29 ;
    END
    ANTENNADIFFAREA 0.197 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.98 0.19 1.1 0.5 ;
      RECT  0.55 0.5 1.1 0.595 ;
      RECT  0.55 0.595 0.65 1.21 ;
      RECT  0.55 1.21 1.1 1.3 ;
      RECT  0.98 1.3 1.1 1.61 ;
  END
END SEN_ND2B_V1DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1DG_2
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1DG_2
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.19 1.225 1.75 ;
      RECT  1.605 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.605 0.05 1.74 0.39 ;
      RECT  0.845 0.05 0.975 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.47 0.45 1.11 ;
      RECT  0.34 1.11 0.965 1.29 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.24 0.73 0.36 ;
      RECT  0.065 0.36 0.185 0.42 ;
      RECT  0.64 0.36 0.73 0.505 ;
      RECT  0.64 0.505 1.265 0.625 ;
      RECT  1.355 0.19 1.46 0.785 ;
      RECT  0.82 0.785 1.46 0.895 ;
      RECT  1.355 0.895 1.46 1.51 ;
  END
END SEN_ND2B_V1DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1DG_4
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1DG_4
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.185 1.75 ;
      RECT  0.0 1.75 2.8 1.85 ;
      RECT  0.575 1.39 0.695 1.75 ;
      RECT  1.095 1.39 1.215 1.75 ;
      RECT  1.615 1.39 1.735 1.75 ;
      RECT  2.14 1.19 2.255 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      RECT  1.355 0.05 1.475 0.385 ;
      RECT  1.875 0.05 1.995 0.385 ;
      RECT  2.605 0.05 2.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.265 0.44 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.11 ;
      RECT  0.35 1.11 2.05 1.29 ;
      RECT  0.35 1.29 0.45 1.315 ;
      RECT  0.315 1.315 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.225 1.24 0.345 ;
      RECT  0.055 0.345 0.175 0.42 ;
      RECT  1.14 0.345 1.24 0.485 ;
      RECT  1.14 0.485 2.255 0.605 ;
      RECT  2.135 0.605 2.255 0.68 ;
      RECT  2.345 0.19 2.46 0.785 ;
      RECT  1.475 0.785 2.46 0.895 ;
      RECT  2.37 0.895 2.46 1.24 ;
      RECT  2.37 1.24 2.565 1.36 ;
  END
END SEN_ND2B_V1DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_S_0P5
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_S_0P5
  CLASS CORE ;
  FOREIGN SEN_ND2B_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.71 0.255 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0216 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.475 0.505 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.94 1.44 1.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.33 0.05 0.45 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.205 1.05 1.26 ;
      RECT  0.75 1.26 1.05 1.31 ;
      RECT  0.63 1.31 1.05 1.35 ;
      RECT  0.63 1.35 0.85 1.49 ;
    END
    ANTENNADIFFAREA 0.106 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.185 0.19 0.505 ;
      RECT  0.07 0.505 0.45 0.595 ;
      RECT  0.36 0.595 0.45 1.08 ;
      RECT  0.36 1.08 0.855 1.17 ;
      RECT  0.745 0.915 0.855 1.08 ;
      RECT  0.36 1.17 0.45 1.26 ;
      RECT  0.07 1.26 0.45 1.38 ;
      RECT  0.07 1.38 0.19 1.625 ;
  END
END SEN_ND2B_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_S_1
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_S_1
  CLASS CORE ;
  FOREIGN SEN_ND2B_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.71 0.255 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0318 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.475 0.505 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.94 1.44 1.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.33 0.05 0.45 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.31 1.05 0.6 ;
      RECT  0.95 0.6 1.12 0.69 ;
      RECT  1.02 0.69 1.12 1.26 ;
      RECT  0.665 1.26 1.12 1.35 ;
      RECT  0.665 1.35 0.85 1.49 ;
    END
    ANTENNADIFFAREA 0.211 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.18 0.19 0.495 ;
      RECT  0.07 0.495 0.45 0.585 ;
      RECT  0.36 0.585 0.45 1.07 ;
      RECT  0.36 1.07 0.93 1.16 ;
      RECT  0.82 0.78 0.93 1.07 ;
      RECT  0.36 1.16 0.45 1.26 ;
      RECT  0.07 1.26 0.45 1.38 ;
      RECT  0.07 1.38 0.19 1.48 ;
  END
END SEN_ND2B_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_S_12
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_S_12
  CLASS CORE ;
  FOREIGN SEN_ND2B_S_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.25 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3264 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.71 8.05 0.89 ;
      RECT  7.95 0.89 8.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.625 1.24 0.745 1.75 ;
      RECT  1.155 1.235 1.275 1.75 ;
      RECT  1.675 1.21 1.795 1.75 ;
      RECT  2.195 1.415 2.315 1.75 ;
      RECT  2.715 1.415 2.835 1.75 ;
      RECT  3.235 1.415 3.355 1.75 ;
      RECT  3.755 1.415 3.875 1.75 ;
      RECT  4.275 1.415 4.395 1.75 ;
      RECT  4.795 1.415 4.915 1.75 ;
      RECT  5.35 1.415 5.47 1.75 ;
      RECT  5.87 1.415 5.99 1.75 ;
      RECT  6.39 1.415 6.51 1.75 ;
      RECT  6.91 1.415 7.03 1.75 ;
      RECT  7.43 1.415 7.55 1.75 ;
      RECT  7.975 1.21 8.09 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  5.09 0.05 5.21 0.35 ;
      RECT  5.61 0.05 5.73 0.35 ;
      RECT  6.13 0.05 6.25 0.35 ;
      RECT  6.65 0.05 6.77 0.35 ;
      RECT  7.17 0.05 7.29 0.35 ;
      RECT  7.69 0.05 7.81 0.35 ;
      RECT  0.865 0.05 0.985 0.37 ;
      RECT  1.425 0.05 1.545 0.37 ;
      RECT  0.24 0.05 0.36 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.94 0.51 4.66 0.69 ;
      RECT  3.95 0.69 4.66 0.72 ;
      RECT  4.41 0.72 4.66 1.08 ;
      RECT  3.95 1.08 5.25 1.11 ;
      RECT  1.94 1.11 7.85 1.29 ;
    END
    ANTENNADIFFAREA 2.038 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.21 0.16 5.0 0.24 ;
      RECT  1.635 0.24 5.0 0.37 ;
      RECT  4.75 0.37 5.0 0.44 ;
      RECT  4.75 0.44 8.12 0.56 ;
      RECT  4.75 0.56 6.535 0.61 ;
      RECT  4.75 0.61 5.47 0.65 ;
      RECT  0.535 0.46 1.56 0.58 ;
      RECT  1.43 0.58 1.56 0.78 ;
      RECT  1.43 0.78 3.805 0.81 ;
      RECT  1.43 0.81 4.265 0.905 ;
      RECT  1.43 0.905 1.56 1.005 ;
      RECT  0.34 1.005 1.56 1.135 ;
  END
END SEN_ND2B_S_12
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_S_2
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_S_2
  CLASS CORE ;
  FOREIGN SEN_ND2B_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0609 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.18 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.58 1.24 0.7 1.75 ;
      RECT  1.1 1.44 1.22 1.75 ;
      RECT  1.62 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.36 0.05 1.48 0.35 ;
      RECT  0.06 0.05 0.18 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.79 0.44 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.11 ;
      RECT  0.84 1.11 1.45 1.29 ;
      RECT  1.35 1.29 1.45 1.41 ;
      RECT  1.35 1.41 1.465 1.59 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.545 0.24 1.26 0.35 ;
      RECT  1.14 0.35 1.26 0.44 ;
      RECT  1.14 0.44 1.73 0.56 ;
      RECT  1.63 0.18 1.73 0.44 ;
      RECT  0.335 0.215 0.45 0.385 ;
      RECT  0.35 0.385 0.45 0.755 ;
      RECT  0.35 0.755 0.85 0.925 ;
      RECT  0.35 0.925 0.45 1.415 ;
      RECT  0.335 1.415 0.45 1.585 ;
  END
END SEN_ND2B_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_S_4
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_S_4
  CLASS CORE ;
  FOREIGN SEN_ND2B_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1098 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.095 1.21 0.215 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.635 1.22 0.755 1.75 ;
      RECT  0.895 1.21 1.015 1.75 ;
      RECT  1.415 1.38 1.535 1.75 ;
      RECT  1.935 1.38 2.055 1.75 ;
      RECT  2.455 1.38 2.575 1.75 ;
      RECT  2.99 1.21 3.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.61 0.05 0.78 0.32 ;
      RECT  2.195 0.05 2.315 0.35 ;
      RECT  2.715 0.05 2.835 0.35 ;
      RECT  0.085 0.05 0.225 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.85 0.69 ;
      RECT  1.75 0.69 1.85 1.11 ;
      RECT  1.15 1.11 2.85 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.87 0.24 2.055 0.36 ;
      RECT  1.95 0.36 2.055 0.44 ;
      RECT  1.95 0.44 3.095 0.56 ;
      RECT  2.975 0.34 3.095 0.44 ;
      RECT  0.32 0.41 0.73 0.515 ;
      RECT  0.64 0.515 0.73 0.785 ;
      RECT  0.64 0.785 1.585 0.895 ;
      RECT  0.64 0.895 0.73 1.01 ;
      RECT  0.34 1.01 0.73 1.13 ;
  END
END SEN_ND2B_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_S_8
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_S_8
  CLASS CORE ;
  FOREIGN SEN_ND2B_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2169 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.05 0.71 5.45 0.89 ;
      RECT  5.35 0.89 5.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.095 1.21 0.215 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.635 1.235 0.755 1.75 ;
      RECT  1.155 1.21 1.275 1.75 ;
      RECT  1.675 1.38 1.795 1.75 ;
      RECT  2.195 1.38 2.315 1.75 ;
      RECT  2.715 1.38 2.835 1.75 ;
      RECT  3.235 1.38 3.355 1.75 ;
      RECT  3.755 1.38 3.875 1.75 ;
      RECT  4.275 1.38 4.395 1.75 ;
      RECT  4.795 1.38 4.915 1.75 ;
      RECT  5.34 1.21 5.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.61 0.05 0.78 0.32 ;
      RECT  3.495 0.05 3.615 0.35 ;
      RECT  4.015 0.05 4.135 0.35 ;
      RECT  4.535 0.05 4.655 0.35 ;
      RECT  5.055 0.05 5.175 0.35 ;
      RECT  0.095 0.05 0.215 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.42 0.51 3.095 0.69 ;
      RECT  2.88 0.69 3.05 1.11 ;
      RECT  1.42 1.11 5.175 1.29 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.69 0.19 3.38 0.24 ;
      RECT  1.115 0.24 3.38 0.36 ;
      RECT  3.21 0.36 3.38 0.44 ;
      RECT  3.21 0.44 5.485 0.56 ;
      RECT  3.21 0.56 3.9 0.61 ;
      RECT  0.325 0.41 1.04 0.515 ;
      RECT  0.95 0.515 1.04 0.785 ;
      RECT  0.95 0.785 2.715 0.895 ;
      RECT  0.95 0.895 1.04 1.01 ;
      RECT  0.35 1.01 1.04 1.13 ;
  END
END SEN_ND2B_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1_1
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1_1
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.655 1.415 0.795 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.65 0.05 0.79 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.08 0.18 0.2 0.3 ;
      RECT  0.08 0.3 0.46 0.4 ;
      RECT  0.34 0.4 0.46 1.3 ;
    END
    ANTENNADIFFAREA 0.187 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.98 0.2 1.1 0.495 ;
      RECT  0.55 0.495 1.1 0.59 ;
      RECT  0.55 0.59 0.65 1.215 ;
      RECT  0.55 1.215 1.1 1.305 ;
      RECT  0.98 1.305 1.1 1.585 ;
  END
END SEN_ND2B_V1_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1_2
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1_2
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  1.105 1.155 1.225 1.75 ;
      RECT  1.615 1.21 1.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.61 0.05 1.74 0.39 ;
      RECT  0.835 0.05 0.975 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.45 0.45 1.11 ;
      RECT  0.34 1.11 0.99 1.29 ;
    END
    ANTENNADIFFAREA 0.316 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.185 0.705 0.305 ;
      RECT  0.065 0.305 0.185 0.41 ;
      RECT  0.585 0.305 0.705 0.5 ;
      RECT  0.585 0.5 1.25 0.62 ;
      RECT  1.355 0.36 1.46 0.81 ;
      RECT  0.79 0.81 1.46 0.92 ;
      RECT  1.355 0.92 1.46 1.32 ;
  END
END SEN_ND2B_V1_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1_3
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1_3
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0918 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.92 ;
      RECT  0.15 0.92 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1854 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.59 1.39 0.71 1.75 ;
      RECT  1.1 1.39 1.24 1.75 ;
      RECT  1.645 1.415 1.785 1.75 ;
      RECT  2.2 1.21 2.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.12 0.05 1.24 0.385 ;
      RECT  1.645 0.05 1.785 0.385 ;
      RECT  2.2 0.05 2.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.07 0.325 0.19 0.44 ;
      RECT  0.07 0.44 0.85 0.56 ;
      RECT  0.75 0.56 0.85 1.11 ;
      RECT  0.34 1.11 1.48 1.29 ;
    END
    ANTENNADIFFAREA 0.503 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.23 1.03 0.35 ;
      RECT  0.94 0.35 1.03 0.48 ;
      RECT  0.94 0.48 1.48 0.6 ;
      RECT  1.37 0.38 1.48 0.48 ;
      RECT  1.94 0.26 2.06 0.495 ;
      RECT  1.57 0.495 2.06 0.585 ;
      RECT  1.57 0.585 1.66 0.81 ;
      RECT  1.11 0.81 1.66 0.92 ;
      RECT  1.57 0.92 1.66 1.2 ;
      RECT  1.57 1.2 2.085 1.32 ;
  END
END SEN_ND2B_V1_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND2B_V1_4
#      Description : "2-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND2B_V1_4
  CLASS CORE ;
  FOREIGN SEN_ND2B_V1_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.92 ;
      RECT  2.55 0.92 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.92 ;
      RECT  0.15 0.92 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.6 1.415 0.72 1.75 ;
      RECT  1.12 1.415 1.24 1.75 ;
      RECT  1.64 1.415 1.76 1.75 ;
      RECT  2.16 1.16 2.28 1.75 ;
      RECT  2.415 1.415 2.555 1.75 ;
      RECT  2.96 1.21 3.08 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  1.38 0.05 1.5 0.385 ;
      RECT  1.9 0.05 2.02 0.385 ;
      RECT  2.425 0.05 2.545 0.385 ;
      RECT  2.96 0.05 3.08 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.29 0.44 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.11 ;
      RECT  0.34 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.632 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.23 1.265 0.35 ;
      RECT  0.08 0.35 0.2 0.455 ;
      RECT  1.165 0.35 1.265 0.48 ;
      RECT  1.165 0.48 2.28 0.6 ;
      RECT  2.16 0.375 2.28 0.48 ;
      RECT  2.37 0.48 2.855 0.6 ;
      RECT  2.37 0.6 2.46 0.81 ;
      RECT  1.435 0.81 2.46 0.92 ;
      RECT  2.37 0.92 2.46 1.2 ;
      RECT  2.37 1.2 2.855 1.32 ;
  END
END SEN_ND2B_V1_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_0P5
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_0P5
  CLASS CORE ;
  FOREIGN SEN_ND3_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.64 1.395 0.76 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.07 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.17 1.06 0.3 ;
      RECT  0.75 0.3 1.06 0.39 ;
      RECT  0.75 0.39 0.85 1.11 ;
      RECT  0.34 1.11 0.85 1.2 ;
      RECT  0.34 1.2 1.06 1.29 ;
      RECT  0.34 1.29 0.46 1.52 ;
      RECT  0.94 1.29 1.06 1.52 ;
    END
    ANTENNADIFFAREA 0.159 ;
  END X
END SEN_ND3_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_1
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_1
  CLASS CORE ;
  FOREIGN SEN_ND3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 0.71 ;
      RECT  0.35 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.64 1.395 0.76 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.07 0.05 0.2 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.17 1.06 0.3 ;
      RECT  0.75 0.3 1.06 0.39 ;
      RECT  0.75 0.39 0.85 1.11 ;
      RECT  0.35 1.11 0.85 1.18 ;
      RECT  0.35 1.18 1.06 1.29 ;
      RECT  0.94 1.29 1.06 1.49 ;
    END
    ANTENNADIFFAREA 0.304 ;
  END X
END SEN_ND3_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_2
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_2
  CLASS CORE ;
  FOREIGN SEN_ND3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.585 1.42 0.705 1.75 ;
      RECT  1.19 1.42 1.31 1.75 ;
      RECT  1.81 1.215 1.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.315 0.05 0.435 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.465 1.705 0.585 ;
      RECT  1.35 0.585 1.45 1.21 ;
      RECT  0.295 1.21 1.695 1.33 ;
    END
    ANTENNADIFFAREA 0.45 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.78 0.215 1.94 0.335 ;
      RECT  1.82 0.335 1.94 0.39 ;
      RECT  0.055 0.19 0.175 0.5 ;
      RECT  0.055 0.5 1.25 0.62 ;
  END
END SEN_ND3_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_3
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_3
  CLASS CORE ;
  FOREIGN SEN_ND3_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  1.105 1.415 1.225 1.75 ;
      RECT  1.625 1.415 1.745 1.75 ;
      RECT  2.145 1.415 2.265 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.585 0.05 0.705 0.38 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.405 0.37 2.525 0.47 ;
      RECT  1.75 0.47 2.525 0.59 ;
      RECT  1.75 0.59 1.85 1.205 ;
      RECT  0.295 1.205 2.535 1.325 ;
      RECT  2.415 1.325 2.535 1.43 ;
    END
    ANTENNADIFFAREA 0.75 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.08 0.22 2.32 0.34 ;
      RECT  0.295 0.47 1.54 0.59 ;
  END
END SEN_ND3_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_4
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_4
  CLASS CORE ;
  FOREIGN SEN_ND3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  1.105 1.415 1.225 1.75 ;
      RECT  1.625 1.415 1.745 1.75 ;
      RECT  2.25 1.415 2.37 1.75 ;
      RECT  2.87 1.415 2.99 1.75 ;
      RECT  3.41 1.21 3.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.325 0.05 0.445 0.385 ;
      RECT  0.845 0.05 0.965 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.44 3.28 0.56 ;
      RECT  2.55 0.56 2.65 1.11 ;
      RECT  2.55 1.11 3.25 1.205 ;
      RECT  0.3 1.205 3.25 1.325 ;
    END
    ANTENNADIFFAREA 0.9 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.31 0.23 3.51 0.35 ;
      RECT  3.39 0.35 3.51 0.45 ;
      RECT  0.065 0.38 0.185 0.49 ;
      RECT  0.065 0.49 2.32 0.61 ;
  END
END SEN_ND3_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_6
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_6
  CLASS CORE ;
  FOREIGN SEN_ND3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.51 5.05 0.71 ;
      RECT  4.02 0.71 5.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3852 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.85 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3852 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3852 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.585 1.43 0.705 1.75 ;
      RECT  1.105 1.43 1.225 1.75 ;
      RECT  1.625 1.43 1.745 1.75 ;
      RECT  2.145 1.43 2.265 1.75 ;
      RECT  2.675 1.43 2.795 1.75 ;
      RECT  3.325 1.43 3.445 1.75 ;
      RECT  3.97 1.43 4.09 1.75 ;
      RECT  4.49 1.43 4.61 1.75 ;
      RECT  5.01 1.21 5.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  0.325 0.05 0.445 0.37 ;
      RECT  0.845 0.05 0.965 0.37 ;
      RECT  1.365 0.05 1.485 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.41 4.855 0.46 ;
      RECT  3.68 0.46 4.855 0.58 ;
      RECT  3.75 0.58 3.88 1.11 ;
      RECT  3.75 1.11 4.9 1.21 ;
      RECT  0.295 1.21 4.9 1.34 ;
    END
    ANTENNADIFFAREA 1.35 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.9 0.22 3.595 0.23 ;
      RECT  1.83 0.23 5.13 0.32 ;
      RECT  1.83 0.32 4.64 0.35 ;
      RECT  5.01 0.32 5.13 0.4 ;
      RECT  0.065 0.36 0.185 0.46 ;
      RECT  0.065 0.46 3.37 0.58 ;
  END
END SEN_ND3_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_8
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_8
  CLASS CORE ;
  FOREIGN SEN_ND3_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.055 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5136 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.51 4.65 0.71 ;
      RECT  2.95 0.71 4.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5136 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.85 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5136 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 6.8 1.85 ;
      RECT  0.65 1.415 0.77 1.75 ;
      RECT  1.22 1.41 1.34 1.75 ;
      RECT  1.74 1.41 1.86 1.75 ;
      RECT  2.26 1.41 2.38 1.75 ;
      RECT  2.78 1.41 2.9 1.75 ;
      RECT  3.3 1.41 3.42 1.75 ;
      RECT  3.85 1.41 3.97 1.75 ;
      RECT  4.44 1.41 4.56 1.75 ;
      RECT  5.005 1.41 5.125 1.75 ;
      RECT  5.53 1.41 5.65 1.75 ;
      RECT  6.05 1.41 6.17 1.75 ;
      RECT  6.59 1.21 6.71 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      RECT  1.4 0.05 1.52 0.36 ;
      RECT  1.92 0.05 2.04 0.36 ;
      RECT  0.36 0.05 0.48 0.365 ;
      RECT  0.88 0.05 1.0 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.745 0.475 6.5 0.595 ;
      RECT  4.745 0.595 4.9 1.11 ;
      RECT  0.95 1.11 6.455 1.225 ;
      RECT  0.34 1.225 6.455 1.29 ;
      RECT  0.34 1.29 1.08 1.325 ;
      RECT  0.34 1.325 0.46 1.5 ;
    END
    ANTENNADIFFAREA 1.8 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.975 0.17 4.655 0.19 ;
      RECT  2.935 0.19 5.695 0.22 ;
      RECT  2.39 0.22 6.735 0.34 ;
      RECT  0.1 0.35 0.22 0.455 ;
      RECT  0.1 0.455 4.43 0.575 ;
      RECT  1.15 0.575 3.365 0.585 ;
      RECT  2.155 0.585 3.365 0.59 ;
      RECT  2.155 0.59 2.845 0.605 ;
  END
END SEN_ND3_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_S_0P5
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_S_0P5
  CLASS CORE ;
  FOREIGN SEN_ND3_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.5 0.92 0.89 ;
      RECT  0.82 0.89 0.92 1.265 ;
      RECT  0.625 1.265 0.92 1.365 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.175 1.75 ;
      RECT  0.0 1.75 1.0 1.85 ;
      RECT  0.55 1.48 0.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      RECT  0.785 0.05 0.915 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.17 0.175 0.31 ;
      RECT  0.065 0.31 0.45 0.49 ;
      RECT  0.35 0.49 0.45 1.0 ;
      RECT  0.35 1.0 0.73 1.1 ;
      RECT  0.63 1.1 0.73 1.175 ;
      RECT  0.35 1.1 0.46 1.475 ;
      RECT  0.265 1.475 0.46 1.575 ;
    END
    ANTENNADIFFAREA 0.156 ;
  END X
END SEN_ND3_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_S_1
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_S_1
  CLASS CORE ;
  FOREIGN SEN_ND3_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0456 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.51 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0456 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.91 ;
      RECT  0.75 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0456 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.64 1.4 0.76 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.94 0.05 1.06 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.07 0.17 0.19 0.29 ;
      RECT  0.07 0.29 0.45 0.39 ;
      RECT  0.35 0.39 0.45 1.21 ;
      RECT  0.35 1.21 1.06 1.31 ;
      RECT  0.94 1.31 1.06 1.555 ;
      RECT  0.35 1.31 0.45 1.575 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
END SEN_ND3_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_S_12
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_S_12
  CLASS CORE ;
  FOREIGN SEN_ND3_S_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.71 6.45 0.91 ;
      RECT  5.275 0.91 6.85 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5472 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 4.85 0.91 ;
      RECT  2.75 0.91 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5472 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.945 0.71 1.05 0.91 ;
      RECT  0.35 0.91 2.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5472 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.435 0.465 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  0.835 1.43 0.985 1.75 ;
      RECT  1.355 1.43 1.505 1.75 ;
      RECT  1.875 1.43 2.025 1.75 ;
      RECT  2.4 1.43 2.55 1.75 ;
      RECT  2.915 1.43 3.065 1.75 ;
      RECT  3.435 1.43 3.585 1.75 ;
      RECT  3.955 1.43 4.105 1.75 ;
      RECT  4.475 1.44 4.625 1.75 ;
      RECT  4.995 1.44 5.145 1.75 ;
      RECT  5.515 1.43 5.665 1.75 ;
      RECT  6.035 1.43 6.185 1.75 ;
      RECT  6.555 1.43 6.705 1.75 ;
      RECT  7.12 1.21 7.24 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  0.575 0.05 0.725 0.38 ;
      RECT  1.1 0.05 1.24 0.38 ;
      RECT  1.615 0.05 1.765 0.38 ;
      RECT  2.14 0.05 2.29 0.38 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.09 0.31 7.25 0.48 ;
      RECT  4.94 0.48 7.25 0.59 ;
      RECT  4.94 0.59 6.25 0.69 ;
      RECT  4.94 0.69 5.17 1.2 ;
      RECT  4.94 1.2 5.45 1.21 ;
      RECT  2.125 1.21 5.45 1.225 ;
      RECT  2.125 1.225 7.005 1.23 ;
      RECT  0.07 1.23 7.005 1.34 ;
      RECT  0.07 1.34 0.19 1.465 ;
    END
    ANTENNADIFFAREA 1.636 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.115 0.17 5.435 0.2 ;
      RECT  3.67 0.2 5.98 0.26 ;
      RECT  2.605 0.26 6.485 0.27 ;
      RECT  2.605 0.27 7.0 0.37 ;
      RECT  0.285 0.5 4.66 0.61 ;
      RECT  1.33 0.61 3.64 0.67 ;
      RECT  1.775 0.67 3.095 0.7 ;
  END
END SEN_ND3_S_12
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_S_2
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_S_2
  CLASS CORE ;
  FOREIGN SEN_ND3_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.91 ;
      RECT  0.55 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.705 1.85 0.91 ;
      RECT  1.55 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.58 1.43 0.72 1.75 ;
      RECT  1.185 1.415 1.335 1.75 ;
      RECT  1.815 1.37 1.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.555 0.05 1.675 0.405 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.345 0.475 0.45 1.23 ;
      RECT  0.345 1.23 1.675 1.32 ;
      RECT  0.86 1.32 1.05 1.57 ;
      RECT  1.55 1.32 1.675 1.57 ;
      RECT  0.345 1.32 0.45 1.575 ;
    END
    ANTENNADIFFAREA 0.264 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.235 1.28 0.355 ;
      RECT  0.08 0.355 0.18 0.465 ;
      RECT  1.825 0.375 1.925 0.505 ;
      RECT  0.8 0.505 1.925 0.615 ;
  END
END SEN_ND3_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_S_4
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_S_4
  CLASS CORE ;
  FOREIGN SEN_ND3_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  2.15 0.91 2.65 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1824 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 0.91 ;
      RECT  1.15 0.91 1.85 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1824 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.945 0.71 1.05 0.91 ;
      RECT  0.55 0.91 1.05 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1824 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.56 1.435 0.68 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.08 1.435 1.2 1.75 ;
      RECT  1.6 1.435 1.72 1.75 ;
      RECT  2.12 1.435 2.24 1.75 ;
      RECT  2.72 1.23 2.84 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.81 0.05 0.95 0.43 ;
      RECT  0.275 0.05 0.4 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.64 0.32 2.76 0.495 ;
      RECT  1.945 0.495 2.76 0.595 ;
      RECT  1.945 0.595 2.05 1.235 ;
      RECT  0.3 1.235 2.53 1.345 ;
      RECT  0.3 1.345 0.45 1.495 ;
    END
    ANTENNADIFFAREA 0.588 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.29 0.285 2.55 0.385 ;
      RECT  0.51 0.52 1.77 0.62 ;
  END
END SEN_ND3_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_S_8
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_S_8
  CLASS CORE ;
  FOREIGN SEN_ND3_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 4.85 0.91 ;
      RECT  3.81 0.91 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.05 0.91 ;
      RECT  1.95 0.91 3.05 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.71 0.85 0.91 ;
      RECT  0.35 0.91 1.45 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3648 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.09 1.21 0.21 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.61 1.44 0.73 1.75 ;
      RECT  1.13 1.44 1.25 1.75 ;
      RECT  1.65 1.44 1.77 1.75 ;
      RECT  2.17 1.44 2.29 1.75 ;
      RECT  2.69 1.44 2.81 1.75 ;
      RECT  3.3 1.44 3.42 1.75 ;
      RECT  3.915 1.44 4.035 1.75 ;
      RECT  4.435 1.44 4.555 1.75 ;
      RECT  4.97 1.21 5.09 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  0.35 0.05 0.47 0.405 ;
      RECT  0.87 0.05 0.99 0.405 ;
      RECT  1.39 0.05 1.51 0.405 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.485 4.875 0.605 ;
      RECT  3.55 0.605 4.65 0.69 ;
      RECT  3.55 0.69 3.7 1.21 ;
      RECT  1.35 1.21 3.79 1.22 ;
      RECT  1.35 1.22 4.85 1.23 ;
      RECT  0.315 1.23 4.85 1.35 ;
    END
    ANTENNADIFFAREA 1.058 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.82 0.2 4.085 0.26 ;
      RECT  1.86 0.26 4.085 0.27 ;
      RECT  1.86 0.27 5.075 0.375 ;
      RECT  4.955 0.165 5.075 0.27 ;
      RECT  0.09 0.315 0.21 0.52 ;
      RECT  0.09 0.52 3.32 0.62 ;
      RECT  1.075 0.62 2.34 0.67 ;
      RECT  3.22 0.62 3.32 0.7 ;
  END
END SEN_ND3_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_0P5
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_0P5
  CLASS CORE ;
  FOREIGN SEN_ND3_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.9 ;
      RECT  0.35 0.9 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.21 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.59 1.415 0.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.07 0.05 0.21 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.8 0.265 1.05 0.38 ;
      RECT  0.95 0.38 1.05 1.225 ;
      RECT  0.34 1.225 1.05 1.325 ;
      RECT  0.86 1.325 0.98 1.595 ;
      RECT  0.34 1.325 0.46 1.61 ;
    END
    ANTENNADIFFAREA 0.128 ;
  END X
END SEN_ND3_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_0P65
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_0P65
  CLASS CORE ;
  FOREIGN SEN_ND3_T_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0384 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.21 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.6 1.415 0.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.07 0.05 0.21 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.79 0.26 1.05 0.38 ;
      RECT  0.95 0.38 1.05 1.225 ;
      RECT  0.34 1.225 1.05 1.325 ;
      RECT  0.34 1.325 0.46 1.525 ;
      RECT  0.86 1.325 0.98 1.54 ;
    END
    ANTENNADIFFAREA 0.166 ;
  END X
END SEN_ND3_T_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_0P8
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_0P8
  CLASS CORE ;
  FOREIGN SEN_ND3_T_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0585 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0585 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.35 1.41 0.49 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.915 1.415 1.035 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.355 0.05 0.48 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.175 0.165 1.295 0.26 ;
      RECT  0.95 0.26 1.295 0.38 ;
      RECT  0.95 0.38 1.05 1.225 ;
      RECT  0.655 1.225 1.295 1.325 ;
      RECT  0.655 1.325 0.775 1.52 ;
      RECT  1.15 1.325 1.295 1.52 ;
    END
    ANTENNADIFFAREA 0.214 ;
  END X
END SEN_ND3_T_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_1
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_1
  CLASS CORE ;
  FOREIGN SEN_ND3_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0588 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.75 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0738 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.63 1.415 0.77 1.75 ;
      RECT  1.37 1.41 1.51 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.095 0.05 1.215 0.37 ;
      RECT  1.605 0.05 1.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.265 0.185 0.44 ;
      RECT  0.065 0.44 0.45 0.56 ;
      RECT  0.35 0.56 0.45 1.215 ;
      RECT  0.35 1.215 1.26 1.325 ;
      RECT  0.35 1.325 0.45 1.405 ;
      RECT  0.325 1.405 0.45 1.585 ;
    END
    ANTENNADIFFAREA 0.264 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.225 1.005 0.345 ;
      RECT  0.56 0.46 1.525 0.565 ;
  END
END SEN_ND3_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_12
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_12
  CLASS CORE ;
  FOREIGN SEN_ND3_T_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.45 0.81 ;
      RECT  0.15 0.81 2.585 0.92 ;
      RECT  0.15 0.92 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7056 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.25 0.895 ;
      RECT  5.15 0.895 6.305 0.91 ;
      RECT  3.95 0.91 6.305 1.0 ;
      RECT  3.95 1.0 5.25 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8844 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.75 0.71 10.85 0.91 ;
      RECT  7.685 0.91 10.85 1.025 ;
      RECT  9.35 1.025 10.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8844 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 11.0 1.85 ;
      RECT  0.585 1.45 0.705 1.75 ;
      RECT  1.105 1.45 1.225 1.75 ;
      RECT  1.625 1.45 1.745 1.75 ;
      RECT  2.145 1.45 2.265 1.75 ;
      RECT  2.665 1.45 2.785 1.75 ;
      RECT  3.185 1.45 3.305 1.75 ;
      RECT  3.705 1.45 3.825 1.75 ;
      RECT  4.225 1.45 4.345 1.75 ;
      RECT  4.745 1.45 4.865 1.75 ;
      RECT  5.265 1.45 5.385 1.75 ;
      RECT  5.785 1.45 5.905 1.75 ;
      RECT  6.305 1.45 6.425 1.75 ;
      RECT  6.825 1.45 6.945 1.75 ;
      RECT  7.345 1.45 7.465 1.75 ;
      RECT  7.865 1.45 7.985 1.75 ;
      RECT  8.385 1.45 8.505 1.75 ;
      RECT  8.905 1.45 9.025 1.75 ;
      RECT  9.425 1.45 9.545 1.75 ;
      RECT  9.945 1.45 10.065 1.75 ;
      RECT  10.465 1.45 10.585 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      RECT  7.085 0.05 7.205 0.385 ;
      RECT  7.605 0.05 7.725 0.385 ;
      RECT  8.125 0.05 8.245 0.385 ;
      RECT  8.645 0.05 8.765 0.385 ;
      RECT  9.165 0.05 9.285 0.385 ;
      RECT  9.685 0.05 9.805 0.385 ;
      RECT  10.205 0.05 10.325 0.385 ;
      RECT  10.76 0.05 10.88 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 1.11 7.655 1.135 ;
      RECT  5.35 1.135 9.25 1.2 ;
      RECT  0.275 0.49 3.05 0.6 ;
      RECT  1.55 0.6 3.05 0.69 ;
      RECT  2.75 0.69 3.05 1.11 ;
      RECT  0.34 1.11 3.85 1.2 ;
      RECT  0.34 1.2 9.25 1.23 ;
      RECT  0.34 1.23 10.87 1.36 ;
    END
    ANTENNADIFFAREA 2.404 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.15 0.16 4.84 0.21 ;
      RECT  0.065 0.21 6.955 0.38 ;
      RECT  10.465 0.395 10.585 0.49 ;
      RECT  3.385 0.49 10.585 0.62 ;
      RECT  5.35 0.62 10.585 0.66 ;
      RECT  5.35 0.66 8.67 0.74 ;
  END
END SEN_ND3_T_12
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_16
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_16
  CLASS CORE ;
  FOREIGN SEN_ND3_T_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 14.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.905 ;
      RECT  0.15 0.905 3.7 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9396 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.25 0.885 ;
      RECT  5.15 0.885 7.65 0.905 ;
      RECT  5.15 0.905 8.5 1.0 ;
      RECT  5.15 1.0 7.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1763 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  14.15 0.71 14.25 0.905 ;
      RECT  10.315 0.905 14.25 1.0 ;
      RECT  11.95 1.0 14.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1763 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 14.4 1.85 ;
      RECT  0.56 1.46 0.73 1.75 ;
      RECT  1.08 1.46 1.25 1.75 ;
      RECT  1.6 1.46 1.77 1.75 ;
      RECT  2.12 1.49 2.29 1.75 ;
      RECT  2.64 1.49 2.81 1.75 ;
      RECT  3.16 1.49 3.33 1.75 ;
      RECT  3.68 1.49 3.85 1.75 ;
      RECT  4.205 1.49 4.375 1.75 ;
      RECT  4.725 1.49 4.895 1.75 ;
      RECT  5.245 1.49 5.415 1.75 ;
      RECT  5.765 1.49 5.935 1.75 ;
      RECT  6.285 1.49 6.455 1.75 ;
      RECT  6.805 1.49 6.975 1.75 ;
      RECT  7.325 1.49 7.495 1.75 ;
      RECT  7.845 1.49 8.015 1.75 ;
      RECT  8.365 1.49 8.535 1.75 ;
      RECT  8.885 1.49 9.055 1.75 ;
      RECT  9.405 1.49 9.575 1.75 ;
      RECT  9.925 1.49 10.095 1.75 ;
      RECT  10.445 1.49 10.615 1.75 ;
      RECT  10.965 1.49 11.135 1.75 ;
      RECT  11.485 1.49 11.655 1.75 ;
      RECT  12.005 1.49 12.175 1.75 ;
      RECT  12.525 1.49 12.695 1.75 ;
      RECT  13.045 1.49 13.215 1.75 ;
      RECT  13.565 1.49 13.735 1.75 ;
      RECT  14.15 1.21 14.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 14.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 14.4 0.05 ;
      RECT  9.43 0.05 9.55 0.385 ;
      RECT  9.95 0.05 10.07 0.385 ;
      RECT  10.47 0.05 10.59 0.385 ;
      RECT  10.99 0.05 11.11 0.385 ;
      RECT  11.51 0.05 11.63 0.385 ;
      RECT  12.03 0.05 12.15 0.385 ;
      RECT  12.55 0.05 12.67 0.385 ;
      RECT  13.07 0.05 13.19 0.385 ;
      RECT  13.59 0.05 13.71 0.385 ;
      RECT  14.15 0.05 14.27 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 14.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 1.09 10.25 1.11 ;
      RECT  7.75 1.11 11.85 1.2 ;
      RECT  0.34 0.51 4.25 0.69 ;
      RECT  2.35 0.69 4.25 0.795 ;
      RECT  3.93 0.795 4.25 1.08 ;
      RECT  3.93 1.08 5.05 1.2 ;
      RECT  0.325 1.2 13.955 1.37 ;
      RECT  2.385 1.37 13.955 1.4 ;
    END
    ANTENNADIFFAREA 3.197 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.35 0.16 6.45 0.19 ;
      RECT  2.35 0.19 9.015 0.215 ;
      RECT  0.08 0.215 9.015 0.4 ;
      RECT  4.44 0.51 14.015 0.62 ;
      RECT  5.975 0.62 14.015 0.68 ;
      RECT  11.745 0.68 11.915 0.685 ;
      RECT  7.75 0.68 11.45 0.795 ;
      RECT  8.55 0.795 10.25 0.82 ;
  END
END SEN_ND3_T_16
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_1P5
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_1P5
  CLASS CORE ;
  FOREIGN SEN_ND3_T_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.95 ;
      RECT  0.15 0.95 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.087 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.34 0.94 ;
      RECT  0.95 0.94 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1101 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.625 0.71 2.05 0.95 ;
      RECT  1.95 0.95 2.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1101 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.21 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.59 1.445 0.73 1.75 ;
      RECT  1.245 1.445 1.38 1.75 ;
      RECT  1.91 1.41 2.05 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.64 0.05 1.76 0.355 ;
      RECT  2.175 0.05 2.305 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.31 0.435 0.65 0.555 ;
      RECT  0.55 0.555 0.65 1.23 ;
      RECT  0.55 1.23 1.825 1.235 ;
      RECT  0.34 1.235 1.825 1.355 ;
      RECT  0.34 1.355 0.46 1.53 ;
    END
    ANTENNADIFFAREA 0.294 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.225 1.295 0.345 ;
      RECT  0.08 0.345 0.2 0.46 ;
      RECT  0.81 0.445 2.07 0.565 ;
  END
END SEN_ND3_T_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_2
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_2
  CLASS CORE ;
  FOREIGN SEN_ND3_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.95 ;
      RECT  0.15 0.95 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1176 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.34 0.945 ;
      RECT  0.95 0.945 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1476 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.64 0.71 2.05 0.945 ;
      RECT  1.95 0.945 2.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1476 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.21 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.59 1.44 0.73 1.75 ;
      RECT  1.24 1.44 1.38 1.75 ;
      RECT  1.92 1.41 2.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.64 0.05 1.76 0.355 ;
      RECT  2.17 0.05 2.29 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.29 0.44 0.65 0.56 ;
      RECT  0.55 0.56 0.65 1.22 ;
      RECT  0.55 1.22 1.81 1.235 ;
      RECT  0.34 1.235 1.81 1.35 ;
      RECT  0.34 1.35 0.46 1.49 ;
    END
    ANTENNADIFFAREA 0.396 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.225 1.29 0.345 ;
      RECT  0.08 0.345 0.2 0.5 ;
      RECT  1.9 0.34 2.02 0.445 ;
      RECT  0.81 0.445 2.02 0.565 ;
  END
END SEN_ND3_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_3
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_3
  CLASS CORE ;
  FOREIGN SEN_ND3_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.945 ;
      RECT  0.15 0.945 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1764 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.695 0.965 ;
      RECT  1.35 0.965 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.5 0.71 2.85 0.985 ;
      RECT  2.75 0.985 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.575 1.415 0.715 1.75 ;
      RECT  1.095 1.415 1.235 1.75 ;
      RECT  1.66 1.415 1.8 1.75 ;
      RECT  2.395 1.415 2.515 1.75 ;
      RECT  2.925 1.21 3.045 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  2.135 0.05 2.255 0.37 ;
      RECT  2.655 0.05 2.775 0.37 ;
      RECT  3.185 0.05 3.305 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.065 0.285 0.185 0.44 ;
      RECT  0.065 0.44 0.85 0.56 ;
      RECT  0.75 0.56 0.85 1.215 ;
      RECT  0.275 1.215 2.825 1.325 ;
    END
    ANTENNADIFFAREA 0.653 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 0.225 2.03 0.345 ;
      RECT  2.915 0.36 3.035 0.46 ;
      RECT  1.055 0.46 3.035 0.58 ;
  END
END SEN_ND3_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_4
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_4
  CLASS CORE ;
  FOREIGN SEN_ND3_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.65 0.945 ;
      RECT  3.55 0.945 3.65 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2352 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.55 0.91 2.295 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2943 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 1.085 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2943 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.585 1.445 0.705 1.75 ;
      RECT  1.105 1.445 1.225 1.75 ;
      RECT  1.625 1.445 1.745 1.75 ;
      RECT  2.145 1.445 2.265 1.75 ;
      RECT  2.665 1.445 2.785 1.75 ;
      RECT  3.185 1.445 3.305 1.75 ;
      RECT  3.74 1.215 3.86 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.445 3.615 0.555 ;
      RECT  2.75 0.555 2.85 1.235 ;
      RECT  0.275 1.235 3.615 1.355 ;
    END
    ANTENNADIFFAREA 0.79 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.6 0.22 3.825 0.33 ;
      RECT  3.705 0.33 3.825 0.48 ;
      RECT  0.275 0.44 2.575 0.56 ;
  END
END SEN_ND3_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_6
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_6
  CLASS CORE ;
  FOREIGN SEN_ND3_T_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.71 6.25 0.945 ;
      RECT  6.15 0.945 6.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3528 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.25 0.91 ;
      RECT  3.15 0.91 4.495 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.441 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.91 ;
      RECT  0.935 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.441 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.42 1.48 0.59 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.98 1.48 1.15 1.75 ;
      RECT  1.5 1.48 1.67 1.75 ;
      RECT  2.02 1.48 2.19 1.75 ;
      RECT  2.54 1.48 2.71 1.75 ;
      RECT  3.06 1.48 3.23 1.75 ;
      RECT  3.58 1.48 3.75 1.75 ;
      RECT  4.1 1.48 4.27 1.75 ;
      RECT  4.62 1.48 4.79 1.75 ;
      RECT  5.165 1.415 5.285 1.75 ;
      RECT  5.685 1.415 5.8 1.75 ;
      RECT  6.205 1.21 6.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  0.445 0.05 0.565 0.355 ;
      RECT  1.005 0.05 1.125 0.355 ;
      RECT  1.525 0.05 1.645 0.355 ;
      RECT  2.045 0.05 2.165 0.355 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.72 0.47 6.115 0.595 ;
      RECT  4.72 0.595 4.85 1.11 ;
      RECT  4.72 1.11 6.06 1.26 ;
      RECT  0.095 1.26 6.06 1.29 ;
      RECT  0.095 1.29 4.85 1.39 ;
    END
    ANTENNADIFFAREA 1.215 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.54 0.21 6.325 0.34 ;
      RECT  6.205 0.34 6.325 0.455 ;
      RECT  0.095 0.45 4.555 0.62 ;
  END
END SEN_ND3_T_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3_T_8
#      Description : "3-Input NAND"
#      Equation    : X=!(A1&A2&A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3_T_8
  CLASS CORE ;
  FOREIGN SEN_ND3_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.915 0.925 ;
      RECT  0.15 0.925 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4698 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.05 0.91 ;
      RECT  2.95 0.91 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5904 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.25 0.895 ;
      RECT  5.75 0.895 7.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5904 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  0.59 1.415 0.71 1.75 ;
      RECT  1.11 1.415 1.23 1.75 ;
      RECT  1.63 1.42 1.75 1.75 ;
      RECT  2.15 1.435 2.27 1.75 ;
      RECT  2.67 1.435 2.79 1.75 ;
      RECT  3.19 1.435 3.31 1.75 ;
      RECT  3.71 1.435 3.83 1.75 ;
      RECT  4.23 1.43 4.35 1.75 ;
      RECT  4.75 1.435 4.87 1.75 ;
      RECT  5.27 1.435 5.39 1.75 ;
      RECT  5.79 1.435 5.91 1.75 ;
      RECT  6.31 1.435 6.43 1.75 ;
      RECT  6.85 1.42 6.97 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  4.75 0.05 4.87 0.36 ;
      RECT  5.27 0.05 5.39 0.36 ;
      RECT  5.79 0.05 5.91 0.36 ;
      RECT  6.31 0.05 6.43 0.36 ;
      RECT  6.85 0.05 6.97 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.43 2.255 0.47 ;
      RECT  0.28 0.47 2.255 0.6 ;
      RECT  2.085 0.6 2.255 1.11 ;
      RECT  0.34 1.11 2.85 1.2 ;
      RECT  0.34 1.2 7.25 1.29 ;
      RECT  4.15 1.11 5.65 1.2 ;
      RECT  1.75 1.29 7.25 1.33 ;
      RECT  7.15 1.33 7.25 1.49 ;
    END
    ANTENNADIFFAREA 1.616 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.4 0.16 3.02 0.19 ;
      RECT  1.4 0.19 4.4 0.2 ;
      RECT  0.07 0.2 4.4 0.32 ;
      RECT  0.07 0.32 0.19 0.475 ;
      RECT  3.765 0.45 5.625 0.49 ;
      RECT  2.36 0.49 7.26 0.62 ;
      RECT  7.14 0.345 7.26 0.49 ;
  END
END SEN_ND3_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_0P5
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_0P5
  CLASS CORE ;
  FOREIGN SEN_ND3B_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.13 0.7 0.25 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.85 0.98 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.705 ;
      RECT  0.52 0.705 0.65 0.98 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.425 0.445 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.845 1.455 0.965 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.325 0.05 0.445 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.105 0.175 1.25 0.375 ;
      RECT  1.15 0.375 1.25 1.255 ;
      RECT  0.55 1.255 1.25 1.345 ;
      RECT  0.55 1.345 0.705 1.59 ;
      RECT  1.105 1.345 1.25 1.605 ;
    END
    ANTENNADIFFAREA 0.129 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.205 0.185 0.475 ;
      RECT  0.065 0.475 0.43 0.59 ;
      RECT  0.34 0.59 0.43 1.075 ;
      RECT  0.34 1.075 1.06 1.165 ;
      RECT  0.96 0.485 1.06 1.075 ;
      RECT  0.34 1.165 0.43 1.21 ;
      RECT  0.065 1.21 0.43 1.315 ;
      RECT  0.065 1.315 0.185 1.61 ;
  END
END SEN_ND3B_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_1
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_1
  CLASS CORE ;
  FOREIGN SEN_ND3B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0498 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.865 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.73 ;
      RECT  0.52 0.73 0.65 0.92 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.365 1.45 0.495 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.935 1.445 1.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.305 0.05 0.505 0.21 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.35 0.69 ;
      RECT  1.26 0.69 1.35 1.11 ;
      RECT  1.15 1.11 1.35 1.235 ;
      RECT  0.6 1.235 1.35 1.355 ;
      RECT  1.15 1.355 1.35 1.49 ;
    END
    ANTENNADIFFAREA 0.298 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.955 0.82 1.17 0.93 ;
      RECT  0.955 0.93 1.045 1.055 ;
      RECT  0.07 0.18 0.19 0.3 ;
      RECT  0.07 0.3 0.43 0.39 ;
      RECT  0.34 0.39 0.43 1.055 ;
      RECT  0.34 1.055 1.045 1.145 ;
      RECT  0.34 1.145 0.43 1.24 ;
      RECT  0.07 1.24 0.43 1.34 ;
      RECT  0.07 1.34 0.19 1.46 ;
  END
END SEN_ND3B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_2
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_2
  CLASS CORE ;
  FOREIGN SEN_ND3B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0996 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 0.71 ;
      RECT  1.55 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.5 0.65 0.71 ;
      RECT  0.55 0.71 1.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.585 1.215 0.705 1.75 ;
      RECT  1.245 1.415 1.385 1.75 ;
      RECT  1.885 1.415 2.025 1.75 ;
      RECT  2.415 1.425 2.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.105 0.05 1.225 0.37 ;
      RECT  0.575 0.05 0.72 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.155 0.465 2.45 0.635 ;
      RECT  2.35 0.635 2.45 1.195 ;
      RECT  0.82 1.195 2.45 1.315 ;
    END
    ANTENNADIFFAREA 0.45 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.415 0.17 2.535 0.245 ;
      RECT  1.335 0.245 2.535 0.365 ;
      RECT  0.79 0.47 1.81 0.59 ;
      RECT  0.34 0.33 0.445 1.01 ;
      RECT  0.34 1.01 2.25 1.1 ;
      RECT  2.15 0.755 2.25 1.01 ;
      RECT  0.34 1.1 0.445 1.38 ;
  END
END SEN_ND3B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_4
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_4
  CLASS CORE ;
  FOREIGN SEN_ND3B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1992 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.45 0.71 ;
      RECT  2.85 0.71 3.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.5 1.25 0.71 ;
      RECT  1.15 0.71 1.725 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.185 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.585 1.41 0.705 1.75 ;
      RECT  1.105 1.41 1.225 1.75 ;
      RECT  1.625 1.435 1.745 1.75 ;
      RECT  2.24 1.435 2.36 1.75 ;
      RECT  2.865 1.435 2.985 1.75 ;
      RECT  3.385 1.435 3.505 1.75 ;
      RECT  3.905 1.435 4.03 1.75 ;
      RECT  4.425 1.44 4.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.585 0.05 0.705 0.36 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  1.625 0.05 1.745 0.365 ;
      RECT  2.145 0.05 2.265 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.51 4.45 0.69 ;
      RECT  4.35 0.69 4.45 1.21 ;
      RECT  1.31 1.21 4.45 1.34 ;
    END
    ANTENNADIFFAREA 0.9 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.355 0.2 4.545 0.32 ;
      RECT  4.425 0.32 4.545 0.39 ;
      RECT  2.355 0.32 2.465 0.68 ;
      RECT  2.605 0.425 3.245 0.545 ;
      RECT  3.125 0.545 3.245 0.595 ;
      RECT  2.605 0.545 2.725 0.77 ;
      RECT  1.34 0.475 2.02 0.595 ;
      RECT  1.885 0.595 2.02 0.77 ;
      RECT  1.885 0.77 2.725 0.89 ;
      RECT  3.635 0.785 4.26 0.895 ;
      RECT  3.635 0.895 3.745 0.98 ;
      RECT  0.295 0.45 1.05 0.57 ;
      RECT  0.96 0.57 1.05 0.98 ;
      RECT  0.96 0.98 3.745 1.07 ;
      RECT  0.96 1.07 1.05 1.135 ;
      RECT  0.34 1.135 1.05 1.26 ;
      RECT  0.34 1.26 0.445 1.38 ;
  END
END SEN_ND3B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_8
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_8
  CLASS CORE ;
  FOREIGN SEN_ND3B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 0.87 ;
      RECT  3.15 0.87 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4698 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.65 0.895 ;
      RECT  5.15 0.895 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4698 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.445 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.845 1.415 0.965 1.75 ;
      RECT  1.34 1.48 1.51 1.75 ;
      RECT  1.86 1.48 2.03 1.75 ;
      RECT  2.38 1.48 2.55 1.75 ;
      RECT  2.9 1.48 3.07 1.75 ;
      RECT  3.42 1.48 3.59 1.75 ;
      RECT  3.94 1.48 4.11 1.75 ;
      RECT  4.46 1.48 4.63 1.75 ;
      RECT  4.98 1.48 5.15 1.75 ;
      RECT  5.5 1.48 5.67 1.75 ;
      RECT  6.02 1.48 6.19 1.75 ;
      RECT  6.54 1.48 6.71 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  5.005 0.05 5.125 0.345 ;
      RECT  5.525 0.05 5.645 0.345 ;
      RECT  6.045 0.05 6.165 0.345 ;
      RECT  6.565 0.05 6.685 0.345 ;
      RECT  0.865 0.05 0.985 0.36 ;
      RECT  0.325 0.05 0.445 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 3.05 0.69 ;
      RECT  2.88 0.69 3.05 1.11 ;
      RECT  0.95 1.11 3.05 1.21 ;
      RECT  0.95 1.21 6.945 1.3 ;
      RECT  2.88 1.3 6.945 1.33 ;
      RECT  2.88 1.33 5.945 1.34 ;
      RECT  6.825 1.33 6.945 1.46 ;
      RECT  2.88 1.34 5.44 1.38 ;
    END
    ANTENNADIFFAREA 1.62 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.26 0.2 4.655 0.32 ;
      RECT  2.235 0.32 3.68 0.33 ;
      RECT  6.825 0.31 6.945 0.435 ;
      RECT  3.185 0.435 6.945 0.555 ;
      RECT  4.12 0.555 5.495 0.565 ;
      RECT  3.185 0.555 3.305 0.605 ;
      RECT  0.065 0.335 0.185 0.46 ;
      RECT  0.065 0.46 0.85 0.58 ;
      RECT  0.745 0.58 0.85 0.87 ;
      RECT  0.745 0.87 2.73 0.98 ;
      RECT  0.745 0.98 0.85 1.18 ;
      RECT  0.065 1.18 0.85 1.3 ;
      RECT  0.065 1.3 0.185 1.48 ;
  END
END SEN_ND3B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_V1DG_8
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_V1DG_8
  CLASS CORE ;
  FOREIGN SEN_ND3B_V1DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.71 6.85 0.89 ;
      RECT  6.75 0.89 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.16 4.45 0.25 ;
      RECT  3.55 0.25 3.65 0.455 ;
      RECT  4.35 0.25 4.45 0.455 ;
      RECT  1.95 0.16 3.05 0.25 ;
      RECT  1.95 0.25 2.05 0.45 ;
      RECT  2.95 0.25 3.05 0.455 ;
      RECT  0.95 0.45 2.05 0.53 ;
      RECT  2.95 0.455 3.65 0.53 ;
      RECT  4.35 0.455 5.65 0.545 ;
      RECT  0.95 0.53 2.45 0.55 ;
      RECT  2.95 0.53 4.05 0.545 ;
      RECT  3.55 0.545 4.05 0.62 ;
      RECT  5.55 0.545 5.65 0.925 ;
      RECT  1.95 0.55 2.45 0.62 ;
      RECT  0.95 0.55 1.05 0.925 ;
      RECT  2.35 0.62 2.45 0.925 ;
      RECT  3.95 0.62 4.05 0.925 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.505 6.05 0.925 ;
      RECT  5.15 0.71 5.45 0.925 ;
      RECT  4.35 0.71 4.65 0.925 ;
      RECT  3.55 0.71 3.85 0.925 ;
      RECT  2.75 0.71 3.05 0.925 ;
      RECT  1.95 0.71 2.25 0.925 ;
      RECT  1.25 0.71 1.55 0.925 ;
      RECT  0.49 0.505 0.595 0.925 ;
      LAYER M2 ;
      RECT  0.45 0.75 6.09 0.85 ;
      LAYER V1 ;
      RECT  5.95 0.75 6.05 0.85 ;
      RECT  5.15 0.75 5.25 0.85 ;
      RECT  5.35 0.75 5.45 0.85 ;
      RECT  4.35 0.75 4.45 0.85 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  1.25 0.75 1.35 0.85 ;
      RECT  1.45 0.75 1.55 0.85 ;
      RECT  0.49 0.75 0.59 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.585 1.45 0.705 1.75 ;
      RECT  1.12 1.44 1.21 1.75 ;
      RECT  1.64 1.44 1.73 1.75 ;
      RECT  2.16 1.44 2.25 1.75 ;
      RECT  2.68 1.44 2.77 1.75 ;
      RECT  3.2 1.44 3.29 1.75 ;
      RECT  3.72 1.42 3.81 1.75 ;
      RECT  4.24 1.42 4.33 1.75 ;
      RECT  4.76 1.44 4.85 1.75 ;
      RECT  5.28 1.38 5.37 1.75 ;
      RECT  5.8 1.38 5.89 1.75 ;
      RECT  6.305 1.455 6.425 1.75 ;
      RECT  6.825 1.41 6.945 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  6.305 0.05 6.425 0.35 ;
      RECT  1.625 0.05 1.745 0.36 ;
      RECT  3.185 0.05 3.305 0.365 ;
      RECT  4.745 0.05 4.865 0.365 ;
      RECT  6.825 0.05 6.945 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.47 0.24 5.85 0.36 ;
      RECT  5.75 0.36 5.85 1.11 ;
      RECT  5.005 1.11 6.165 1.14 ;
      RECT  3.915 0.34 4.25 0.44 ;
      RECT  4.15 0.44 4.25 1.11 ;
      RECT  3.445 1.11 4.65 1.14 ;
      RECT  2.355 0.34 2.65 0.44 ;
      RECT  2.55 0.44 2.65 1.11 ;
      RECT  1.95 1.11 3.05 1.14 ;
      RECT  0.75 0.24 1.02 0.36 ;
      RECT  0.75 0.36 0.85 1.11 ;
      RECT  0.34 1.11 1.605 1.14 ;
      RECT  0.34 1.14 6.165 1.29 ;
    END
    ANTENNADIFFAREA 1.824 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.35 0.44 6.735 0.56 ;
      RECT  6.35 0.56 6.45 0.755 ;
      RECT  6.205 0.755 6.45 0.925 ;
      RECT  6.34 0.925 6.45 1.245 ;
      RECT  6.34 1.245 6.735 1.365 ;
      RECT  1.675 0.675 1.775 0.95 ;
      RECT  1.675 0.95 1.855 1.05 ;
      RECT  3.15 0.675 3.25 0.95 ;
      RECT  3.15 0.95 3.33 1.05 ;
      RECT  4.75 0.675 4.85 0.95 ;
      RECT  4.75 0.95 4.93 1.05 ;
      RECT  0.13 0.68 0.25 1.1 ;
      LAYER M2 ;
      RECT  0.11 0.95 6.49 1.05 ;
      LAYER V1 ;
      RECT  0.15 0.95 0.25 1.05 ;
      RECT  1.715 0.95 1.815 1.05 ;
      RECT  3.19 0.95 3.29 1.05 ;
      RECT  4.79 0.95 4.89 1.05 ;
      RECT  6.35 0.95 6.45 1.05 ;
  END
END SEN_ND3B_V1DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_V1DG_1
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_V1DG_1
  CLASS CORE ;
  FOREIGN SEN_ND3B_V1DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.65 0.25 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.45 1.25 1.02 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.85 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.445 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.845 1.39 0.965 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.315 0.05 0.455 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.24 1.285 0.36 ;
      RECT  0.95 0.36 1.05 1.11 ;
      RECT  0.55 1.11 1.25 1.29 ;
    END
    ANTENNADIFFAREA 0.293 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.195 0.185 0.45 ;
      RECT  0.065 0.45 0.45 0.55 ;
      RECT  0.35 0.55 0.45 0.755 ;
      RECT  0.35 0.755 0.545 0.925 ;
      RECT  0.35 0.925 0.455 1.25 ;
      RECT  0.065 1.25 0.455 1.35 ;
      RECT  0.065 1.35 0.185 1.58 ;
  END
END SEN_ND3B_V1DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_V1DG_2
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_V1DG_2
  CLASS CORE ;
  FOREIGN SEN_ND3B_V1DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.64 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.71 ;
      RECT  1.95 0.71 2.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 0.71 ;
      RECT  1.35 0.71 1.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.535 1.38 0.655 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.095 1.38 1.215 1.75 ;
      RECT  1.615 1.38 1.735 1.75 ;
      RECT  2.165 1.21 2.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.445 2.045 0.555 ;
      RECT  1.75 0.555 1.85 1.11 ;
      RECT  0.75 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.48 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.07 0.245 2.28 0.355 ;
      RECT  0.065 0.21 0.185 0.45 ;
      RECT  0.065 0.45 0.45 0.55 ;
      RECT  0.35 0.55 0.45 0.785 ;
      RECT  0.35 0.785 0.87 0.895 ;
      RECT  0.35 0.895 0.45 1.26 ;
      RECT  0.065 1.26 0.45 1.35 ;
      RECT  0.065 1.35 0.185 1.59 ;
      RECT  0.54 0.45 1.46 0.57 ;
      RECT  1.355 0.57 1.46 0.62 ;
  END
END SEN_ND3B_V1DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND3B_V1DG_4
#      Description : "3-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND3B_V1DG_4
  CLASS CORE ;
  FOREIGN SEN_ND3B_V1DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.65 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.685 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  1.15 0.71 1.895 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.085 1.21 0.205 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  0.63 1.39 0.75 1.75 ;
      RECT  1.15 1.39 1.27 1.75 ;
      RECT  1.84 1.39 1.96 1.75 ;
      RECT  2.4 1.39 2.52 1.75 ;
      RECT  2.96 1.39 3.08 1.75 ;
      RECT  3.48 1.45 3.6 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  3.48 0.05 3.6 0.35 ;
      RECT  2.44 0.05 2.56 0.36 ;
      RECT  2.96 0.05 3.08 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.345 0.445 1.05 0.555 ;
      RECT  0.95 0.555 1.05 1.11 ;
      RECT  0.35 1.11 3.355 1.29 ;
    END
    ANTENNADIFFAREA 1.014 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.11 0.245 2.335 0.355 ;
      RECT  0.11 0.355 0.23 0.49 ;
      RECT  1.36 0.45 3.39 0.56 ;
      RECT  3.555 0.44 3.885 0.56 ;
      RECT  3.555 0.56 3.645 0.785 ;
      RECT  2.92 0.785 3.645 0.895 ;
      RECT  3.555 0.895 3.645 1.24 ;
      RECT  3.555 1.24 3.885 1.36 ;
  END
END SEN_ND3B_V1DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_1
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_1
  CLASS CORE ;
  FOREIGN SEN_ND4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.71 ;
      RECT  0.35 0.71 0.65 0.915 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.085 1.41 0.215 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.665 1.41 0.795 1.75 ;
      RECT  1.195 1.41 1.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.085 0.05 0.215 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.25 1.345 0.37 ;
      RECT  0.95 0.37 1.05 1.21 ;
      RECT  0.34 1.21 1.05 1.32 ;
    END
    ANTENNADIFFAREA 0.322 ;
  END X
END SEN_ND4_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_2
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_2
  CLASS CORE ;
  FOREIGN SEN_ND4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.585 1.41 0.715 1.75 ;
      RECT  1.24 1.41 1.37 1.75 ;
      RECT  1.875 1.41 2.005 1.75 ;
      RECT  2.4 1.21 2.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.325 0.05 0.455 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.41 2.25 1.21 ;
      RECT  0.345 1.21 2.25 1.31 ;
      RECT  0.345 1.31 0.45 1.5 ;
    END
    ANTENNADIFFAREA 0.544 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.895 0.19 2.52 0.29 ;
      RECT  2.4 0.29 2.52 0.39 ;
      RECT  1.895 0.29 2.01 0.48 ;
      RECT  1.36 0.48 2.01 0.59 ;
      RECT  1.36 0.59 1.48 0.65 ;
      RECT  0.8 0.24 1.785 0.36 ;
      RECT  0.07 0.36 0.19 0.48 ;
      RECT  0.07 0.48 1.23 0.58 ;
      RECT  1.12 0.58 1.23 0.65 ;
  END
END SEN_ND4_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_4
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_4
  CLASS CORE ;
  FOREIGN SEN_ND4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  2.75 0.89 2.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.585 1.455 0.715 1.75 ;
      RECT  1.11 1.455 1.23 1.75 ;
      RECT  1.625 1.455 1.755 1.75 ;
      RECT  2.235 1.455 2.365 1.75 ;
      RECT  2.85 1.455 2.98 1.75 ;
      RECT  3.37 1.455 3.5 1.75 ;
      RECT  3.9 1.455 4.03 1.75 ;
      RECT  4.42 1.41 4.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.325 0.05 0.455 0.385 ;
      RECT  0.845 0.05 0.975 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.615 0.45 4.31 0.57 ;
      RECT  3.75 0.57 3.85 1.235 ;
      RECT  3.75 1.235 4.33 1.24 ;
      RECT  0.33 1.24 4.33 1.365 ;
      RECT  0.33 1.365 0.45 1.49 ;
    END
    ANTENNADIFFAREA 1.098 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.95 0.14 2.665 0.23 ;
      RECT  1.95 0.23 2.06 0.24 ;
      RECT  2.57 0.23 2.665 0.24 ;
      RECT  1.32 0.24 2.06 0.36 ;
      RECT  2.57 0.24 3.265 0.36 ;
      RECT  3.375 0.235 4.535 0.355 ;
      RECT  4.425 0.355 4.535 0.43 ;
      RECT  3.375 0.355 3.495 0.48 ;
      RECT  2.28 0.32 2.48 0.425 ;
      RECT  2.39 0.425 2.48 0.48 ;
      RECT  2.39 0.48 3.495 0.6 ;
      RECT  0.07 0.37 0.19 0.48 ;
      RECT  0.07 0.48 2.16 0.545 ;
      RECT  0.07 0.545 2.295 0.59 ;
      RECT  2.075 0.59 2.295 0.665 ;
  END
END SEN_ND4_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_8
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_8
  CLASS CORE ;
  FOREIGN SEN_ND4_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.75 0.51 8.85 0.71 ;
      RECT  7.35 0.71 8.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.85 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 4.05 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.65 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 9.0 1.85 ;
      RECT  0.565 1.28 0.735 1.75 ;
      RECT  1.085 1.28 1.255 1.75 ;
      RECT  1.605 1.28 1.775 1.75 ;
      RECT  2.125 1.28 2.295 1.75 ;
      RECT  2.665 1.29 2.795 1.75 ;
      RECT  3.165 1.465 3.335 1.75 ;
      RECT  3.685 1.465 3.855 1.75 ;
      RECT  4.205 1.465 4.375 1.75 ;
      RECT  4.725 1.465 4.895 1.75 ;
      RECT  5.245 1.465 5.415 1.75 ;
      RECT  5.765 1.465 5.935 1.75 ;
      RECT  6.285 1.465 6.455 1.75 ;
      RECT  6.825 1.38 6.955 1.75 ;
      RECT  7.345 1.38 7.475 1.75 ;
      RECT  7.865 1.38 7.995 1.75 ;
      RECT  8.435 1.38 8.565 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      RECT  1.345 0.05 1.515 0.335 ;
      RECT  1.865 0.05 2.035 0.335 ;
      RECT  0.33 0.05 0.45 0.4 ;
      RECT  0.85 0.05 0.97 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.865 0.44 8.61 0.59 ;
      RECT  6.865 0.59 7.05 1.11 ;
      RECT  5.95 1.11 8.85 1.205 ;
      RECT  0.34 1.03 3.06 1.19 ;
      RECT  2.89 1.19 3.06 1.205 ;
      RECT  0.34 1.19 0.45 1.29 ;
      RECT  2.89 1.205 8.85 1.29 ;
      RECT  2.89 1.29 6.095 1.375 ;
    END
    ANTENNADIFFAREA 2.236 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.315 0.16 6.46 0.2 ;
      RECT  2.385 0.2 6.46 0.33 ;
      RECT  6.56 0.18 8.885 0.35 ;
      RECT  6.56 0.35 6.73 0.425 ;
      RECT  4.47 0.425 6.73 0.585 ;
      RECT  0.07 0.39 0.19 0.49 ;
      RECT  0.07 0.49 4.375 0.61 ;
      RECT  1.62 0.47 4.375 0.49 ;
      RECT  1.08 0.61 4.375 0.62 ;
  END
END SEN_ND4_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_S_0P5
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_S_0P5
  CLASS CORE ;
  FOREIGN SEN_ND4_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.145 0.51 1.255 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.89 ;
      RECT  0.35 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0237 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.635 1.44 0.755 1.75 ;
      RECT  1.19 1.41 1.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.06 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.2 0.175 1.32 0.29 ;
      RECT  0.95 0.29 1.32 0.4 ;
      RECT  0.95 0.4 1.05 1.235 ;
      RECT  0.35 1.235 1.05 1.325 ;
      RECT  0.35 1.325 0.45 1.64 ;
      RECT  0.95 1.325 1.05 1.64 ;
    END
    ANTENNADIFFAREA 0.114 ;
  END X
END SEN_ND4_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_S_1
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_S_1
  CLASS CORE ;
  FOREIGN SEN_ND4_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.85 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 0.91 ;
      RECT  0.35 0.91 0.65 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0426 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.21 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.68 1.455 0.8 1.75 ;
      RECT  1.19 1.41 1.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.07 0.05 0.21 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.2 0.15 1.32 0.285 ;
      RECT  0.95 0.285 1.32 0.39 ;
      RECT  0.95 0.39 1.05 1.275 ;
      RECT  0.35 1.275 1.05 1.365 ;
      RECT  0.35 1.365 0.45 1.59 ;
      RECT  0.95 1.365 1.05 1.59 ;
    END
    ANTENNADIFFAREA 0.179 ;
  END X
END SEN_ND4_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_S_1P5
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_S_1P5
  CLASS CORE ;
  FOREIGN SEN_ND4_S_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.34 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0633 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.46 1.075 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0633 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0633 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0633 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.23 1.41 0.37 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.79 1.48 0.96 1.75 ;
      RECT  1.415 1.475 1.585 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.315 0.05 0.455 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.41 1.45 1.255 ;
      RECT  0.5 1.255 1.45 1.375 ;
    END
    ANTENNADIFFAREA 0.208 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.02 0.2 1.72 0.32 ;
      RECT  1.6 0.32 1.72 0.42 ;
      RECT  0.065 0.31 0.185 0.435 ;
      RECT  0.065 0.435 0.755 0.555 ;
  END
END SEN_ND4_S_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_S_2
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_S_2
  CLASS CORE ;
  FOREIGN SEN_ND4_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.85 0.45 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0852 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 0.85 ;
      RECT  0.75 0.85 1.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0852 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.85 ;
      RECT  1.55 0.85 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0852 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0852 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.23 1.41 0.37 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.24 1.455 1.36 1.75 ;
      RECT  2.23 1.41 2.37 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  2.135 0.05 2.255 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.265 0.44 0.65 0.56 ;
      RECT  0.55 0.56 0.65 1.24 ;
      RECT  0.55 1.24 1.94 1.36 ;
    END
    ANTENNADIFFAREA 0.52 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.2 1.24 0.335 ;
      RECT  0.055 0.335 0.175 0.41 ;
      RECT  1.33 0.215 1.995 0.335 ;
      RECT  1.875 0.335 1.995 0.44 ;
      RECT  1.875 0.44 2.515 0.56 ;
      RECT  2.395 0.32 2.515 0.44 ;
      RECT  0.785 0.44 1.785 0.56 ;
  END
END SEN_ND4_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_S_3
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_S_3
  CLASS CORE ;
  FOREIGN SEN_ND4_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 2.85 0.885 ;
      RECT  2.55 0.885 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1278 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.05 0.91 ;
      RECT  1.75 0.91 2.05 1.145 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1278 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 0.91 ;
      RECT  0.95 0.91 1.45 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1278 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.31 0.91 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1278 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.23 1.41 0.37 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.915 1.48 1.085 1.75 ;
      RECT  1.595 1.48 1.765 1.75 ;
      RECT  2.115 1.48 2.285 1.75 ;
      RECT  2.71 1.41 2.85 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.59 0.05 0.71 0.345 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.94 0.305 3.06 0.44 ;
      RECT  2.35 0.44 3.06 0.56 ;
      RECT  2.35 0.56 2.45 1.27 ;
      RECT  0.535 1.27 2.575 1.39 ;
    END
    ANTENNADIFFAREA 0.455 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.14 0.205 2.85 0.32 ;
      RECT  2.14 0.32 2.26 0.44 ;
      RECT  1.62 0.44 2.26 0.56 ;
      RECT  1.62 0.56 1.74 0.705 ;
      RECT  1.055 0.23 2.05 0.35 ;
      RECT  0.28 0.44 1.49 0.56 ;
      RECT  1.37 0.56 1.49 0.71 ;
  END
END SEN_ND4_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_S_4
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_S_4
  CLASS CORE ;
  FOREIGN SEN_ND4_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.25 0.91 ;
      RECT  2.75 0.91 3.25 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1704 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  1.75 0.91 2.25 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1704 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.91 ;
      RECT  1.15 0.91 1.65 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1704 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.35 0.91 0.85 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1704 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.585 1.49 0.755 1.75 ;
      RECT  1.105 1.49 1.275 1.75 ;
      RECT  1.625 1.49 1.795 1.75 ;
      RECT  2.145 1.49 2.315 1.75 ;
      RECT  2.685 1.49 2.855 1.75 ;
      RECT  3.27 1.41 3.41 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.61 0.05 0.73 0.345 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.44 3.375 0.56 ;
      RECT  2.55 0.56 2.65 1.27 ;
      RECT  0.335 1.27 3.09 1.4 ;
      RECT  0.335 1.4 0.46 1.54 ;
      RECT  1.91 1.4 2.05 1.54 ;
      RECT  2.95 1.4 3.09 1.54 ;
    END
    ANTENNADIFFAREA 0.605 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.08 0.23 1.77 0.35 ;
      RECT  1.65 0.35 1.77 0.44 ;
      RECT  1.65 0.44 2.345 0.56 ;
      RECT  1.86 0.23 3.145 0.35 ;
      RECT  0.285 0.44 1.535 0.56 ;
  END
END SEN_ND4_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_S_6
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_S_6
  CLASS CORE ;
  FOREIGN SEN_ND4_S_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 1.11 ;
      RECT  3.95 1.11 4.65 1.22 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2556 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.25 0.91 ;
      RECT  2.75 0.91 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2556 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  1.75 0.91 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2556 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.11 ;
      RECT  0.35 1.11 1.05 1.22 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2556 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.585 1.495 0.755 1.75 ;
      RECT  1.105 1.495 1.275 1.75 ;
      RECT  1.625 1.495 1.795 1.75 ;
      RECT  2.145 1.495 2.315 1.75 ;
      RECT  2.665 1.495 2.835 1.75 ;
      RECT  3.185 1.495 3.355 1.75 ;
      RECT  3.715 1.495 3.885 1.75 ;
      RECT  4.235 1.495 4.405 1.75 ;
      RECT  4.79 1.41 4.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.35 0.05 0.47 0.345 ;
      RECT  0.87 0.05 0.99 0.345 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.44 4.7 0.56 ;
      RECT  3.75 0.56 3.85 1.31 ;
      RECT  0.35 1.31 4.66 1.4 ;
      RECT  2.405 1.4 2.575 1.46 ;
      RECT  0.845 1.4 1.015 1.47 ;
      RECT  3.445 1.4 3.615 1.47 ;
      RECT  3.975 1.4 4.145 1.47 ;
      RECT  1.91 1.4 2.05 1.53 ;
      RECT  2.95 1.4 3.07 1.53 ;
      RECT  0.35 1.4 0.47 1.55 ;
      RECT  1.365 1.4 1.51 1.55 ;
      RECT  4.54 1.4 4.66 1.55 ;
    END
    ANTENNADIFFAREA 0.866 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.13 0.23 2.345 0.35 ;
      RECT  1.13 0.35 1.25 0.44 ;
      RECT  0.09 0.31 0.21 0.44 ;
      RECT  0.09 0.44 1.25 0.56 ;
      RECT  2.635 0.23 4.92 0.35 ;
      RECT  4.8 0.35 4.92 0.46 ;
      RECT  1.34 0.44 3.64 0.56 ;
  END
END SEN_ND4_S_6
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4_S_8
#      Description : "4-Input NAND"
#      Equation    : X=!(A1&A2&A3&A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4_S_8
  CLASS CORE ;
  FOREIGN SEN_ND4_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.25 0.91 ;
      RECT  5.34 0.91 6.25 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3408 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 4.865 0.91 ;
      RECT  3.71 0.91 4.865 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3408 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.05 0.91 ;
      RECT  2.15 0.91 3.05 1.19 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3408 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.91 1.45 1.145 ;
      RECT  0.15 1.145 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3408 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.09 1.41 0.23 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  0.61 1.49 0.78 1.75 ;
      RECT  1.13 1.49 1.3 1.75 ;
      RECT  1.65 1.49 1.82 1.75 ;
      RECT  2.17 1.49 2.34 1.75 ;
      RECT  2.69 1.49 2.86 1.75 ;
      RECT  3.21 1.49 3.38 1.75 ;
      RECT  3.73 1.49 3.9 1.75 ;
      RECT  4.25 1.49 4.42 1.75 ;
      RECT  4.77 1.49 4.94 1.75 ;
      RECT  5.29 1.49 5.46 1.75 ;
      RECT  5.81 1.49 5.98 1.75 ;
      RECT  6.37 1.41 6.51 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.375 0.05 0.495 0.415 ;
      RECT  0.895 0.05 1.015 0.415 ;
      RECT  1.415 0.05 1.535 0.415 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.055 0.44 6.28 0.56 ;
      RECT  5.055 0.56 5.25 1.3 ;
      RECT  0.35 1.3 6.25 1.4 ;
      RECT  0.35 1.4 0.495 1.52 ;
      RECT  0.895 1.4 1.015 1.52 ;
      RECT  1.415 1.4 1.535 1.52 ;
      RECT  1.935 1.4 2.055 1.52 ;
      RECT  2.455 1.4 2.575 1.52 ;
      RECT  2.95 1.4 3.095 1.52 ;
      RECT  3.495 1.4 3.615 1.52 ;
      RECT  4.015 1.4 4.135 1.52 ;
      RECT  4.535 1.4 4.655 1.52 ;
      RECT  5.055 1.4 5.175 1.52 ;
      RECT  5.55 1.4 5.695 1.52 ;
      RECT  6.095 1.4 6.25 1.52 ;
    END
    ANTENNADIFFAREA 1.134 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.88 0.195 4.695 0.315 ;
      RECT  1.88 0.315 4.16 0.32 ;
      RECT  2.43 0.32 4.16 0.345 ;
      RECT  2.95 0.345 3.615 0.365 ;
      RECT  4.785 0.195 6.505 0.32 ;
      RECT  4.785 0.32 5.46 0.345 ;
      RECT  6.385 0.32 6.505 0.425 ;
      RECT  4.785 0.345 4.935 0.445 ;
      RECT  4.25 0.445 4.935 0.475 ;
      RECT  3.175 0.475 4.935 0.595 ;
      RECT  0.09 0.385 0.215 0.54 ;
      RECT  0.09 0.54 2.34 0.55 ;
      RECT  1.13 0.52 2.34 0.54 ;
      RECT  0.09 0.55 2.865 0.67 ;
  END
END SEN_ND4_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4B_1
#      Description : "4-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4B_1
  CLASS CORE ;
  FOREIGN SEN_ND4B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0474 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.755 ;
      RECT  0.695 0.755 0.85 0.935 ;
      RECT  0.75 0.935 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.76 ;
      RECT  0.35 0.76 0.53 0.935 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.58 1.39 0.71 1.75 ;
      RECT  1.215 1.39 1.385 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  1.61 0.05 1.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.25 1.265 0.355 ;
      RECT  0.95 0.355 1.05 1.21 ;
      RECT  0.335 1.21 1.05 1.3 ;
      RECT  0.335 1.3 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.288 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.355 0.38 1.46 0.7 ;
      RECT  1.15 0.7 1.46 0.79 ;
      RECT  1.15 0.79 1.25 1.21 ;
      RECT  1.15 1.21 1.71 1.3 ;
  END
END SEN_ND4B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4B_2
#      Description : "4-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4B_2
  CLASS CORE ;
  FOREIGN SEN_ND4B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.66 3.05 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0948 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.985 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.05 1.41 0.18 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.57 1.42 0.7 1.75 ;
      RECT  1.145 1.425 1.305 1.75 ;
      RECT  1.845 1.42 1.975 1.75 ;
      RECT  2.44 1.21 2.56 1.75 ;
      RECT  2.98 1.21 3.1 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.31 0.05 0.44 0.385 ;
      RECT  2.515 0.05 2.63 0.39 ;
      RECT  3.025 0.05 3.145 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.575 2.205 0.665 ;
      RECT  1.95 0.665 2.05 1.11 ;
      RECT  1.95 1.11 2.285 1.21 ;
      RECT  0.26 1.21 2.285 1.33 ;
    END
    ANTENNADIFFAREA 0.544 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.85 0.14 1.645 0.23 ;
      RECT  0.85 0.23 0.94 0.345 ;
      RECT  1.555 0.23 1.645 0.345 ;
      RECT  1.255 0.32 1.425 0.41 ;
      RECT  1.335 0.41 1.425 0.485 ;
      RECT  1.335 0.485 1.82 0.575 ;
      RECT  1.73 0.395 2.425 0.485 ;
      RECT  2.335 0.485 2.425 0.665 ;
      RECT  0.055 0.33 0.175 0.49 ;
      RECT  0.055 0.49 1.2 0.58 ;
      RECT  1.11 0.58 1.2 0.69 ;
      RECT  2.725 0.44 2.91 0.56 ;
      RECT  2.725 0.56 2.84 0.795 ;
      RECT  2.175 0.795 2.84 0.895 ;
      RECT  2.725 0.895 2.84 1.42 ;
  END
END SEN_ND4B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4B_4
#      Description : "4-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4B_4
  CLASS CORE ;
  FOREIGN SEN_ND4B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.03 0.71 5.65 0.895 ;
      RECT  5.55 0.895 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1893 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.895 ;
      RECT  2.55 0.895 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.895 ;
      RECT  1.35 0.895 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.895 ;
      RECT  0.35 0.895 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.18 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.57 1.42 0.7 1.75 ;
      RECT  1.09 1.42 1.22 1.75 ;
      RECT  1.61 1.42 1.74 1.75 ;
      RECT  2.235 1.425 2.365 1.75 ;
      RECT  2.835 1.42 2.965 1.75 ;
      RECT  3.38 1.425 3.51 1.75 ;
      RECT  3.96 1.415 4.09 1.75 ;
      RECT  4.545 1.21 4.665 1.75 ;
      RECT  5.14 1.44 5.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  5.1 0.05 5.23 0.355 ;
      RECT  0.31 0.05 0.44 0.385 ;
      RECT  0.83 0.05 0.96 0.385 ;
      RECT  5.62 0.05 5.74 0.39 ;
      RECT  4.595 0.05 4.69 0.63 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.51 4.285 0.69 ;
      RECT  3.75 0.69 3.85 1.11 ;
      RECT  3.75 1.11 4.355 1.21 ;
      RECT  0.26 1.21 4.355 1.29 ;
      RECT  0.26 1.29 3.91 1.33 ;
    END
    ANTENNADIFFAREA 1.088 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.965 0.14 2.65 0.215 ;
      RECT  1.3 0.215 3.245 0.23 ;
      RECT  1.3 0.23 2.055 0.305 ;
      RECT  2.555 0.23 3.245 0.305 ;
      RECT  3.375 0.19 4.505 0.32 ;
      RECT  4.405 0.32 4.505 0.39 ;
      RECT  3.375 0.32 3.465 0.4 ;
      RECT  2.27 0.32 2.465 0.4 ;
      RECT  2.27 0.4 3.465 0.41 ;
      RECT  2.375 0.41 3.465 0.49 ;
      RECT  0.055 0.33 0.175 0.475 ;
      RECT  0.055 0.475 2.18 0.56 ;
      RECT  0.055 0.56 2.31 0.595 ;
      RECT  2.08 0.595 2.31 0.65 ;
      RECT  4.805 0.445 5.51 0.56 ;
      RECT  4.805 0.56 4.92 0.795 ;
      RECT  3.96 0.795 4.92 0.895 ;
      RECT  4.805 0.895 4.92 1.23 ;
      RECT  4.805 1.23 5.615 1.35 ;
  END
END SEN_ND4B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_ND4B_8
#      Description : "4-Input NAND (A inverted input)"
#      Equation    : X=!(!A&B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_ND4B_8
  CLASS CORE ;
  FOREIGN SEN_ND4B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.51 0.925 ;
      RECT  0.15 0.925 0.25 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 0.89 ;
      RECT  4.55 0.89 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4392 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.05 0.89 ;
      RECT  3.15 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4392 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 0.895 ;
      RECT  0.95 0.895 2.13 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4392 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.445 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  0.845 1.185 0.965 1.75 ;
      RECT  1.365 1.445 1.485 1.75 ;
      RECT  1.885 1.445 2.005 1.75 ;
      RECT  2.405 1.445 2.525 1.75 ;
      RECT  2.925 1.445 3.045 1.75 ;
      RECT  3.445 1.445 3.565 1.75 ;
      RECT  3.965 1.445 4.085 1.75 ;
      RECT  4.485 1.445 4.605 1.75 ;
      RECT  5.005 1.445 5.125 1.75 ;
      RECT  5.525 1.445 5.645 1.75 ;
      RECT  6.045 1.445 6.165 1.75 ;
      RECT  6.565 1.445 6.685 1.75 ;
      RECT  7.085 1.44 7.205 1.75 ;
      RECT  7.605 1.44 7.725 1.75 ;
      RECT  8.15 1.21 8.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  1.365 0.05 1.485 0.375 ;
      RECT  0.325 0.05 0.445 0.395 ;
      RECT  1.885 0.05 2.005 0.545 ;
      RECT  2.405 0.05 2.525 0.545 ;
      RECT  0.845 0.05 0.965 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.145 0.31 8.265 0.51 ;
      RECT  6.55 0.51 8.265 0.69 ;
      RECT  7.75 0.69 8.05 1.18 ;
      RECT  6.75 0.69 6.93 1.185 ;
      RECT  7.295 1.18 8.05 1.35 ;
      RECT  1.105 1.185 6.93 1.355 ;
    END
    ANTENNADIFFAREA 1.815 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.87 0.17 6.195 0.34 ;
      RECT  6.285 0.19 7.985 0.37 ;
      RECT  6.285 0.37 6.455 0.485 ;
      RECT  4.745 0.485 6.455 0.655 ;
      RECT  0.065 0.345 0.185 0.49 ;
      RECT  0.065 0.49 0.73 0.62 ;
      RECT  0.63 0.62 0.73 1.225 ;
      RECT  0.065 1.225 0.73 1.345 ;
      RECT  0.065 1.345 0.185 1.485 ;
      RECT  2.64 0.44 4.395 0.61 ;
      RECT  2.64 0.61 2.81 0.635 ;
      RECT  1.055 0.465 1.785 0.6 ;
      RECT  1.645 0.6 1.785 0.635 ;
      RECT  1.645 0.635 2.81 0.805 ;
      RECT  7.02 0.86 7.66 1.09 ;
      RECT  7.02 1.09 7.15 1.29 ;
      LAYER M2 ;
      RECT  0.59 1.15 7.16 1.25 ;
      LAYER V1 ;
      RECT  0.63 1.15 0.73 1.25 ;
      RECT  7.02 1.15 7.12 1.25 ;
  END
END SEN_ND4B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_0P5
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_0P5
  CLASS CORE ;
  FOREIGN SEN_NR2_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.205 0.39 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.2 0.45 1.44 ;
      RECT  0.35 1.44 0.745 1.56 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
END SEN_NR2_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_1
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_1
  CLASS CORE ;
  FOREIGN SEN_NR2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.205 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.205 0.39 ;
      RECT  0.595 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 1.44 ;
      RECT  0.35 1.44 0.745 1.56 ;
    END
    ANTENNADIFFAREA 0.199 ;
  END X
END SEN_NR2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_2
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_2
  CLASS CORE ;
  FOREIGN SEN_NR2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.935 1.41 1.065 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.635 0.05 0.765 0.385 ;
      RECT  0.08 0.05 0.2 0.59 ;
      RECT  1.2 0.05 1.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.31 0.46 0.5 ;
      RECT  0.34 0.5 1.06 0.59 ;
      RECT  0.94 0.31 1.06 0.5 ;
      RECT  0.55 0.59 0.65 1.0 ;
      RECT  0.35 1.0 0.65 1.09 ;
      RECT  0.35 1.09 0.45 1.3 ;
    END
    ANTENNADIFFAREA 0.308 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.64 1.21 1.345 1.31 ;
      RECT  0.64 1.31 0.76 1.49 ;
      RECT  0.08 1.41 0.2 1.49 ;
      RECT  0.08 1.49 0.76 1.61 ;
  END
END SEN_NR2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_3
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_3
  CLASS CORE ;
  FOREIGN SEN_NR2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.09 1.41 1.22 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.615 1.21 1.735 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.31 0.05 0.44 0.39 ;
      RECT  0.83 0.05 0.96 0.39 ;
      RECT  1.35 0.05 1.48 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.055 0.19 0.175 0.48 ;
      RECT  0.055 0.48 1.735 0.59 ;
      RECT  1.615 0.37 1.735 0.48 ;
      RECT  0.75 0.59 0.85 1.0 ;
      RECT  0.55 1.0 0.85 1.09 ;
      RECT  0.55 1.09 0.695 1.21 ;
      RECT  0.055 1.21 0.695 1.3 ;
      RECT  0.055 1.3 0.175 1.61 ;
    END
    ANTENNADIFFAREA 0.522 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.835 1.21 1.5 1.32 ;
      RECT  0.835 1.32 0.955 1.41 ;
      RECT  0.29 1.41 0.955 1.53 ;
  END
END SEN_NR2_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_4
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_4
  CLASS CORE ;
  FOREIGN SEN_NR2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.5 2.25 0.71 ;
      RECT  1.55 0.71 2.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.41 1.21 1.54 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.935 1.21 2.065 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.15 0.05 1.28 0.385 ;
      RECT  1.675 0.05 1.805 0.385 ;
      RECT  0.605 0.05 0.735 0.39 ;
      RECT  2.205 0.05 2.335 0.39 ;
      RECT  0.08 0.05 0.2 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.94 0.31 2.06 0.48 ;
      RECT  0.325 0.48 2.06 0.59 ;
      RECT  0.95 0.59 1.05 1.11 ;
      RECT  0.35 1.11 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.624 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.15 1.01 2.32 1.12 ;
      RECT  2.2 1.12 2.32 1.23 ;
      RECT  1.15 1.12 1.28 1.44 ;
      RECT  0.06 1.44 1.28 1.56 ;
  END
END SEN_NR2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_6
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_6
  CLASS CORE ;
  FOREIGN SEN_NR2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 1.195 0.9 ;
      RECT  0.15 0.9 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3852 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 0.71 ;
      RECT  2.15 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3852 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.9 1.21 2.02 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  2.42 1.21 2.54 1.75 ;
      RECT  2.94 1.21 3.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.595 0.05 0.725 0.39 ;
      RECT  1.115 0.05 1.245 0.39 ;
      RECT  1.635 0.05 1.765 0.39 ;
      RECT  2.155 0.05 2.285 0.39 ;
      RECT  2.675 0.05 2.805 0.39 ;
      RECT  3.205 0.05 3.335 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.94 0.31 3.06 0.48 ;
      RECT  0.315 0.48 3.06 0.59 ;
      RECT  1.33 0.59 2.05 0.69 ;
      RECT  1.33 0.69 1.46 1.11 ;
      RECT  0.34 1.11 1.5 1.29 ;
    END
    ANTENNADIFFAREA 0.924 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.64 1.01 3.32 1.12 ;
      RECT  3.2 1.12 3.32 1.23 ;
      RECT  1.64 1.12 1.76 1.44 ;
      RECT  0.08 1.34 0.2 1.44 ;
      RECT  0.08 1.44 1.76 1.56 ;
  END
END SEN_NR2_6
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_8
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_8
  CLASS CORE ;
  FOREIGN SEN_NR2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 1.68 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5136 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.5 4.45 0.71 ;
      RECT  2.95 0.71 4.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5136 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.46 1.21 2.58 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  2.99 1.21 3.11 1.75 ;
      RECT  3.545 1.21 3.665 1.75 ;
      RECT  4.115 1.21 4.235 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.615 0.05 0.745 0.39 ;
      RECT  1.155 0.05 1.285 0.39 ;
      RECT  1.675 0.05 1.805 0.39 ;
      RECT  2.195 0.05 2.325 0.39 ;
      RECT  2.725 0.05 2.855 0.39 ;
      RECT  3.28 0.05 3.41 0.39 ;
      RECT  3.85 0.05 3.98 0.39 ;
      RECT  4.405 0.05 4.535 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.31 0.46 0.48 ;
      RECT  0.34 0.48 4.26 0.59 ;
      RECT  2.475 0.475 2.565 0.48 ;
      RECT  4.14 0.31 4.26 0.48 ;
      RECT  1.89 0.59 2.85 0.69 ;
      RECT  1.89 0.69 2.06 1.11 ;
      RECT  0.34 1.11 2.06 1.29 ;
    END
    ANTENNADIFFAREA 1.232 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.195 1.01 4.52 1.12 ;
      RECT  4.4 1.12 4.52 1.23 ;
      RECT  2.195 1.12 2.325 1.44 ;
      RECT  0.08 1.34 0.2 1.44 ;
      RECT  0.08 1.44 2.325 1.56 ;
  END
END SEN_NR2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_16
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_16
  CLASS CORE ;
  FOREIGN SEN_NR2_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.67 8.05 1.09 ;
      RECT  6.75 0.7 6.85 1.12 ;
      RECT  5.72 0.78 5.82 1.2 ;
      RECT  4.72 0.8 4.82 1.22 ;
      RECT  3.75 0.8 3.85 1.22 ;
      RECT  2.75 0.78 2.85 1.2 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 8.09 1.05 ;
      LAYER V1 ;
      RECT  7.95 0.95 8.05 1.05 ;
      RECT  6.75 0.95 6.85 1.05 ;
      RECT  5.72 0.95 5.82 1.05 ;
      RECT  4.72 0.95 4.82 1.05 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.981 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.71 8.45 0.89 ;
      RECT  8.15 0.89 8.25 1.455 ;
      RECT  7.15 0.71 7.65 0.89 ;
      RECT  7.15 0.89 7.25 1.455 ;
      RECT  7.55 0.89 7.65 1.455 ;
      RECT  6.12 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.455 ;
      RECT  6.12 0.89 6.22 1.505 ;
      RECT  6.55 1.455 7.25 1.545 ;
      RECT  7.55 1.455 8.25 1.545 ;
      RECT  5.1 0.8 5.585 0.905 ;
      RECT  5.485 0.905 5.585 1.505 ;
      RECT  5.1 0.905 5.19 1.525 ;
      RECT  5.485 1.505 6.22 1.595 ;
      RECT  3.945 0.835 4.625 0.935 ;
      RECT  3.945 0.935 4.05 1.525 ;
      RECT  4.52 0.935 4.625 1.525 ;
      RECT  2.95 0.8 3.47 0.9 ;
      RECT  2.95 0.9 3.05 1.505 ;
      RECT  3.38 0.9 3.47 1.525 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.505 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.505 3.05 1.595 ;
      RECT  3.38 1.525 4.05 1.615 ;
      RECT  4.52 1.525 5.19 1.615 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.981 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  1.12 1.185 1.225 1.75 ;
      RECT  2.145 1.185 2.26 1.75 ;
      RECT  3.185 1.23 3.29 1.75 ;
      RECT  4.225 1.18 4.345 1.75 ;
      RECT  5.28 1.18 5.385 1.75 ;
      RECT  6.31 1.185 6.425 1.75 ;
      RECT  7.345 1.175 7.46 1.75 ;
      RECT  8.385 1.21 8.505 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  3.68 0.05 3.865 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.72 0.05 4.89 0.305 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  5.265 0.05 5.385 0.35 ;
      RECT  5.785 0.05 5.905 0.35 ;
      RECT  6.305 0.05 6.425 0.35 ;
      RECT  6.825 0.05 6.945 0.35 ;
      RECT  7.345 0.05 7.465 0.35 ;
      RECT  7.865 0.05 7.985 0.35 ;
      RECT  0.54 0.05 0.66 0.58 ;
      RECT  8.385 0.05 8.505 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.395 5.01 0.44 ;
      RECT  0.75 0.44 8.295 0.56 ;
      RECT  0.75 0.56 7.85 0.57 ;
      RECT  1.75 0.57 7.05 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  7.75 0.57 7.85 1.24 ;
      RECT  2.55 0.61 6.02 0.69 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  6.95 0.61 7.05 1.24 ;
      RECT  3.56 0.69 5.01 0.71 ;
      RECT  2.55 0.69 2.65 1.29 ;
      RECT  5.92 0.69 6.02 1.29 ;
      RECT  3.56 0.71 3.66 1.31 ;
      RECT  4.91 0.71 5.01 1.31 ;
      RECT  0.54 1.24 0.85 1.36 ;
      RECT  1.565 1.24 1.85 1.36 ;
      RECT  6.76 1.24 7.05 1.36 ;
      RECT  7.75 1.24 8.05 1.36 ;
      RECT  2.55 1.29 2.835 1.41 ;
      RECT  5.725 1.29 6.02 1.41 ;
      RECT  3.56 1.31 3.855 1.43 ;
      RECT  4.72 1.31 5.01 1.43 ;
    END
    ANTENNADIFFAREA 2.31 ;
  END X
END SEN_NR2_16
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_8
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_8
  CLASS CORE ;
  FOREIGN SEN_NR2_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.67 3.85 1.09 ;
      RECT  2.75 0.67 2.85 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 3.89 1.05 ;
      LAYER V1 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3717 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.945 0.71 4.25 0.89 ;
      RECT  3.945 0.89 4.05 1.455 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  2.95 0.89 3.05 1.455 ;
      RECT  3.38 0.89 3.47 1.455 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.455 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.455 3.05 1.545 ;
      RECT  3.38 1.455 4.05 1.545 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3717 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  1.12 1.165 1.225 1.75 ;
      RECT  2.145 1.165 2.26 1.75 ;
      RECT  3.185 1.16 3.29 1.75 ;
      RECT  4.215 1.41 4.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  1.08 0.05 1.2 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.69 0.05 2.81 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.44 3.66 0.57 ;
      RECT  1.75 0.57 2.65 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  3.56 0.57 3.66 1.24 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  2.55 0.61 2.65 1.24 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.57 1.24 1.85 1.36 ;
      RECT  2.55 1.24 2.84 1.36 ;
      RECT  3.56 1.24 3.85 1.36 ;
    END
    ANTENNADIFFAREA 0.762 ;
  END X
END SEN_NR2_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_12
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_12
  CLASS CORE ;
  FOREIGN SEN_NR2_G_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.84 0.67 5.94 1.09 ;
      RECT  4.84 0.67 4.94 1.09 ;
      RECT  3.64 0.78 3.74 1.2 ;
      RECT  2.75 0.78 2.85 1.2 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 5.98 1.05 ;
      LAYER V1 ;
      RECT  5.84 0.95 5.94 1.05 ;
      RECT  4.84 0.95 4.94 1.05 ;
      RECT  3.64 0.95 3.74 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.04 0.71 6.34 0.89 ;
      RECT  6.04 0.89 6.14 1.455 ;
      RECT  5.04 0.71 5.55 0.89 ;
      RECT  5.04 0.89 5.14 1.455 ;
      RECT  5.46 0.89 5.55 1.455 ;
      RECT  4.04 0.71 4.54 0.89 ;
      RECT  4.44 0.89 4.54 1.455 ;
      RECT  4.04 0.89 4.14 1.505 ;
      RECT  4.44 1.455 5.14 1.545 ;
      RECT  5.46 1.455 6.14 1.545 ;
      RECT  2.95 0.8 3.54 0.9 ;
      RECT  2.95 0.9 3.05 1.505 ;
      RECT  3.44 0.9 3.54 1.505 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.505 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.505 3.05 1.595 ;
      RECT  3.44 1.505 4.14 1.595 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.12 1.23 1.225 1.75 ;
      RECT  2.145 1.19 2.26 1.75 ;
      RECT  3.185 1.185 3.305 1.75 ;
      RECT  4.23 1.18 4.345 1.75 ;
      RECT  5.265 1.18 5.37 1.75 ;
      RECT  6.32 1.21 6.44 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  4.225 0.05 4.345 0.35 ;
      RECT  4.745 0.05 4.865 0.35 ;
      RECT  5.265 0.05 5.385 0.35 ;
      RECT  5.785 0.05 5.905 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.32 0.05 6.44 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.44 6.215 0.56 ;
      RECT  0.75 0.56 5.74 0.57 ;
      RECT  1.75 0.57 4.74 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  5.64 0.57 5.74 1.24 ;
      RECT  2.55 0.61 3.94 0.69 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  4.64 0.61 4.74 1.24 ;
      RECT  2.55 0.69 2.65 1.29 ;
      RECT  3.84 0.69 3.94 1.29 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.555 1.24 1.85 1.36 ;
      RECT  4.64 1.24 4.925 1.36 ;
      RECT  5.64 1.24 5.94 1.36 ;
      RECT  2.55 1.29 2.84 1.41 ;
      RECT  3.645 1.29 3.94 1.41 ;
    END
    ANTENNADIFFAREA 1.872 ;
  END X
END SEN_NR2_G_12
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_16
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_16
  CLASS CORE ;
  FOREIGN SEN_NR2_G_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.67 8.05 1.09 ;
      RECT  6.75 0.7 6.85 1.12 ;
      RECT  5.72 0.78 5.82 1.2 ;
      RECT  4.72 0.8 4.82 1.22 ;
      RECT  3.75 0.8 3.85 1.22 ;
      RECT  2.75 0.78 2.85 1.2 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 8.09 1.05 ;
      LAYER V1 ;
      RECT  7.95 0.95 8.05 1.05 ;
      RECT  6.75 0.95 6.85 1.05 ;
      RECT  5.72 0.95 5.82 1.05 ;
      RECT  4.72 0.95 4.82 1.05 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.71 8.45 0.89 ;
      RECT  8.15 0.89 8.25 1.455 ;
      RECT  7.15 0.71 7.65 0.89 ;
      RECT  7.15 0.89 7.25 1.455 ;
      RECT  7.55 0.89 7.65 1.455 ;
      RECT  6.12 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.455 ;
      RECT  6.12 0.89 6.22 1.505 ;
      RECT  6.55 1.455 7.25 1.545 ;
      RECT  7.55 1.455 8.25 1.545 ;
      RECT  5.1 0.8 5.585 0.905 ;
      RECT  5.485 0.905 5.585 1.505 ;
      RECT  5.1 0.905 5.19 1.525 ;
      RECT  5.485 1.505 6.22 1.595 ;
      RECT  3.945 0.835 4.625 0.935 ;
      RECT  3.945 0.935 4.05 1.525 ;
      RECT  4.52 0.935 4.625 1.525 ;
      RECT  2.95 0.8 3.47 0.9 ;
      RECT  2.95 0.9 3.05 1.505 ;
      RECT  3.38 0.9 3.47 1.525 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.505 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.505 3.05 1.595 ;
      RECT  3.38 1.525 4.05 1.615 ;
      RECT  4.52 1.525 5.19 1.615 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  1.12 1.18 1.225 1.75 ;
      RECT  2.145 1.165 2.26 1.75 ;
      RECT  3.185 1.175 3.29 1.75 ;
      RECT  4.225 1.18 4.345 1.75 ;
      RECT  5.28 1.185 5.385 1.75 ;
      RECT  6.31 1.18 6.425 1.75 ;
      RECT  7.345 1.165 7.46 1.75 ;
      RECT  8.4 1.21 8.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  3.68 0.05 3.865 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.72 0.05 4.89 0.305 ;
      RECT  0.585 0.05 0.705 0.345 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  5.265 0.05 5.385 0.35 ;
      RECT  5.785 0.05 5.905 0.35 ;
      RECT  6.305 0.05 6.425 0.35 ;
      RECT  6.825 0.05 6.945 0.35 ;
      RECT  7.345 0.05 7.465 0.35 ;
      RECT  7.865 0.05 7.985 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  8.4 0.05 8.52 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.395 5.01 0.44 ;
      RECT  0.275 0.44 8.295 0.56 ;
      RECT  0.75 0.56 7.85 0.57 ;
      RECT  1.75 0.57 7.05 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  7.75 0.57 7.85 1.24 ;
      RECT  2.55 0.61 6.02 0.69 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  6.95 0.61 7.05 1.24 ;
      RECT  3.56 0.69 5.01 0.71 ;
      RECT  2.55 0.69 2.65 1.29 ;
      RECT  5.92 0.69 6.02 1.29 ;
      RECT  3.56 0.71 3.66 1.31 ;
      RECT  4.91 0.71 5.01 1.31 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.56 1.24 1.85 1.36 ;
      RECT  6.76 1.24 7.05 1.36 ;
      RECT  7.75 1.24 8.045 1.36 ;
      RECT  2.55 1.29 2.845 1.41 ;
      RECT  5.69 1.29 6.02 1.41 ;
      RECT  3.56 1.31 3.85 1.43 ;
      RECT  4.72 1.31 5.01 1.43 ;
    END
    ANTENNADIFFAREA 2.496 ;
  END X
END SEN_NR2_G_16
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_24
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_24
  CLASS CORE ;
  FOREIGN SEN_NR2_G_24 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.08 0.51 12.18 0.93 ;
      RECT  10.995 0.51 11.095 0.93 ;
      RECT  9.88 0.51 9.98 0.95 ;
      RECT  8.88 0.51 8.98 0.95 ;
      RECT  7.88 0.51 7.98 0.93 ;
      RECT  6.88 0.46 6.98 0.88 ;
      RECT  5.75 0.46 5.85 0.89 ;
      RECT  4.75 0.51 4.85 0.93 ;
      RECT  3.75 0.51 3.85 0.95 ;
      RECT  2.75 0.51 2.85 0.95 ;
      RECT  1.635 0.51 1.735 0.93 ;
      RECT  0.55 0.51 0.65 0.93 ;
      LAYER M2 ;
      RECT  0.51 0.55 12.22 0.65 ;
      LAYER V1 ;
      RECT  12.08 0.55 12.18 0.65 ;
      RECT  10.995 0.55 11.095 0.65 ;
      RECT  9.88 0.55 9.98 0.65 ;
      RECT  8.88 0.55 8.98 0.65 ;
      RECT  7.88 0.55 7.98 0.65 ;
      RECT  6.88 0.55 6.98 0.65 ;
      RECT  5.75 0.55 5.85 0.65 ;
      RECT  4.75 0.55 4.85 0.65 ;
      RECT  3.75 0.55 3.85 0.65 ;
      RECT  2.75 0.55 2.85 0.65 ;
      RECT  1.635 0.55 1.735 0.65 ;
      RECT  0.55 0.55 0.65 0.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5552 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.48 0.68 12.58 1.12 ;
      RECT  11.48 0.71 11.78 0.89 ;
      RECT  10.28 0.71 10.58 0.89 ;
      RECT  9.28 0.71 9.58 0.89 ;
      RECT  8.28 0.71 8.58 0.89 ;
      RECT  7.23 0.71 7.58 0.85 ;
      RECT  6.15 0.71 6.58 0.86 ;
      RECT  5.15 0.725 5.5 0.895 ;
      RECT  4.15 0.71 4.45 0.89 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.15 0.68 0.25 1.12 ;
      LAYER M2 ;
      RECT  0.11 0.75 12.62 0.85 ;
      LAYER V1 ;
      RECT  12.48 0.75 12.58 0.85 ;
      RECT  11.48 0.75 11.58 0.85 ;
      RECT  11.68 0.75 11.78 0.85 ;
      RECT  10.28 0.75 10.38 0.85 ;
      RECT  10.48 0.75 10.58 0.85 ;
      RECT  9.28 0.75 9.38 0.85 ;
      RECT  9.48 0.75 9.58 0.85 ;
      RECT  8.28 0.75 8.38 0.85 ;
      RECT  8.48 0.75 8.58 0.85 ;
      RECT  7.325 0.75 7.425 0.85 ;
      RECT  6.37 0.75 6.47 0.85 ;
      RECT  5.305 0.75 5.405 0.85 ;
      RECT  4.15 0.75 4.25 0.85 ;
      RECT  4.35 0.75 4.45 0.85 ;
      RECT  3.15 0.75 3.25 0.85 ;
      RECT  3.35 0.75 3.45 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  2.35 0.75 2.45 0.85 ;
      RECT  0.95 0.75 1.05 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  0.15 0.75 0.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.5552 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  1.105 1.455 1.225 1.75 ;
      RECT  2.145 1.415 2.26 1.75 ;
      RECT  3.185 1.415 3.305 1.75 ;
      RECT  4.2 1.495 4.37 1.75 ;
      RECT  5.24 1.495 5.41 1.75 ;
      RECT  6.28 1.495 6.45 1.75 ;
      RECT  7.32 1.495 7.49 1.75 ;
      RECT  8.36 1.495 8.53 1.75 ;
      RECT  9.425 1.415 9.545 1.75 ;
      RECT  10.47 1.415 10.585 1.75 ;
      RECT  11.505 1.455 11.625 1.75 ;
      RECT  12.56 1.21 12.68 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  4.225 0.05 4.345 0.35 ;
      RECT  5.265 0.05 5.385 0.35 ;
      RECT  5.785 0.05 5.905 0.35 ;
      RECT  6.825 0.05 6.945 0.35 ;
      RECT  7.335 0.05 7.465 0.35 ;
      RECT  7.865 0.05 7.985 0.35 ;
      RECT  8.385 0.05 8.505 0.35 ;
      RECT  8.905 0.05 9.025 0.35 ;
      RECT  9.425 0.05 9.545 0.35 ;
      RECT  9.945 0.05 10.065 0.35 ;
      RECT  10.465 0.05 10.585 0.35 ;
      RECT  10.985 0.05 11.105 0.35 ;
      RECT  11.505 0.05 11.625 0.35 ;
      RECT  12.025 0.05 12.145 0.35 ;
      RECT  1.625 0.05 1.745 0.365 ;
      RECT  4.745 0.05 4.865 0.395 ;
      RECT  6.305 0.05 6.425 0.57 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  12.56 0.05 12.68 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  12.28 0.31 12.45 0.49 ;
      RECT  12.28 0.49 12.38 1.11 ;
      RECT  11.22 0.44 11.98 0.56 ;
      RECT  11.88 0.56 11.98 1.11 ;
      RECT  10.08 0.44 10.905 0.56 ;
      RECT  10.08 0.56 10.18 1.04 ;
      RECT  9.68 0.275 9.79 0.44 ;
      RECT  9.08 0.44 9.79 0.56 ;
      RECT  9.08 0.56 9.18 1.04 ;
      RECT  9.08 1.04 10.18 1.085 ;
      RECT  8.08 0.44 8.79 0.56 ;
      RECT  8.08 0.56 8.18 1.085 ;
      RECT  7.08 0.26 7.205 0.44 ;
      RECT  7.08 0.44 7.78 0.56 ;
      RECT  7.68 0.56 7.78 0.97 ;
      RECT  6.515 0.44 6.78 0.56 ;
      RECT  6.68 0.56 6.78 0.97 ;
      RECT  5.95 0.44 6.215 0.56 ;
      RECT  5.95 0.56 6.05 0.97 ;
      RECT  5.95 0.97 7.78 1.0 ;
      RECT  5.525 0.275 5.65 0.44 ;
      RECT  4.95 0.44 5.65 0.56 ;
      RECT  4.95 0.56 5.05 1.0 ;
      RECT  4.95 1.0 7.78 1.085 ;
      RECT  3.94 0.44 4.65 0.56 ;
      RECT  4.55 0.56 4.65 1.085 ;
      RECT  2.94 0.285 3.05 0.44 ;
      RECT  2.94 0.44 3.65 0.56 ;
      RECT  3.55 0.56 3.65 1.04 ;
      RECT  1.83 0.44 2.65 0.56 ;
      RECT  2.55 0.56 2.65 1.04 ;
      RECT  2.55 1.04 3.65 1.085 ;
      RECT  2.55 1.085 10.18 1.11 ;
      RECT  0.75 0.44 1.51 0.56 ;
      RECT  0.75 0.56 0.85 1.11 ;
      RECT  0.3 0.31 0.45 0.485 ;
      RECT  0.35 0.485 0.45 1.11 ;
      RECT  0.35 1.11 12.38 1.29 ;
      RECT  3.7 1.29 9.25 1.39 ;
    END
    ANTENNADIFFAREA 3.744 ;
  END X
END SEN_NR2_G_24
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_6
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_6
  CLASS CORE ;
  FOREIGN SEN_NR2_G_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.67 2.85 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 2.89 1.05 ;
      LAYER V1 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.25 0.89 ;
      RECT  2.95 0.89 3.05 1.455 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.455 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.455 3.05 1.545 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  1.12 1.19 1.225 1.75 ;
      RECT  2.145 1.185 2.26 1.75 ;
      RECT  3.2 1.21 3.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.2 0.05 3.32 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.44 3.095 0.56 ;
      RECT  0.75 0.56 0.85 1.24 ;
      RECT  1.75 0.56 1.85 1.24 ;
      RECT  2.55 0.56 2.65 1.24 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.57 1.24 1.85 1.36 ;
      RECT  2.55 1.24 2.84 1.36 ;
    END
    ANTENNADIFFAREA 0.936 ;
  END X
END SEN_NR2_G_6
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_8
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_8
  CLASS CORE ;
  FOREIGN SEN_NR2_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.67 3.85 1.09 ;
      RECT  2.75 0.67 2.85 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 3.89 1.05 ;
      LAYER V1 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.945 0.71 4.25 0.89 ;
      RECT  3.945 0.89 4.05 1.455 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  2.95 0.89 3.05 1.455 ;
      RECT  3.38 0.89 3.47 1.455 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.455 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.455 3.05 1.545 ;
      RECT  3.38 1.455 4.05 1.545 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  1.12 1.185 1.225 1.75 ;
      RECT  2.145 1.18 2.26 1.75 ;
      RECT  3.185 1.18 3.29 1.75 ;
      RECT  4.215 1.41 4.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  4.215 0.05 4.345 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.44 4.135 0.56 ;
      RECT  0.75 0.56 3.66 0.57 ;
      RECT  1.75 0.57 2.65 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  3.56 0.57 3.66 1.24 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  2.55 0.61 2.65 1.24 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.57 1.24 1.85 1.36 ;
      RECT  2.55 1.24 2.84 1.36 ;
      RECT  3.56 1.24 3.85 1.36 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
END SEN_NR2_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_0P65
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_0P65
  CLASS CORE ;
  FOREIGN SEN_NR2_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0399 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0399 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.065 0.05 0.205 0.39 ;
      RECT  0.595 0.05 0.735 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.23 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.12 ;
  END X
END SEN_NR2_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_0P8
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_0P8
  CLASS CORE ;
  FOREIGN SEN_NR2_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0489 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0489 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.065 0.05 0.205 0.39 ;
      RECT  0.595 0.05 0.735 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.245 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.147 ;
  END X
END SEN_NR2_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_0P5
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_0P5
  CLASS CORE ;
  FOREIGN SEN_NR2_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.027 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.415 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.195 0.385 ;
      RECT  0.605 0.05 0.725 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.21 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.08 ;
  END X
END SEN_NR2_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_0P65
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_0P65
  CLASS CORE ;
  FOREIGN SEN_NR2_S_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.215 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.195 0.385 ;
      RECT  0.605 0.05 0.725 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.21 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.094 ;
  END X
END SEN_NR2_S_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_0P8
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_0P8
  CLASS CORE ;
  FOREIGN SEN_NR2_S_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0378 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.215 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.195 0.385 ;
      RECT  0.605 0.05 0.725 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.21 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.109 ;
  END X
END SEN_NR2_S_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_1
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_1
  CLASS CORE ;
  FOREIGN SEN_NR2_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0465 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0465 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.215 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.195 0.385 ;
      RECT  0.605 0.05 0.725 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.21 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.132 ;
  END X
END SEN_NR2_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_2
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_2
  CLASS CORE ;
  FOREIGN SEN_NR2_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.5 1.25 0.71 ;
      RECT  0.95 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.093 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.093 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.365 1.415 0.505 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.35 0.05 0.47 0.585 ;
      RECT  0.94 0.05 1.06 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.635 0.285 0.85 0.515 ;
      RECT  0.75 0.515 0.85 1.0 ;
      RECT  0.75 1.0 1.04 1.115 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.115 1.21 1.28 1.32 ;
      RECT  0.115 1.32 0.235 1.43 ;
      RECT  1.16 1.32 1.28 1.47 ;
  END
END SEN_NR2_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_3
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_3
  CLASS CORE ;
  FOREIGN SEN_NR2_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1392 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1392 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.565 1.415 0.705 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.835 0.05 0.955 0.385 ;
      RECT  0.28 0.05 0.42 0.39 ;
      RECT  1.37 0.05 1.51 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.27 0.695 0.475 ;
      RECT  0.55 0.475 1.25 0.565 ;
      RECT  1.095 0.275 1.25 0.475 ;
      RECT  1.15 0.565 1.25 1.24 ;
      RECT  1.045 1.24 1.735 1.36 ;
      RECT  1.615 1.36 1.735 1.46 ;
    END
    ANTENNADIFFAREA 0.32 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.265 1.205 0.955 1.325 ;
      RECT  0.835 1.325 0.955 1.45 ;
      RECT  0.835 1.45 1.525 1.57 ;
  END
END SEN_NR2_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_4
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_4
  CLASS CORE ;
  FOREIGN SEN_NR2_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.05 0.71 ;
      RECT  1.55 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.186 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.186 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.46 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.84 1.415 0.98 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.11 0.05 1.23 0.345 ;
      RECT  0.56 0.05 0.68 0.585 ;
      RECT  1.66 0.05 1.78 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.8 0.435 1.54 0.55 ;
      RECT  1.35 0.55 1.45 1.11 ;
      RECT  1.35 1.11 2.06 1.29 ;
    END
    ANTENNADIFFAREA 0.38 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.205 1.23 1.325 ;
      RECT  1.11 1.325 1.23 1.44 ;
      RECT  0.075 1.325 0.19 1.45 ;
      RECT  1.11 1.44 2.27 1.56 ;
      RECT  2.15 1.35 2.27 1.44 ;
  END
END SEN_NR2_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_S_5
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_S_5
  CLASS CORE ;
  FOREIGN SEN_NR2_S_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 0.62 ;
      RECT  1.57 0.62 2.25 0.725 ;
      RECT  2.15 0.725 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2322 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.4 0.62 0.85 0.72 ;
      RECT  0.75 0.72 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2322 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.34 1.415 0.48 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.86 1.415 1.0 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.61 0.05 0.73 0.35 ;
      RECT  1.13 0.05 1.25 0.35 ;
      RECT  1.65 0.05 1.77 0.35 ;
      RECT  0.08 0.05 0.22 0.39 ;
      RECT  2.17 0.05 2.31 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.2 0.47 0.44 ;
      RECT  0.35 0.44 2.05 0.53 ;
      RECT  0.87 0.21 0.99 0.44 ;
      RECT  1.35 0.21 1.51 0.44 ;
      RECT  1.91 0.2 2.05 0.44 ;
      RECT  1.35 0.53 1.465 1.11 ;
      RECT  1.35 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.477 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.09 1.205 1.25 1.325 ;
      RECT  1.13 1.325 1.25 1.44 ;
      RECT  0.09 1.325 0.21 1.46 ;
      RECT  1.13 1.44 2.29 1.56 ;
      RECT  2.17 1.31 2.29 1.44 ;
  END
END SEN_NR2_S_5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_0P5
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_0P5
  CLASS CORE ;
  FOREIGN SEN_NR2_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0492 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.21 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.07 0.05 0.21 0.39 ;
      RECT  0.59 0.05 0.73 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.2 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.093 ;
  END X
END SEN_NR2_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_1
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_1
  CLASS CORE ;
  FOREIGN SEN_NR2_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.31 0.25 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.225 0.48 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.99 0.05 1.13 0.39 ;
      RECT  0.41 0.05 0.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.85 1.24 ;
      RECT  0.75 1.24 1.115 1.36 ;
      RECT  0.995 1.36 1.115 1.47 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.1 1.015 0.66 1.135 ;
      RECT  0.1 1.135 0.22 1.255 ;
      RECT  0.57 1.135 0.66 1.46 ;
      RECT  0.57 1.46 0.885 1.58 ;
  END
END SEN_NR2_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_12
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_12
  CLASS CORE ;
  FOREIGN SEN_NR2_T_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.71 8.25 0.89 ;
      RECT  8.15 0.89 8.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7356 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.225 0.645 4.05 0.75 ;
      RECT  2.95 0.75 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.1676 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.09 1.21 0.21 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  0.63 1.455 0.75 1.75 ;
      RECT  1.15 1.455 1.27 1.75 ;
      RECT  1.67 1.455 1.79 1.75 ;
      RECT  2.185 1.455 2.31 1.75 ;
      RECT  2.705 1.45 2.83 1.75 ;
      RECT  3.23 1.455 3.35 1.75 ;
      RECT  3.75 1.45 3.87 1.75 ;
      RECT  4.27 1.45 4.39 1.75 ;
      RECT  4.79 1.45 4.91 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  3.465 0.05 3.635 0.305 ;
      RECT  3.985 0.05 4.155 0.305 ;
      RECT  4.505 0.05 4.675 0.305 ;
      RECT  5.045 0.05 5.215 0.305 ;
      RECT  5.575 0.05 5.745 0.305 ;
      RECT  0.89 0.05 1.01 0.35 ;
      RECT  1.41 0.05 1.53 0.35 ;
      RECT  1.93 0.05 2.065 0.35 ;
      RECT  2.45 0.05 2.57 0.35 ;
      RECT  2.97 0.05 3.09 0.35 ;
      RECT  7.16 0.05 7.28 0.36 ;
      RECT  7.68 0.05 7.8 0.36 ;
      RECT  6.65 0.05 6.77 0.37 ;
      RECT  6.12 0.05 6.24 0.38 ;
      RECT  0.33 0.05 0.47 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.79 0.255 4.91 0.405 ;
      RECT  4.79 0.405 6.015 0.44 ;
      RECT  3.23 0.27 3.35 0.395 ;
      RECT  3.23 0.395 4.39 0.44 ;
      RECT  3.75 0.26 3.87 0.395 ;
      RECT  4.27 0.275 4.39 0.395 ;
      RECT  0.63 0.26 0.75 0.44 ;
      RECT  0.63 0.44 6.015 0.47 ;
      RECT  1.15 0.265 1.27 0.44 ;
      RECT  1.67 0.27 1.79 0.44 ;
      RECT  2.19 0.26 2.31 0.44 ;
      RECT  2.71 0.265 2.85 0.44 ;
      RECT  0.63 0.47 8.07 0.555 ;
      RECT  7.95 0.285 8.07 0.47 ;
      RECT  4.15 0.555 8.07 0.59 ;
      RECT  4.15 0.59 5.66 0.69 ;
      RECT  5.35 0.69 5.66 1.11 ;
      RECT  5.35 1.11 8.06 1.29 ;
    END
    ANTENNADIFFAREA 1.776 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.43 1.11 5.25 1.19 ;
      RECT  1.87 1.19 5.25 1.24 ;
      RECT  0.315 1.24 5.25 1.36 ;
      RECT  5.0 1.36 5.25 1.4 ;
      RECT  5.0 1.4 7.315 1.44 ;
      RECT  5.0 1.44 8.33 1.58 ;
      RECT  8.2 1.33 8.33 1.44 ;
      RECT  5.0 1.58 6.305 1.64 ;
  END
END SEN_NR2_T_12
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_16
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_16
  CLASS CORE ;
  FOREIGN SEN_NR2_T_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.75 0.71 10.85 0.79 ;
      RECT  8.295 0.79 10.85 0.89 ;
      RECT  10.75 0.89 10.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.981 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.635 5.095 0.74 ;
      RECT  0.15 0.74 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.557 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 11.0 1.85 ;
      RECT  0.61 1.255 0.73 1.75 ;
      RECT  1.13 1.255 1.25 1.75 ;
      RECT  1.65 1.255 1.77 1.75 ;
      RECT  2.185 1.255 2.305 1.75 ;
      RECT  2.705 1.255 2.825 1.75 ;
      RECT  3.225 1.255 3.345 1.75 ;
      RECT  3.74 1.455 3.865 1.75 ;
      RECT  4.26 1.45 4.385 1.75 ;
      RECT  4.785 1.455 4.905 1.75 ;
      RECT  5.305 1.45 5.425 1.75 ;
      RECT  5.825 1.45 5.945 1.75 ;
      RECT  6.345 1.455 6.45 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      RECT  2.94 0.05 3.11 0.305 ;
      RECT  3.46 0.05 3.63 0.305 ;
      RECT  3.98 0.05 4.15 0.305 ;
      RECT  4.5 0.05 4.67 0.305 ;
      RECT  5.02 0.05 5.19 0.305 ;
      RECT  5.535 0.05 5.71 0.305 ;
      RECT  6.06 0.05 6.23 0.305 ;
      RECT  6.58 0.05 6.75 0.305 ;
      RECT  7.11 0.05 7.28 0.305 ;
      RECT  7.63 0.05 7.8 0.305 ;
      RECT  0.35 0.05 0.47 0.345 ;
      RECT  0.87 0.05 0.99 0.345 ;
      RECT  1.39 0.05 1.51 0.345 ;
      RECT  1.925 0.05 2.065 0.345 ;
      RECT  2.445 0.05 2.565 0.35 ;
      RECT  8.705 0.05 8.825 0.36 ;
      RECT  9.225 0.05 9.345 0.36 ;
      RECT  9.745 0.05 9.865 0.36 ;
      RECT  10.265 0.05 10.385 0.36 ;
      RECT  8.185 0.05 8.305 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.705 0.27 2.85 0.395 ;
      RECT  2.705 0.395 6.465 0.405 ;
      RECT  3.225 0.27 3.345 0.395 ;
      RECT  3.745 0.24 3.865 0.395 ;
      RECT  4.265 0.24 4.405 0.395 ;
      RECT  4.785 0.24 4.905 0.395 ;
      RECT  5.305 0.24 5.425 0.395 ;
      RECT  5.825 0.25 5.945 0.395 ;
      RECT  6.345 0.24 6.465 0.395 ;
      RECT  2.705 0.405 8.065 0.44 ;
      RECT  0.065 0.255 0.185 0.44 ;
      RECT  0.065 0.44 8.065 0.47 ;
      RECT  0.61 0.27 0.73 0.44 ;
      RECT  1.13 0.26 1.25 0.44 ;
      RECT  1.65 0.27 1.77 0.44 ;
      RECT  2.185 0.27 2.305 0.44 ;
      RECT  0.065 0.47 10.695 0.545 ;
      RECT  5.35 0.545 10.695 0.59 ;
      RECT  5.35 0.59 8.65 0.69 ;
      RECT  6.85 0.69 7.25 0.91 ;
      RECT  6.85 0.91 8.05 1.005 ;
      RECT  6.85 1.005 10.65 1.11 ;
      RECT  6.95 1.11 10.65 1.18 ;
      RECT  6.95 1.18 8.65 1.25 ;
      LAYER M2 ;
      RECT  3.71 0.35 5.98 0.45 ;
      LAYER V1 ;
      RECT  3.75 0.35 3.85 0.45 ;
      RECT  4.28 0.35 4.38 0.45 ;
      RECT  4.795 0.35 4.895 0.45 ;
      RECT  5.315 0.35 5.415 0.45 ;
      RECT  5.84 0.35 5.94 0.45 ;
    END
    ANTENNADIFFAREA 2.363 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.91 0.975 6.76 1.045 ;
      RECT  0.34 1.045 6.76 1.165 ;
      RECT  3.75 1.165 6.76 1.2 ;
      RECT  0.34 1.165 0.46 1.43 ;
      RECT  3.75 1.2 6.86 1.315 ;
      RECT  6.35 1.315 6.86 1.36 ;
      RECT  6.35 1.36 10.905 1.365 ;
      RECT  10.78 1.245 10.905 1.36 ;
      RECT  6.54 1.365 10.905 1.5 ;
      RECT  6.54 1.5 8.85 1.64 ;
  END
END SEN_NR2_T_16
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_1P5
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_1P5
  CLASS CORE ;
  FOREIGN SEN_NR2_T_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.705 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0912 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1458 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.575 1.455 0.715 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.82 0.05 0.99 0.315 ;
      RECT  1.355 0.05 1.525 0.315 ;
      RECT  0.29 0.05 0.43 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.535 0.405 1.45 0.515 ;
      RECT  1.35 0.515 1.45 1.24 ;
      RECT  1.08 1.24 1.45 1.35 ;
    END
    ANTENNADIFFAREA 0.218 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 1.245 0.965 1.36 ;
      RECT  0.845 1.36 0.965 1.44 ;
      RECT  0.845 1.44 1.485 1.56 ;
      RECT  1.37 1.56 1.485 1.635 ;
  END
END SEN_NR2_T_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_2
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_2
  CLASS CORE ;
  FOREIGN SEN_NR2_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.705 1.45 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.455 0.435 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.835 1.455 0.955 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.095 0.05 1.215 0.36 ;
      RECT  1.615 0.05 1.735 0.36 ;
      RECT  0.55 0.05 0.67 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.785 0.45 1.65 0.56 ;
      RECT  1.55 0.56 1.65 1.11 ;
      RECT  1.35 1.11 1.65 1.29 ;
    END
    ANTENNADIFFAREA 0.288 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 1.245 1.215 1.36 ;
      RECT  1.095 1.36 1.215 1.41 ;
      RECT  0.055 1.36 0.175 1.61 ;
      RECT  1.095 1.41 1.735 1.5 ;
      RECT  1.615 1.5 1.735 1.62 ;
  END
END SEN_NR2_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_3
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_3
  CLASS CORE ;
  FOREIGN SEN_NR2_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1836 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.59 0.63 1.45 0.74 ;
      RECT  1.35 0.74 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2916 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.64 1.45 0.76 1.75 ;
      RECT  1.22 1.455 1.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.64 0.05 0.76 0.345 ;
      RECT  1.22 0.05 1.34 0.345 ;
      RECT  1.86 0.05 1.98 0.345 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  2.39 0.05 2.51 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.335 0.23 0.455 0.435 ;
      RECT  0.335 0.435 2.29 0.525 ;
      RECT  0.93 0.23 1.05 0.435 ;
      RECT  1.55 0.24 1.67 0.435 ;
      RECT  1.75 0.525 2.29 0.555 ;
      RECT  1.75 0.555 1.85 1.235 ;
      RECT  1.75 1.235 2.5 1.355 ;
      RECT  2.38 1.355 2.5 1.46 ;
    END
    ANTENNADIFFAREA 0.5 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 1.24 1.655 1.36 ;
      RECT  1.535 1.36 1.655 1.445 ;
      RECT  1.535 1.445 2.29 1.56 ;
  END
END SEN_NR2_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_4
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_4
  CLASS CORE ;
  FOREIGN SEN_NR2_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.65 0.62 1.65 0.735 ;
      RECT  1.55 0.735 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.585 1.425 0.705 1.75 ;
      RECT  1.105 1.425 1.225 1.75 ;
      RECT  1.625 1.425 1.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.845 0.05 0.965 0.345 ;
      RECT  1.365 0.05 1.485 0.345 ;
      RECT  1.975 0.05 2.095 0.345 ;
      RECT  2.495 0.05 2.615 0.345 ;
      RECT  0.29 0.05 0.43 0.39 ;
      RECT  3.015 0.05 3.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.255 0.705 0.44 ;
      RECT  0.55 0.44 2.9 0.53 ;
      RECT  1.105 0.255 1.25 0.44 ;
      RECT  1.715 0.255 1.85 0.44 ;
      RECT  2.235 0.27 2.355 0.44 ;
      RECT  2.35 0.53 2.9 0.56 ;
      RECT  2.35 0.56 2.45 1.23 ;
      RECT  2.185 1.23 2.925 1.35 ;
    END
    ANTENNADIFFAREA 0.602 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 1.215 2.095 1.335 ;
      RECT  1.975 1.335 2.095 1.44 ;
      RECT  1.975 1.44 3.135 1.56 ;
      RECT  3.015 1.56 3.135 1.64 ;
  END
END SEN_NR2_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_5
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_5
  CLASS CORE ;
  FOREIGN SEN_NR2_T_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.935 0.71 3.45 0.89 ;
      RECT  2.935 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.306 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.655 0.62 1.85 0.735 ;
      RECT  1.75 0.735 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.486 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.345 1.43 0.465 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.87 1.425 0.99 1.75 ;
      RECT  1.39 1.425 1.51 1.75 ;
      RECT  1.955 1.425 2.075 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.61 0.05 0.73 0.345 ;
      RECT  1.13 0.05 1.265 0.345 ;
      RECT  1.65 0.05 1.77 0.345 ;
      RECT  2.26 0.05 2.38 0.345 ;
      RECT  2.78 0.05 2.9 0.345 ;
      RECT  3.3 0.05 3.42 0.35 ;
      RECT  0.07 0.05 0.21 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.24 0.46 0.44 ;
      RECT  0.34 0.44 3.68 0.53 ;
      RECT  0.87 0.24 0.99 0.44 ;
      RECT  1.39 0.24 1.51 0.44 ;
      RECT  1.95 0.24 2.07 0.44 ;
      RECT  2.52 0.28 2.65 0.44 ;
      RECT  3.55 0.3 3.68 0.44 ;
      RECT  1.945 0.53 3.68 0.55 ;
      RECT  2.55 0.55 3.68 0.56 ;
      RECT  2.55 0.56 2.675 1.23 ;
      RECT  2.47 1.23 3.68 1.35 ;
      RECT  3.56 1.35 3.68 1.435 ;
    END
    ANTENNADIFFAREA 0.807 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 1.2 2.38 1.32 ;
      RECT  0.08 1.32 0.2 1.44 ;
      RECT  2.26 1.32 2.38 1.44 ;
      RECT  2.26 1.44 3.47 1.56 ;
  END
END SEN_NR2_T_5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_6
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_6
  CLASS CORE ;
  FOREIGN SEN_NR2_T_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.335 0.71 4.05 0.89 ;
      RECT  3.335 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3672 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.83 0.62 2.25 0.735 ;
      RECT  2.15 0.735 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5832 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.425 0.435 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.835 1.425 0.955 1.75 ;
      RECT  1.355 1.42 1.475 1.75 ;
      RECT  1.875 1.42 1.995 1.75 ;
      RECT  2.395 1.42 2.515 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  2.11 0.05 2.28 0.305 ;
      RECT  0.575 0.05 0.695 0.345 ;
      RECT  1.095 0.05 1.215 0.345 ;
      RECT  1.615 0.05 1.735 0.345 ;
      RECT  2.655 0.05 2.775 0.345 ;
      RECT  3.175 0.05 3.295 0.345 ;
      RECT  3.695 0.05 3.815 0.35 ;
      RECT  4.215 0.05 4.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.875 0.245 1.995 0.42 ;
      RECT  1.875 0.42 2.515 0.44 ;
      RECT  2.395 0.245 2.515 0.42 ;
      RECT  0.315 0.255 0.45 0.44 ;
      RECT  0.315 0.44 4.125 0.53 ;
      RECT  0.835 0.245 0.955 0.44 ;
      RECT  1.35 0.245 1.475 0.44 ;
      RECT  2.375 0.53 4.125 0.56 ;
      RECT  2.375 0.56 3.08 0.57 ;
      RECT  2.95 0.57 3.08 1.23 ;
      RECT  2.875 1.23 4.135 1.35 ;
    END
    ANTENNADIFFAREA 0.881 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 1.2 2.785 1.33 ;
      RECT  2.655 1.33 2.785 1.44 ;
      RECT  0.055 1.33 0.175 1.625 ;
      RECT  2.655 1.44 4.335 1.57 ;
      RECT  4.215 1.57 4.335 1.64 ;
  END
END SEN_NR2_T_6
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_T_8
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_T_8
  CLASS CORE ;
  FOREIGN SEN_NR2_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.92 0.62 2.85 0.735 ;
      RECT  2.75 0.735 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.605 1.455 0.73 1.75 ;
      RECT  1.125 1.45 1.25 1.75 ;
      RECT  1.675 1.455 1.795 1.75 ;
      RECT  2.195 1.45 2.315 1.75 ;
      RECT  2.715 1.45 2.835 1.75 ;
      RECT  3.235 1.45 3.355 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  2.95 0.05 3.12 0.305 ;
      RECT  3.49 0.05 3.66 0.305 ;
      RECT  4.01 0.05 4.18 0.305 ;
      RECT  2.455 0.05 2.575 0.345 ;
      RECT  0.87 0.05 0.99 0.35 ;
      RECT  1.39 0.05 1.51 0.35 ;
      RECT  1.935 0.05 2.055 0.35 ;
      RECT  5.09 0.05 5.21 0.37 ;
      RECT  4.555 0.05 4.675 0.38 ;
      RECT  0.31 0.05 0.45 0.39 ;
      RECT  5.61 0.05 5.73 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.715 0.24 2.85 0.4 ;
      RECT  2.715 0.4 3.355 0.42 ;
      RECT  3.235 0.25 3.355 0.4 ;
      RECT  2.715 0.42 4.45 0.44 ;
      RECT  0.61 0.24 0.73 0.44 ;
      RECT  0.61 0.44 4.45 0.47 ;
      RECT  1.13 0.24 1.25 0.44 ;
      RECT  1.675 0.24 1.795 0.44 ;
      RECT  2.205 0.24 2.315 0.44 ;
      RECT  0.61 0.47 5.52 0.53 ;
      RECT  3.15 0.53 5.52 0.59 ;
      RECT  3.75 0.59 4.05 0.69 ;
      RECT  3.75 0.69 3.92 1.11 ;
      RECT  3.75 1.11 5.46 1.29 ;
    END
    ANTENNADIFFAREA 1.158 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.43 1.19 3.66 1.24 ;
      RECT  0.3 1.24 3.66 1.36 ;
      RECT  3.49 1.36 3.66 1.44 ;
      RECT  3.49 1.44 5.73 1.58 ;
      RECT  5.61 1.355 5.73 1.44 ;
  END
END SEN_NR2_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_0P5
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_0P5
  CLASS CORE ;
  FOREIGN SEN_NR2_G_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.415 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.195 0.385 ;
      RECT  0.605 0.05 0.725 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.17 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
END SEN_NR2_G_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_0P65
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_0P65
  CLASS CORE ;
  FOREIGN SEN_NR2_G_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0423 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0423 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.195 0.39 ;
      RECT  0.605 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.27 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.128 ;
  END X
END SEN_NR2_G_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_0P8
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_0P8
  CLASS CORE ;
  FOREIGN SEN_NR2_G_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0519 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.195 0.39 ;
      RECT  0.605 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.255 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.157 ;
  END X
END SEN_NR2_G_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_1
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_1
  CLASS CORE ;
  FOREIGN SEN_NR2_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.21 0.195 1.75 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      RECT  0.075 0.05 0.195 0.39 ;
      RECT  0.605 0.05 0.725 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.3 0.45 1.31 ;
      RECT  0.35 1.31 0.725 1.49 ;
    END
    ANTENNADIFFAREA 0.196 ;
  END X
END SEN_NR2_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_2
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_2
  CLASS CORE ;
  FOREIGN SEN_NR2_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.705 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.375 1.41 0.495 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.64 0.05 0.76 0.385 ;
      RECT  0.1 0.05 0.22 0.59 ;
      RECT  1.18 0.05 1.3 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.325 0.475 1.075 0.595 ;
      RECT  0.75 0.595 0.85 1.015 ;
      RECT  0.75 1.015 1.06 1.13 ;
    END
    ANTENNADIFFAREA 0.312 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.115 1.22 0.76 1.31 ;
      RECT  0.64 1.31 0.76 1.41 ;
      RECT  0.115 1.31 0.235 1.43 ;
      RECT  0.64 1.41 1.285 1.53 ;
      RECT  1.165 1.53 1.285 1.63 ;
  END
END SEN_NR2_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_3
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_3
  CLASS CORE ;
  FOREIGN SEN_NR2_G_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.575 1.395 0.695 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.575 0.05 0.695 0.385 ;
      RECT  1.095 0.05 1.215 0.385 ;
      RECT  0.055 0.05 0.185 0.39 ;
      RECT  1.615 0.05 1.735 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.265 0.475 1.525 0.595 ;
      RECT  1.15 0.595 1.25 1.235 ;
      RECT  1.045 1.235 1.735 1.355 ;
      RECT  1.615 1.355 1.735 1.49 ;
    END
    ANTENNADIFFAREA 0.504 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.29 1.185 0.955 1.305 ;
      RECT  0.835 1.305 0.955 1.445 ;
      RECT  0.835 1.445 1.525 1.56 ;
  END
END SEN_NR2_G_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2_G_4
#      Description : "2-Input NOR"
#      Equation    : X=!(A1|A2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2_G_4
  CLASS CORE ;
  FOREIGN SEN_NR2_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.4 0.45 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.85 1.4 0.97 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.59 0.05 0.71 0.38 ;
      RECT  1.11 0.05 1.23 0.38 ;
      RECT  1.63 0.05 1.75 0.38 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  2.17 0.05 2.29 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.28 0.47 2.06 0.59 ;
      RECT  1.35 0.59 1.45 1.1 ;
      RECT  1.35 1.1 2.05 1.3 ;
    END
    ANTENNADIFFAREA 0.624 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.19 1.23 1.31 ;
      RECT  0.07 1.31 0.19 1.42 ;
      RECT  1.11 1.31 1.23 1.44 ;
      RECT  1.11 1.44 2.27 1.56 ;
      RECT  2.15 1.34 2.27 1.44 ;
  END
END SEN_NR2_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_1
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_1
  CLASS CORE ;
  FOREIGN SEN_NR2B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0522 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.345 1.59 0.515 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.975 0.05 1.105 0.23 ;
      RECT  0.365 0.05 0.495 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.62 0.32 1.05 0.44 ;
      RECT  0.95 0.44 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.211 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.34 0.19 0.53 ;
      RECT  0.07 0.53 0.86 0.62 ;
      RECT  0.76 0.62 0.86 1.38 ;
      RECT  0.07 1.38 0.86 1.5 ;
      RECT  0.07 1.5 0.19 1.63 ;
  END
END SEN_NR2B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_2
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_2
  CLASS CORE ;
  FOREIGN SEN_NR2B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1044 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  0.58 1.415 0.71 1.75 ;
      RECT  1.545 1.42 1.675 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.285 0.05 1.415 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  0.72 0.05 0.84 0.59 ;
      RECT  1.81 0.05 1.93 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.67 0.5 ;
      RECT  0.95 0.5 1.67 0.59 ;
      RECT  0.95 0.59 1.45 0.69 ;
      RECT  1.35 0.69 1.45 1.0 ;
      RECT  1.005 1.0 1.45 1.12 ;
    END
    ANTENNADIFFAREA 0.308 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.24 0.63 0.36 ;
      RECT  0.54 0.36 0.63 0.78 ;
      RECT  0.54 0.78 1.18 0.89 ;
      RECT  0.54 0.89 0.63 1.195 ;
      RECT  0.3 1.195 0.63 1.315 ;
      RECT  0.77 1.0 0.89 1.21 ;
      RECT  0.77 1.21 1.93 1.33 ;
      RECT  1.81 1.33 1.93 1.43 ;
  END
END SEN_NR2B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_3
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_3
  CLASS CORE ;
  FOREIGN SEN_NR2B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1566 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.95 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.845 1.41 0.975 1.75 ;
      RECT  1.37 1.41 1.5 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  0.845 0.05 0.975 0.36 ;
      RECT  1.37 0.05 1.5 0.39 ;
      RECT  1.89 0.05 2.02 0.39 ;
      RECT  2.41 0.05 2.54 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.09 0.24 1.26 0.36 ;
      RECT  1.15 0.36 1.26 0.51 ;
      RECT  1.15 0.51 2.45 0.6 ;
      RECT  1.55 0.6 2.45 0.69 ;
      RECT  2.35 0.69 2.45 1.11 ;
      RECT  1.895 1.11 2.535 1.29 ;
    END
    ANTENNADIFFAREA 0.498 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.6 0.785 2.24 0.895 ;
      RECT  1.6 0.895 1.69 1.01 ;
      RECT  0.065 0.34 0.185 0.45 ;
      RECT  0.065 0.45 0.85 0.57 ;
      RECT  0.75 0.57 0.85 1.01 ;
      RECT  0.75 1.01 1.69 1.1 ;
      RECT  0.75 1.1 0.85 1.21 ;
      RECT  0.065 1.21 0.85 1.31 ;
      RECT  0.065 1.31 0.185 1.43 ;
      RECT  1.06 1.195 1.755 1.315 ;
      RECT  1.635 1.315 1.755 1.44 ;
      RECT  1.635 1.44 2.33 1.56 ;
  END
END SEN_NR2B_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_4
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_4
  CLASS CORE ;
  FOREIGN SEN_NR2B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2088 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.585 1.41 0.715 1.75 ;
      RECT  1.105 1.41 1.235 1.75 ;
      RECT  2.62 1.41 2.75 1.75 ;
      RECT  3.14 1.41 3.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.585 0.05 0.715 0.36 ;
      RECT  1.84 0.05 1.97 0.39 ;
      RECT  2.36 0.05 2.49 0.39 ;
      RECT  2.88 0.05 3.01 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  1.215 0.05 1.335 0.59 ;
      RECT  3.405 0.05 3.525 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.145 0.31 3.265 0.51 ;
      RECT  1.55 0.51 3.265 0.62 ;
      RECT  1.55 0.62 2.65 0.69 ;
      RECT  2.15 0.69 2.25 1.11 ;
      RECT  1.55 1.11 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.616 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.305 0.45 1.045 0.57 ;
      RECT  0.955 0.57 1.045 0.78 ;
      RECT  0.955 0.78 2.04 0.89 ;
      RECT  0.955 0.89 1.045 1.21 ;
      RECT  0.28 1.21 1.045 1.31 ;
      RECT  2.365 1.21 3.525 1.31 ;
      RECT  3.405 1.31 3.525 1.43 ;
      RECT  2.365 1.31 2.485 1.44 ;
      RECT  1.325 0.99 1.445 1.44 ;
      RECT  1.325 1.44 2.485 1.56 ;
  END
END SEN_NR2B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1DG_12
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1DG_12
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1DG_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.71 7.05 0.89 ;
      RECT  6.95 0.89 7.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.84 0.67 5.94 1.09 ;
      RECT  4.84 0.67 4.94 1.09 ;
      RECT  3.64 0.78 3.74 1.2 ;
      RECT  2.75 0.78 2.85 1.2 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 5.98 1.05 ;
      LAYER V1 ;
      RECT  5.84 0.95 5.94 1.05 ;
      RECT  4.84 0.95 4.94 1.05 ;
      RECT  3.64 0.95 3.74 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.4 1.85 ;
      RECT  1.12 1.2 1.225 1.75 ;
      RECT  2.145 1.2 2.26 1.75 ;
      RECT  3.185 1.2 3.305 1.75 ;
      RECT  4.23 1.2 4.345 1.75 ;
      RECT  5.265 1.2 5.37 1.75 ;
      RECT  6.34 1.455 6.46 1.75 ;
      RECT  6.885 1.455 7.005 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      RECT  6.305 0.05 6.425 0.345 ;
      RECT  6.885 0.05 7.005 0.345 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  4.225 0.05 4.345 0.35 ;
      RECT  4.745 0.05 4.865 0.35 ;
      RECT  5.265 0.05 5.385 0.35 ;
      RECT  5.785 0.05 5.905 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.3 0.44 6.215 0.56 ;
      RECT  0.75 0.56 5.74 0.57 ;
      RECT  1.75 0.57 4.74 0.6 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  5.64 0.57 5.74 1.24 ;
      RECT  2.55 0.6 3.94 0.69 ;
      RECT  1.75 0.6 1.85 1.24 ;
      RECT  4.64 0.6 4.74 1.24 ;
      RECT  2.55 0.69 2.65 1.29 ;
      RECT  3.84 0.69 3.94 1.29 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.555 1.24 1.85 1.36 ;
      RECT  4.64 1.24 4.92 1.36 ;
      RECT  5.64 1.24 5.96 1.36 ;
      RECT  2.55 1.29 2.84 1.41 ;
      RECT  3.64 1.29 3.94 1.41 ;
    END
    ANTENNADIFFAREA 1.872 ;
  END X
  OBS
      LAYER M1 ;
      RECT  7.145 0.265 7.265 0.44 ;
      RECT  6.35 0.44 7.265 0.56 ;
      RECT  6.35 0.56 6.45 0.73 ;
      RECT  6.15 0.73 6.45 0.84 ;
      RECT  6.15 0.84 6.25 1.24 ;
      RECT  6.15 1.24 7.265 1.36 ;
      RECT  6.15 1.36 6.25 1.455 ;
      RECT  7.14 1.36 7.265 1.51 ;
      RECT  5.04 0.71 5.55 0.89 ;
      RECT  5.04 0.89 5.14 1.455 ;
      RECT  5.46 0.89 5.55 1.455 ;
      RECT  4.04 0.71 4.54 0.89 ;
      RECT  4.44 0.89 4.54 1.455 ;
      RECT  4.04 0.89 4.14 1.505 ;
      RECT  4.44 1.455 5.14 1.545 ;
      RECT  5.46 1.455 6.25 1.545 ;
      RECT  2.95 0.8 3.54 0.9 ;
      RECT  2.95 0.9 3.05 1.505 ;
      RECT  3.44 0.9 3.54 1.505 ;
      RECT  1.95 0.71 2.45 0.9 ;
      RECT  1.95 0.9 2.05 1.455 ;
      RECT  2.35 0.9 2.45 1.505 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.505 3.05 1.595 ;
      RECT  3.44 1.505 4.14 1.595 ;
  END
END SEN_NR2B_V1DG_12
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1DG_16
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1DG_16
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1DG_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.895 0.71 9.25 0.89 ;
      RECT  9.15 0.89 9.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.67 8.05 1.09 ;
      RECT  6.75 0.7 6.85 1.12 ;
      RECT  5.72 0.78 5.82 1.2 ;
      RECT  4.72 0.8 4.82 1.22 ;
      RECT  3.75 0.8 3.85 1.22 ;
      RECT  2.75 0.78 2.85 1.2 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 8.09 1.05 ;
      LAYER V1 ;
      RECT  7.95 0.95 8.05 1.05 ;
      RECT  6.75 0.95 6.85 1.05 ;
      RECT  5.72 0.95 5.82 1.05 ;
      RECT  4.72 0.95 4.82 1.05 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  1.12 1.2 1.225 1.75 ;
      RECT  2.145 1.2 2.26 1.75 ;
      RECT  3.185 1.2 3.29 1.75 ;
      RECT  4.225 1.2 4.345 1.75 ;
      RECT  5.28 1.2 5.385 1.75 ;
      RECT  6.31 1.2 6.425 1.75 ;
      RECT  7.345 1.2 7.46 1.75 ;
      RECT  8.385 1.2 8.505 1.75 ;
      RECT  8.905 1.455 9.025 1.75 ;
      RECT  9.415 1.41 9.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  3.68 0.05 3.865 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.72 0.05 4.89 0.305 ;
      RECT  0.585 0.05 0.705 0.345 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  5.265 0.05 5.385 0.35 ;
      RECT  5.785 0.05 5.905 0.35 ;
      RECT  6.305 0.05 6.425 0.35 ;
      RECT  6.825 0.05 6.945 0.35 ;
      RECT  7.345 0.05 7.465 0.35 ;
      RECT  7.865 0.05 7.985 0.35 ;
      RECT  8.905 0.05 9.025 0.35 ;
      RECT  9.415 0.05 9.545 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  8.385 0.05 8.505 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.395 5.01 0.44 ;
      RECT  0.275 0.44 8.295 0.56 ;
      RECT  0.75 0.56 7.85 0.57 ;
      RECT  1.75 0.57 7.05 0.6 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  7.75 0.57 7.85 1.24 ;
      RECT  2.55 0.6 6.02 0.69 ;
      RECT  1.75 0.6 1.85 1.24 ;
      RECT  6.95 0.6 7.05 1.24 ;
      RECT  3.56 0.69 5.01 0.71 ;
      RECT  2.55 0.69 2.65 1.29 ;
      RECT  5.92 0.69 6.02 1.29 ;
      RECT  3.56 0.71 3.66 1.31 ;
      RECT  4.91 0.71 5.01 1.31 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.565 1.24 1.85 1.36 ;
      RECT  6.755 1.24 7.05 1.36 ;
      RECT  7.75 1.24 8.035 1.36 ;
      RECT  2.55 1.29 2.835 1.41 ;
      RECT  5.72 1.29 6.02 1.41 ;
      RECT  3.56 1.31 3.85 1.43 ;
      RECT  4.72 1.31 5.01 1.43 ;
    END
    ANTENNADIFFAREA 2.496 ;
  END X
  OBS
      LAYER M1 ;
      RECT  8.61 0.44 9.335 0.56 ;
      RECT  8.61 0.56 8.7 0.785 ;
      RECT  8.15 0.785 8.7 0.895 ;
      RECT  8.61 0.895 8.7 1.24 ;
      RECT  8.15 0.895 8.25 1.455 ;
      RECT  8.61 1.24 9.31 1.36 ;
      RECT  7.15 0.71 7.65 0.89 ;
      RECT  7.15 0.89 7.25 1.455 ;
      RECT  7.55 0.89 7.65 1.455 ;
      RECT  6.12 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.455 ;
      RECT  6.12 0.89 6.22 1.505 ;
      RECT  6.55 1.455 7.25 1.545 ;
      RECT  7.55 1.455 8.25 1.545 ;
      RECT  5.1 0.8 5.585 0.905 ;
      RECT  5.485 0.905 5.585 1.505 ;
      RECT  5.1 0.905 5.19 1.525 ;
      RECT  5.485 1.505 6.22 1.595 ;
      RECT  3.945 0.82 4.625 0.93 ;
      RECT  3.945 0.93 4.05 1.525 ;
      RECT  4.52 0.93 4.625 1.525 ;
      RECT  2.95 0.8 3.47 0.9 ;
      RECT  2.95 0.9 3.05 1.505 ;
      RECT  3.38 0.9 3.47 1.525 ;
      RECT  1.95 0.71 2.45 0.895 ;
      RECT  1.95 0.895 2.05 1.455 ;
      RECT  2.35 0.895 2.45 1.505 ;
      RECT  0.94 0.725 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.505 3.05 1.595 ;
      RECT  3.38 1.525 4.05 1.615 ;
      RECT  4.52 1.525 5.19 1.615 ;
  END
END SEN_NR2B_V1DG_16
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1DG_6
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1DG_6
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1DG_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.705 3.65 0.91 ;
      RECT  3.55 0.91 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.67 2.85 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 2.89 1.05 ;
      LAYER V1 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  1.105 1.23 1.225 1.75 ;
      RECT  2.145 1.23 2.265 1.75 ;
      RECT  3.195 1.42 3.315 1.75 ;
      RECT  3.76 1.21 3.88 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  3.195 0.05 3.315 0.345 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.76 0.05 3.88 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.44 3.07 0.56 ;
      RECT  0.75 0.56 0.85 1.31 ;
      RECT  1.75 0.56 1.85 1.31 ;
      RECT  2.55 0.56 2.65 1.31 ;
      RECT  0.55 1.31 0.85 1.49 ;
      RECT  1.55 1.31 1.85 1.49 ;
      RECT  2.55 1.31 2.85 1.49 ;
    END
    ANTENNADIFFAREA 0.94 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.16 0.435 3.63 0.555 ;
      RECT  3.16 0.555 3.26 1.18 ;
      RECT  3.16 1.18 3.655 1.3 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  0.15 0.69 0.28 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.75 3.3 0.85 ;
      LAYER V1 ;
      RECT  0.15 0.75 0.25 0.85 ;
      RECT  0.95 0.75 1.05 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  2.35 0.75 2.45 0.85 ;
      RECT  3.16 0.75 3.26 0.85 ;
  END
END SEN_NR2B_V1DG_6
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1DG_8
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1DG_8
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.85 0.89 ;
      RECT  4.55 0.89 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.67 3.85 1.09 ;
      RECT  2.75 0.67 2.85 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 3.89 1.05 ;
      LAYER V1 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.12 1.19 1.225 1.75 ;
      RECT  2.145 1.195 2.26 1.75 ;
      RECT  3.185 1.18 3.29 1.75 ;
      RECT  4.265 1.43 4.385 1.75 ;
      RECT  4.8 1.21 4.92 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  4.265 0.05 4.385 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  4.8 0.05 4.92 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.44 4.085 0.56 ;
      RECT  0.75 0.56 3.66 0.57 ;
      RECT  3.95 0.56 4.085 0.7 ;
      RECT  1.75 0.57 2.65 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  3.56 0.57 3.66 1.24 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  2.55 0.61 2.65 1.24 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.57 1.24 1.85 1.36 ;
      RECT  2.55 1.24 2.84 1.36 ;
      RECT  3.56 1.24 3.85 1.36 ;
    END
    ANTENNADIFFAREA 1.268 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.2 0.44 4.695 0.56 ;
      RECT  4.2 0.56 4.3 1.215 ;
      RECT  3.945 1.215 4.695 1.335 ;
      RECT  3.945 1.335 4.05 1.455 ;
      RECT  2.95 0.725 3.47 0.9 ;
      RECT  2.95 0.9 3.05 1.455 ;
      RECT  3.38 0.9 3.47 1.455 ;
      RECT  1.95 0.725 2.45 0.895 ;
      RECT  1.95 0.895 2.05 1.455 ;
      RECT  2.35 0.895 2.45 1.455 ;
      RECT  0.94 0.725 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.185 0.76 0.45 0.885 ;
      RECT  0.35 0.885 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.455 3.05 1.545 ;
      RECT  3.38 1.455 4.05 1.545 ;
  END
END SEN_NR2B_V1DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1_8
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1_8
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.095 0.89 ;
      RECT  4.75 0.89 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.67 3.85 1.09 ;
      RECT  2.75 0.67 2.85 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  0.55 0.67 0.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 3.89 1.05 ;
      LAYER V1 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  1.12 1.195 1.225 1.75 ;
      RECT  2.145 1.2 2.26 1.75 ;
      RECT  3.185 1.2 3.29 1.75 ;
      RECT  4.225 1.2 4.345 1.75 ;
      RECT  4.745 1.45 4.865 1.75 ;
      RECT  5.29 1.21 5.41 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  4.745 0.05 4.865 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.29 0.05 5.41 0.59 ;
      RECT  4.225 0.05 4.345 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.44 4.085 0.56 ;
      RECT  0.75 0.56 3.66 0.57 ;
      RECT  3.95 0.56 4.085 0.69 ;
      RECT  1.75 0.57 2.65 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  3.56 0.57 3.66 1.24 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  2.55 0.61 2.65 1.24 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.56 1.24 1.85 1.36 ;
      RECT  2.55 1.24 2.845 1.36 ;
      RECT  3.56 1.24 3.85 1.36 ;
    END
    ANTENNADIFFAREA 1.152 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.485 0.44 5.175 0.56 ;
      RECT  4.485 0.56 4.605 0.785 ;
      RECT  3.945 0.785 4.605 0.9 ;
      RECT  4.485 0.9 4.605 1.24 ;
      RECT  3.945 0.9 4.05 1.455 ;
      RECT  4.485 1.24 5.175 1.36 ;
      RECT  2.95 0.725 3.47 0.89 ;
      RECT  2.95 0.89 3.05 1.455 ;
      RECT  3.38 0.89 3.47 1.455 ;
      RECT  1.95 0.725 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.455 ;
      RECT  0.94 0.725 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.195 0.78 0.45 0.9 ;
      RECT  0.35 0.9 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.455 3.05 1.545 ;
      RECT  3.38 1.455 4.05 1.545 ;
  END
END SEN_NR2B_V1_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_12
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_12
  CLASS CORE ;
  FOREIGN SEN_NR2B_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.71 7.65 0.89 ;
      RECT  7.55 0.89 7.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3672 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.04 0.71 5.55 0.89 ;
      RECT  5.04 0.89 5.14 1.455 ;
      RECT  5.46 0.89 5.55 1.455 ;
      RECT  4.04 0.71 4.54 0.89 ;
      RECT  4.44 0.89 4.54 1.455 ;
      RECT  4.04 0.89 4.14 1.505 ;
      RECT  4.44 1.455 5.14 1.545 ;
      RECT  5.46 1.455 6.25 1.545 ;
      RECT  6.15 0.71 6.25 1.455 ;
      RECT  2.95 0.8 3.54 0.9 ;
      RECT  2.95 0.9 3.05 1.505 ;
      RECT  3.44 0.9 3.54 1.505 ;
      RECT  1.95 0.71 2.45 0.895 ;
      RECT  1.95 0.895 2.05 1.455 ;
      RECT  2.35 0.895 2.45 1.505 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.925 ;
      RECT  0.35 0.925 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.505 3.05 1.595 ;
      RECT  3.44 1.505 4.14 1.595 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7344 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  1.12 1.2 1.225 1.75 ;
      RECT  2.145 1.2 2.26 1.75 ;
      RECT  3.185 1.2 3.305 1.75 ;
      RECT  4.23 1.2 4.345 1.75 ;
      RECT  5.265 1.2 5.37 1.75 ;
      RECT  6.34 1.455 6.46 1.75 ;
      RECT  6.885 1.455 7.005 1.75 ;
      RECT  7.405 1.455 7.525 1.75 ;
      RECT  7.94 1.21 8.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  6.305 0.05 6.425 0.345 ;
      RECT  6.885 0.05 7.005 0.345 ;
      RECT  7.405 0.05 7.525 0.345 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  4.225 0.05 4.345 0.35 ;
      RECT  4.745 0.05 4.865 0.35 ;
      RECT  5.265 0.05 5.385 0.35 ;
      RECT  5.785 0.05 5.905 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  7.94 0.05 8.06 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.3 0.44 6.215 0.56 ;
      RECT  0.75 0.56 5.74 0.57 ;
      RECT  1.75 0.57 4.74 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  5.64 0.57 5.74 1.24 ;
      RECT  2.55 0.61 3.94 0.69 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  4.64 0.61 4.74 1.24 ;
      RECT  2.55 0.69 2.65 1.29 ;
      RECT  3.84 0.69 3.94 1.29 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.565 1.24 1.85 1.36 ;
      RECT  4.64 1.24 4.915 1.36 ;
      RECT  5.64 1.24 5.94 1.36 ;
      RECT  2.55 1.29 2.835 1.41 ;
      RECT  3.65 1.29 3.94 1.41 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.35 0.44 7.835 0.57 ;
      RECT  6.35 0.57 6.48 1.23 ;
      RECT  6.35 1.23 7.835 1.36 ;
      RECT  0.55 0.67 0.65 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  4.84 0.67 4.94 1.09 ;
      RECT  5.84 0.67 5.94 1.09 ;
      RECT  2.75 0.78 2.85 1.2 ;
      RECT  3.64 0.78 3.74 1.2 ;
      LAYER M2 ;
      RECT  0.51 0.95 6.49 1.05 ;
      LAYER V1 ;
      RECT  0.55 0.95 0.65 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  3.64 0.95 3.74 1.05 ;
      RECT  4.84 0.95 4.94 1.05 ;
      RECT  5.84 0.95 5.94 1.05 ;
      RECT  6.35 0.95 6.45 1.05 ;
  END
END SEN_NR2B_12
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_16
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_16
  CLASS CORE ;
  FOREIGN SEN_NR2B_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.065 0.71 10.05 0.89 ;
      RECT  9.95 0.89 10.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.705 8.45 0.92 ;
      RECT  8.15 0.92 8.25 1.455 ;
      RECT  7.15 0.71 7.65 0.89 ;
      RECT  7.15 0.89 7.25 1.455 ;
      RECT  7.55 0.89 7.65 1.455 ;
      RECT  6.12 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.455 ;
      RECT  6.12 0.89 6.22 1.505 ;
      RECT  6.55 1.455 7.25 1.545 ;
      RECT  7.55 1.455 8.25 1.545 ;
      RECT  5.1 0.8 5.585 0.905 ;
      RECT  5.485 0.905 5.585 1.505 ;
      RECT  5.1 0.905 5.19 1.525 ;
      RECT  5.485 1.505 6.22 1.595 ;
      RECT  3.945 0.82 4.625 0.92 ;
      RECT  3.945 0.92 4.05 1.525 ;
      RECT  4.52 0.92 4.625 1.525 ;
      RECT  2.95 0.8 3.47 0.9 ;
      RECT  2.95 0.9 3.05 1.505 ;
      RECT  3.38 0.9 3.47 1.525 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.505 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.9 ;
      RECT  0.35 0.9 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.505 3.05 1.595 ;
      RECT  3.38 1.525 4.05 1.615 ;
      RECT  4.52 1.525 5.19 1.615 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9792 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 10.8 1.85 ;
      RECT  1.12 1.2 1.225 1.75 ;
      RECT  2.145 1.2 2.26 1.75 ;
      RECT  3.185 1.2 3.29 1.75 ;
      RECT  4.225 1.23 4.345 1.75 ;
      RECT  5.28 1.23 5.385 1.75 ;
      RECT  6.31 1.23 6.425 1.75 ;
      RECT  7.345 1.23 7.46 1.75 ;
      RECT  8.385 1.23 8.505 1.75 ;
      RECT  8.905 1.42 9.025 1.75 ;
      RECT  9.425 1.42 9.545 1.75 ;
      RECT  9.945 1.42 10.065 1.75 ;
      RECT  10.5 1.21 10.62 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      RECT  3.68 0.05 3.865 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.72 0.05 4.89 0.305 ;
      RECT  8.88 0.05 9.05 0.335 ;
      RECT  9.4 0.05 9.57 0.335 ;
      RECT  9.92 0.05 10.09 0.335 ;
      RECT  0.585 0.05 0.705 0.345 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  5.265 0.05 5.385 0.35 ;
      RECT  5.785 0.05 5.905 0.35 ;
      RECT  6.305 0.05 6.425 0.35 ;
      RECT  6.825 0.05 6.945 0.35 ;
      RECT  7.345 0.05 7.465 0.35 ;
      RECT  7.865 0.05 7.985 0.35 ;
      RECT  8.385 0.05 8.505 0.45 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  10.5 0.05 10.62 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.395 5.01 0.44 ;
      RECT  0.275 0.44 8.295 0.56 ;
      RECT  0.75 0.56 7.85 0.57 ;
      RECT  1.75 0.57 7.05 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  7.75 0.57 7.85 1.24 ;
      RECT  2.55 0.61 6.02 0.69 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  6.95 0.61 7.05 1.24 ;
      RECT  3.56 0.69 5.01 0.71 ;
      RECT  2.55 0.69 2.65 1.29 ;
      RECT  5.92 0.69 6.02 1.29 ;
      RECT  3.56 0.71 3.66 1.31 ;
      RECT  4.91 0.71 5.01 1.31 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.56 1.24 1.85 1.36 ;
      RECT  6.8 1.24 7.05 1.36 ;
      RECT  7.75 1.24 8.02 1.36 ;
      RECT  2.55 1.29 2.84 1.41 ;
      RECT  5.72 1.29 6.02 1.41 ;
      RECT  3.56 1.31 3.85 1.43 ;
      RECT  4.72 1.31 5.01 1.43 ;
    END
    ANTENNADIFFAREA 2.304 ;
  END X
  OBS
      LAYER M1 ;
      RECT  8.62 0.44 10.375 0.56 ;
      RECT  8.62 0.56 9.31 0.61 ;
      RECT  8.62 0.61 8.79 1.16 ;
      RECT  8.62 1.16 9.31 1.21 ;
      RECT  8.62 1.21 10.375 1.33 ;
      RECT  0.55 0.67 0.65 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  7.95 0.67 8.05 1.09 ;
      RECT  6.75 0.7 6.85 1.12 ;
      RECT  2.75 0.78 2.85 1.2 ;
      RECT  5.72 0.78 5.82 1.2 ;
      RECT  3.75 0.8 3.85 1.22 ;
      RECT  4.72 0.8 4.82 1.22 ;
      LAYER M2 ;
      RECT  0.51 0.95 8.775 1.05 ;
      LAYER V1 ;
      RECT  0.55 0.95 0.65 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  4.72 0.95 4.82 1.05 ;
      RECT  5.72 0.95 5.82 1.05 ;
      RECT  6.75 0.95 6.85 1.05 ;
      RECT  7.95 0.95 8.05 1.05 ;
      RECT  8.635 0.95 8.735 1.05 ;
  END
END SEN_NR2B_16
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_6
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_6
  CLASS CORE ;
  FOREIGN SEN_NR2B_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.66 0.705 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1836 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.25 0.89 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.15 0.69 0.285 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.75 3.29 0.85 ;
      LAYER V1 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  3.15 0.75 3.25 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  2.35 0.75 2.45 0.85 ;
      RECT  0.95 0.75 1.05 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  0.15 0.75 0.25 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3672 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  1.105 1.2 1.225 1.75 ;
      RECT  2.145 1.2 2.265 1.75 ;
      RECT  3.185 1.22 3.305 1.75 ;
      RECT  3.705 1.45 3.825 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.185 0.05 3.305 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.44 3.095 0.56 ;
      RECT  0.75 0.56 0.85 1.31 ;
      RECT  1.75 0.56 1.85 1.31 ;
      RECT  2.55 0.56 2.65 1.31 ;
      RECT  0.55 1.31 0.85 1.49 ;
      RECT  1.55 1.31 1.85 1.49 ;
      RECT  2.55 1.31 2.85 1.49 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.95 0.31 4.085 0.44 ;
      RECT  3.42 0.44 4.085 0.56 ;
      RECT  3.42 0.56 3.525 1.015 ;
      RECT  2.75 0.67 2.85 1.015 ;
      RECT  2.75 1.015 3.525 1.13 ;
      RECT  3.42 1.13 3.525 1.24 ;
      RECT  3.42 1.24 4.085 1.36 ;
      RECT  3.97 1.36 4.085 1.49 ;
      RECT  0.55 0.67 0.65 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 2.89 1.05 ;
      LAYER V1 ;
      RECT  0.55 0.95 0.65 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
  END
END SEN_NR2B_6
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_8
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_8
  CLASS CORE ;
  FOREIGN SEN_NR2B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.05 0.9 ;
      RECT  4.75 0.9 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.945 0.71 4.25 0.89 ;
      RECT  3.945 0.89 4.05 1.455 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  2.95 0.89 3.05 1.455 ;
      RECT  3.38 0.89 3.47 1.455 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  1.95 0.89 2.05 1.455 ;
      RECT  2.35 0.89 2.45 1.455 ;
      RECT  0.94 0.71 1.45 0.89 ;
      RECT  0.94 0.89 1.03 1.455 ;
      RECT  1.35 0.89 1.45 1.455 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.455 ;
      RECT  0.35 1.455 1.03 1.545 ;
      RECT  1.35 1.455 2.05 1.545 ;
      RECT  2.35 1.455 3.05 1.545 ;
      RECT  3.38 1.455 4.05 1.545 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  1.12 1.2 1.225 1.75 ;
      RECT  2.145 1.195 2.26 1.75 ;
      RECT  3.185 1.2 3.29 1.75 ;
      RECT  4.225 1.17 4.345 1.75 ;
      RECT  4.745 1.45 4.865 1.75 ;
      RECT  5.3 1.21 5.42 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.35 ;
      RECT  2.145 0.05 2.265 0.35 ;
      RECT  2.665 0.05 2.785 0.35 ;
      RECT  3.185 0.05 3.305 0.35 ;
      RECT  3.705 0.05 3.825 0.35 ;
      RECT  4.745 0.05 4.865 0.35 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  5.3 0.05 5.42 0.59 ;
      RECT  4.225 0.05 4.345 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.44 4.135 0.56 ;
      RECT  0.75 0.56 3.66 0.57 ;
      RECT  1.75 0.57 2.65 0.61 ;
      RECT  0.75 0.57 0.85 1.24 ;
      RECT  3.56 0.57 3.66 1.24 ;
      RECT  1.75 0.61 1.85 1.24 ;
      RECT  2.55 0.61 2.65 1.24 ;
      RECT  0.55 1.24 0.85 1.36 ;
      RECT  1.56 1.24 1.85 1.36 ;
      RECT  2.55 1.24 2.84 1.36 ;
      RECT  3.56 1.24 3.85 1.36 ;
    END
    ANTENNADIFFAREA 1.152 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.485 0.44 5.175 0.56 ;
      RECT  4.485 0.56 4.605 1.24 ;
      RECT  4.485 1.24 5.175 1.36 ;
      RECT  0.55 0.67 0.65 1.09 ;
      RECT  1.55 0.67 1.65 1.09 ;
      RECT  2.75 0.67 2.85 1.09 ;
      RECT  3.75 0.67 3.85 1.09 ;
      LAYER M2 ;
      RECT  0.51 0.95 4.635 1.05 ;
      LAYER V1 ;
      RECT  0.55 0.95 0.65 1.05 ;
      RECT  1.55 0.95 1.65 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  3.75 0.95 3.85 1.05 ;
      RECT  4.495 0.95 4.595 1.05 ;
  END
END SEN_NR2B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1DG_1
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1DG_1
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.37 1.41 0.51 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.37 0.05 0.51 0.385 ;
      RECT  0.985 0.05 1.125 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.85 1.31 ;
      RECT  0.75 1.31 1.115 1.49 ;
    END
    ANTENNADIFFAREA 0.212 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.185 0.185 0.485 ;
      RECT  0.065 0.485 0.65 0.575 ;
      RECT  0.55 0.575 0.65 1.21 ;
      RECT  0.065 1.21 0.65 1.3 ;
      RECT  0.065 1.3 0.185 1.6 ;
  END
END SEN_NR2B_V1DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1DG_2
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1DG_2
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.51 0.255 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.835 1.415 0.975 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.095 0.05 1.235 0.385 ;
      RECT  1.615 0.05 1.745 0.385 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  0.585 0.05 0.705 0.615 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.795 0.475 1.65 0.595 ;
      RECT  1.55 0.595 1.65 1.11 ;
      RECT  1.35 1.11 1.65 1.29 ;
    END
    ANTENNADIFFAREA 0.312 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.36 0.17 0.465 0.785 ;
      RECT  0.36 0.785 1.02 0.895 ;
      RECT  0.36 0.895 0.465 1.525 ;
      RECT  0.56 1.205 1.225 1.32 ;
      RECT  1.105 1.32 1.225 1.415 ;
      RECT  1.105 1.415 1.745 1.505 ;
      RECT  1.625 1.505 1.745 1.615 ;
  END
END SEN_NR2B_V1DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1DG_3
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1DG_3
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.68 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.34 1.415 0.48 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  0.86 1.415 1.0 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.34 0.05 0.48 0.345 ;
      RECT  0.86 0.05 1.0 0.385 ;
      RECT  1.38 0.05 1.52 0.385 ;
      RECT  1.93 0.05 2.05 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.56 0.475 1.82 0.595 ;
      RECT  1.35 0.595 1.45 1.24 ;
      RECT  1.35 1.24 2.05 1.355 ;
      RECT  1.91 1.355 2.05 1.49 ;
    END
    ANTENNADIFFAREA 0.504 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.09 0.325 0.21 0.435 ;
      RECT  0.09 0.435 0.45 0.555 ;
      RECT  0.35 0.555 0.45 0.795 ;
      RECT  0.35 0.795 1.045 0.905 ;
      RECT  0.35 0.905 0.45 1.21 ;
      RECT  0.09 1.21 0.45 1.325 ;
      RECT  0.09 1.325 0.21 1.43 ;
      RECT  0.56 1.205 1.25 1.325 ;
      RECT  1.13 1.325 1.25 1.445 ;
      RECT  1.13 1.445 1.82 1.56 ;
  END
END SEN_NR2B_V1DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1DG_4
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1DG_4
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.215 0.185 1.75 ;
      RECT  0.0 1.75 2.8 1.85 ;
      RECT  0.79 1.23 0.91 1.75 ;
      RECT  1.315 1.23 1.435 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      RECT  1.05 0.05 1.17 0.38 ;
      RECT  1.575 0.05 1.695 0.38 ;
      RECT  2.095 0.05 2.215 0.38 ;
      RECT  0.065 0.05 0.185 0.385 ;
      RECT  0.53 0.05 0.65 0.385 ;
      RECT  2.615 0.05 2.735 0.57 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.765 0.47 2.5 0.59 ;
      RECT  1.75 0.59 1.85 1.235 ;
      RECT  1.75 1.235 2.5 1.35 ;
    END
    ANTENNADIFFAREA 0.624 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.49 0.43 0.79 ;
      RECT  0.34 0.79 1.335 0.91 ;
      RECT  0.34 0.91 0.43 1.58 ;
      RECT  0.545 1.02 1.66 1.14 ;
      RECT  0.545 1.14 0.635 1.195 ;
      RECT  1.54 1.14 1.66 1.44 ;
      RECT  1.54 1.44 2.735 1.555 ;
      RECT  2.615 1.555 2.735 1.61 ;
  END
END SEN_NR2B_V1DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1_1
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1_1
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.37 1.415 0.51 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.37 0.05 0.51 0.385 ;
      RECT  0.99 0.05 1.13 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.31 0.85 1.31 ;
      RECT  0.75 1.31 1.115 1.49 ;
    END
    ANTENNADIFFAREA 0.196 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.19 0.185 0.485 ;
      RECT  0.065 0.485 0.65 0.575 ;
      RECT  0.55 0.575 0.65 1.21 ;
      RECT  0.065 1.21 0.65 1.3 ;
      RECT  0.065 1.3 0.185 1.585 ;
  END
END SEN_NR2B_V1_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1_2
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1_2
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.51 0.255 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.835 1.415 0.975 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.095 0.05 1.235 0.385 ;
      RECT  1.615 0.05 1.745 0.385 ;
      RECT  0.055 0.05 0.185 0.39 ;
      RECT  0.585 0.05 0.705 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.795 0.475 1.65 0.595 ;
      RECT  1.55 0.595 1.65 1.11 ;
      RECT  1.35 1.11 1.65 1.29 ;
    END
    ANTENNADIFFAREA 0.288 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.35 0.155 0.455 0.755 ;
      RECT  0.35 0.755 1.015 0.865 ;
      RECT  0.35 0.865 0.455 1.515 ;
      RECT  0.585 1.205 1.225 1.32 ;
      RECT  1.105 1.32 1.225 1.415 ;
      RECT  0.585 1.32 0.705 1.435 ;
      RECT  1.105 1.415 1.745 1.505 ;
      RECT  1.625 1.505 1.745 1.63 ;
  END
END SEN_NR2B_V1_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR2B_V1_4
#      Description : "2-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR2B_V1_4
  CLASS CORE ;
  FOREIGN SEN_NR2B_V1_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.6 1.43 0.74 1.75 ;
      RECT  1.12 1.25 1.24 1.75 ;
      RECT  1.68 1.25 1.8 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  1.395 0.05 1.535 0.345 ;
      RECT  1.93 0.05 2.07 0.345 ;
      RECT  2.465 0.05 2.605 0.345 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  0.76 0.05 0.88 0.59 ;
      RECT  3.0 0.05 3.12 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.095 0.44 2.88 0.56 ;
      RECT  2.15 0.56 2.25 1.24 ;
      RECT  2.15 1.24 2.88 1.355 ;
    END
    ANTENNADIFFAREA 0.596 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.29 0.26 0.65 0.38 ;
      RECT  0.56 0.38 0.65 0.76 ;
      RECT  0.56 0.76 1.68 0.86 ;
      RECT  0.56 0.86 0.65 1.22 ;
      RECT  0.29 1.22 0.65 1.34 ;
      RECT  0.835 1.04 2.06 1.16 ;
      RECT  1.94 1.16 2.06 1.445 ;
      RECT  1.94 1.445 3.115 1.56 ;
      RECT  2.995 1.34 3.115 1.445 ;
  END
END SEN_NR2B_V1_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_0P5
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_0P5
  CLASS CORE ;
  FOREIGN SEN_NR3_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.705 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0303 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.065 0.05 0.195 0.39 ;
      RECT  0.615 0.05 0.745 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.2 0.46 0.48 ;
      RECT  0.34 0.48 1.05 0.59 ;
      RECT  0.95 0.2 1.05 0.48 ;
      RECT  0.95 0.59 1.05 1.51 ;
    END
    ANTENNADIFFAREA 0.143 ;
  END X
END SEN_NR3_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_1
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_1
  CLASS CORE ;
  FOREIGN SEN_NR3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.705 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.62 0.05 0.74 0.365 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.31 0.455 1.05 0.565 ;
      RECT  0.95 0.565 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.268 ;
  END X
END SEN_NR3_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_2
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_2
  CLASS CORE ;
  FOREIGN SEN_NR3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.45 0.455 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.585 0.05 0.715 0.35 ;
      RECT  1.195 0.05 1.325 0.35 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  1.815 0.05 1.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.305 0.44 1.7 0.56 ;
      RECT  1.35 0.56 1.45 1.11 ;
      RECT  1.35 1.11 1.66 1.29 ;
    END
    ANTENNADIFFAREA 0.366 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 1.015 1.23 1.24 ;
      RECT  0.07 1.24 1.23 1.36 ;
      RECT  0.07 1.36 0.185 1.46 ;
      RECT  1.815 1.34 1.935 1.45 ;
      RECT  0.8 1.45 1.935 1.56 ;
  END
END SEN_NR3_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_4
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_4
  CLASS CORE ;
  FOREIGN SEN_NR3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.45 0.71 ;
      RECT  2.95 0.71 3.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.45 0.455 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.845 1.45 0.975 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.585 0.05 0.715 0.35 ;
      RECT  1.105 0.05 1.235 0.35 ;
      RECT  1.625 0.05 1.755 0.35 ;
      RECT  2.255 0.05 2.385 0.35 ;
      RECT  2.885 0.05 3.015 0.35 ;
      RECT  3.405 0.05 3.535 0.39 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.3 3.26 0.44 ;
      RECT  0.305 0.44 3.26 0.56 ;
      RECT  2.55 0.56 2.65 1.11 ;
      RECT  2.55 1.11 3.27 1.29 ;
    END
    ANTENNADIFFAREA 0.732 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.15 0.98 2.27 1.24 ;
      RECT  0.07 1.24 2.27 1.36 ;
      RECT  0.07 1.36 0.19 1.46 ;
      RECT  3.41 1.34 3.53 1.45 ;
      RECT  1.32 1.45 3.53 1.56 ;
  END
END SEN_NR3_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_8
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_8
  CLASS CORE ;
  FOREIGN SEN_NR3_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.71 5.65 1.29 ;
      RECT  3.95 0.71 4.05 1.29 ;
      RECT  2.35 0.71 2.45 1.29 ;
      RECT  0.95 0.71 1.05 1.29 ;
      LAYER M2 ;
      RECT  0.91 1.15 5.69 1.25 ;
      LAYER V1 ;
      RECT  5.55 1.15 5.65 1.25 ;
      RECT  3.95 1.15 4.05 1.25 ;
      RECT  2.35 1.15 2.45 1.25 ;
      RECT  0.95 1.15 1.05 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.905 0.71 6.005 1.2 ;
      RECT  5.12 0.71 5.25 1.29 ;
      RECT  4.34 0.71 4.45 1.2 ;
      RECT  3.605 0.71 3.705 0.91 ;
      RECT  3.6 0.91 3.705 1.09 ;
      RECT  3.605 1.09 3.705 1.2 ;
      RECT  2.75 0.71 2.85 1.2 ;
      RECT  2.0 0.67 2.1 1.09 ;
      RECT  1.27 0.67 1.37 1.09 ;
      RECT  0.455 0.71 0.65 0.89 ;
      RECT  0.535 0.89 0.65 1.29 ;
      LAYER M2 ;
      RECT  0.51 0.95 6.045 1.05 ;
      LAYER V1 ;
      RECT  5.905 0.95 6.005 1.05 ;
      RECT  5.15 0.95 5.25 1.05 ;
      RECT  4.34 0.95 4.44 1.05 ;
      RECT  3.6 0.95 3.7 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  2.0 0.95 2.1 1.05 ;
      RECT  1.27 0.95 1.37 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.125 0.71 6.45 0.89 ;
      RECT  6.125 0.89 6.215 1.56 ;
      RECT  4.55 0.71 5.03 0.89 ;
      RECT  4.55 0.89 4.65 1.56 ;
      RECT  4.94 0.89 5.03 1.56 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  2.95 0.89 3.05 1.56 ;
      RECT  3.38 0.89 3.47 1.56 ;
      RECT  1.46 0.71 1.91 0.89 ;
      RECT  1.46 0.89 1.55 1.56 ;
      RECT  1.82 0.89 1.91 1.56 ;
      RECT  0.15 0.71 0.365 1.09 ;
      RECT  0.275 1.09 0.365 1.56 ;
      RECT  0.275 1.56 1.55 1.65 ;
      RECT  1.82 1.56 3.05 1.65 ;
      RECT  3.38 1.56 4.65 1.65 ;
      RECT  4.94 1.56 6.215 1.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.64 1.18 1.73 1.75 ;
      RECT  3.185 1.15 3.29 1.75 ;
      RECT  4.76 1.18 4.85 1.75 ;
      RECT  6.33 1.1 6.45 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  1.625 0.05 1.745 0.36 ;
      RECT  2.145 0.05 2.265 0.36 ;
      RECT  2.665 0.05 2.785 0.36 ;
      RECT  3.185 0.05 3.305 0.36 ;
      RECT  3.705 0.05 3.825 0.36 ;
      RECT  4.225 0.05 4.345 0.36 ;
      RECT  4.745 0.05 4.865 0.36 ;
      RECT  5.28 0.05 5.4 0.36 ;
      RECT  0.555 0.05 0.675 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.45 5.45 0.58 ;
      RECT  2.55 0.58 4.25 0.62 ;
      RECT  0.75 0.58 0.85 1.38 ;
      RECT  5.35 0.58 5.45 1.38 ;
      RECT  2.55 0.62 2.65 1.38 ;
      RECT  4.15 0.62 4.25 1.38 ;
      RECT  0.75 1.38 1.025 1.47 ;
      RECT  2.345 1.38 2.65 1.47 ;
      RECT  3.91 1.38 4.25 1.47 ;
      RECT  5.35 1.38 5.67 1.47 ;
    END
    ANTENNADIFFAREA 1.29 ;
  END X
END SEN_NR3_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_G_8
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_G_8
  CLASS CORE ;
  FOREIGN SEN_NR3_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.71 5.65 1.29 ;
      RECT  3.95 0.71 4.05 1.29 ;
      RECT  2.35 0.71 2.45 1.29 ;
      RECT  0.95 0.71 1.05 1.29 ;
      LAYER M2 ;
      RECT  0.91 1.15 5.69 1.25 ;
      LAYER V1 ;
      RECT  5.55 1.15 5.65 1.25 ;
      RECT  3.95 1.15 4.05 1.25 ;
      RECT  2.35 1.15 2.45 1.25 ;
      RECT  0.95 1.15 1.05 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.905 0.71 6.005 1.2 ;
      RECT  5.12 0.71 5.25 1.29 ;
      RECT  4.34 0.71 4.45 1.2 ;
      RECT  3.605 0.71 3.705 0.91 ;
      RECT  3.6 0.91 3.705 1.09 ;
      RECT  3.605 1.09 3.705 1.2 ;
      RECT  2.75 0.71 2.85 1.2 ;
      RECT  2.0 0.67 2.1 1.09 ;
      RECT  1.27 0.67 1.37 1.09 ;
      RECT  0.455 0.71 0.65 0.89 ;
      RECT  0.535 0.89 0.65 1.29 ;
      LAYER M2 ;
      RECT  0.51 0.95 6.045 1.05 ;
      LAYER V1 ;
      RECT  5.905 0.95 6.005 1.05 ;
      RECT  5.15 0.95 5.25 1.05 ;
      RECT  4.34 0.95 4.44 1.05 ;
      RECT  3.6 0.95 3.7 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  2.0 0.95 2.1 1.05 ;
      RECT  1.27 0.95 1.37 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.125 0.71 6.45 0.89 ;
      RECT  6.125 0.89 6.215 1.56 ;
      RECT  4.55 0.71 5.03 0.89 ;
      RECT  4.55 0.89 4.65 1.56 ;
      RECT  4.94 0.89 5.03 1.56 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  2.95 0.89 3.05 1.56 ;
      RECT  3.38 0.89 3.47 1.56 ;
      RECT  1.46 0.71 1.91 0.89 ;
      RECT  1.46 0.89 1.55 1.56 ;
      RECT  1.82 0.89 1.91 1.56 ;
      RECT  0.15 0.71 0.365 1.09 ;
      RECT  0.275 1.09 0.365 1.56 ;
      RECT  0.275 1.56 1.55 1.65 ;
      RECT  1.82 1.56 3.05 1.65 ;
      RECT  3.38 1.56 4.65 1.65 ;
      RECT  4.94 1.56 6.215 1.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.64 1.155 1.73 1.75 ;
      RECT  3.185 1.185 3.29 1.75 ;
      RECT  4.76 1.185 4.85 1.75 ;
      RECT  6.33 1.07 6.45 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.585 0.05 0.705 0.36 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  1.625 0.05 1.745 0.36 ;
      RECT  2.145 0.05 2.265 0.36 ;
      RECT  2.665 0.05 2.785 0.36 ;
      RECT  3.185 0.05 3.305 0.36 ;
      RECT  3.705 0.05 3.825 0.36 ;
      RECT  4.225 0.05 4.345 0.36 ;
      RECT  4.745 0.05 4.865 0.36 ;
      RECT  5.265 0.05 5.385 0.36 ;
      RECT  5.785 0.05 5.905 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.33 0.05 6.45 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.45 6.215 0.57 ;
      RECT  0.75 0.57 5.45 0.58 ;
      RECT  2.55 0.58 4.25 0.62 ;
      RECT  0.75 0.58 0.85 1.38 ;
      RECT  5.35 0.58 5.45 1.38 ;
      RECT  2.55 0.62 2.65 1.38 ;
      RECT  4.15 0.62 4.25 1.38 ;
      RECT  0.75 1.38 1.03 1.47 ;
      RECT  2.35 1.38 2.65 1.47 ;
      RECT  3.9 1.38 4.25 1.47 ;
      RECT  5.35 1.38 5.7 1.47 ;
    END
    ANTENNADIFFAREA 1.632 ;
  END X
END SEN_NR3_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_0P65
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_0P65
  CLASS CORE ;
  FOREIGN SEN_NR3_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.7 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.905 ;
      RECT  0.95 0.905 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.9 1.21 1.02 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.63 0.05 0.76 0.365 ;
      RECT  0.06 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.18 0.45 0.455 ;
      RECT  0.35 0.455 1.05 0.545 ;
      RECT  0.95 0.185 1.05 0.455 ;
      RECT  0.35 0.545 0.45 1.31 ;
      RECT  0.065 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.147 ;
  END X
END SEN_NR3_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_0P8
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_0P8
  CLASS CORE ;
  FOREIGN SEN_NR3_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.685 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.9 1.21 1.02 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.63 0.05 0.77 0.365 ;
      RECT  0.06 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.18 0.45 0.455 ;
      RECT  0.35 0.455 1.05 0.545 ;
      RECT  0.95 0.185 1.05 0.455 ;
      RECT  0.35 0.545 0.45 1.31 ;
      RECT  0.065 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.18 ;
  END X
END SEN_NR3_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_0P5
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_0P5
  CLASS CORE ;
  FOREIGN SEN_NR3_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.67 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0399 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0399 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.91 1.21 1.03 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.63 0.05 0.77 0.365 ;
      RECT  0.06 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.17 0.46 0.455 ;
      RECT  0.35 0.455 1.05 0.545 ;
      RECT  0.95 0.18 1.05 0.455 ;
      RECT  0.35 0.545 0.45 1.31 ;
      RECT  0.065 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.133 ;
  END X
END SEN_NR3_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_0P65
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_0P65
  CLASS CORE ;
  FOREIGN SEN_NR3_T_0P65 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0366 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.635 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.67 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.91 1.21 1.03 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.63 0.05 0.77 0.365 ;
      RECT  0.06 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.155 0.46 0.455 ;
      RECT  0.35 0.455 1.05 0.545 ;
      RECT  0.95 0.195 1.05 0.455 ;
      RECT  0.35 0.545 0.45 1.31 ;
      RECT  0.065 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.147 ;
  END X
END SEN_NR3_T_0P65
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_0P8
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_0P8
  CLASS CORE ;
  FOREIGN SEN_NR3_T_0P8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.165 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.045 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.665 0.66 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0588 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.71 ;
      RECT  0.95 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0588 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.915 1.39 1.045 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.11 0.05 0.25 0.39 ;
      RECT  0.66 0.05 0.78 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.175 0.505 0.485 ;
      RECT  0.35 0.485 1.06 0.575 ;
      RECT  0.94 0.175 1.06 0.485 ;
      RECT  0.35 0.575 0.45 1.31 ;
      RECT  0.15 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.18 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.66 1.21 1.3 1.3 ;
      RECT  0.66 1.3 0.78 1.515 ;
      RECT  1.18 1.3 1.3 1.545 ;
  END
END SEN_NR3_T_0P8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_1
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_1
  CLASS CORE ;
  FOREIGN SEN_NR3_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0561 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0735 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0735 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  0.575 1.44 0.705 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.9 0.05 1.1 0.365 ;
      RECT  1.61 0.05 1.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.215 0.66 0.455 ;
      RECT  0.55 0.455 1.45 0.545 ;
      RECT  1.34 0.25 1.45 0.455 ;
      RECT  1.35 0.545 1.45 1.25 ;
      RECT  1.35 1.25 1.735 1.34 ;
      RECT  1.615 1.34 1.735 1.48 ;
    END
    ANTENNADIFFAREA 0.227 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.275 1.24 1.26 1.35 ;
      RECT  0.81 1.445 1.525 1.56 ;
  END
END SEN_NR3_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_12
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_12
  CLASS CORE ;
  FOREIGN SEN_NR3_T_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.35 0.71 10.65 0.89 ;
      RECT  10.55 0.89 10.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6624 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.825 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8424 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.66 2.85 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8424 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.4 0.445 1.75 ;
      RECT  0.0 1.75 10.8 1.85 ;
      RECT  0.865 1.385 0.985 1.75 ;
      RECT  1.445 1.39 1.565 1.75 ;
      RECT  1.965 1.385 2.085 1.75 ;
      RECT  2.485 1.385 2.605 1.75 ;
      RECT  3.005 1.39 3.125 1.75 ;
      RECT  3.525 1.39 3.645 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      RECT  4.81 0.05 4.98 0.22 ;
      RECT  5.35 0.05 5.52 0.22 ;
      RECT  5.89 0.05 6.06 0.22 ;
      RECT  6.43 0.05 6.6 0.22 ;
      RECT  2.185 0.05 2.325 0.24 ;
      RECT  2.725 0.05 2.865 0.265 ;
      RECT  1.115 0.05 1.235 0.315 ;
      RECT  1.655 0.05 1.775 0.315 ;
      RECT  0.56 0.05 0.73 0.355 ;
      RECT  8.025 0.05 8.145 0.355 ;
      RECT  8.545 0.05 8.665 0.355 ;
      RECT  9.065 0.05 9.185 0.355 ;
      RECT  9.585 0.05 9.705 0.355 ;
      RECT  10.105 0.05 10.225 0.355 ;
      RECT  7.0 0.05 7.11 0.37 ;
      RECT  7.505 0.05 7.625 0.37 ;
      RECT  10.62 0.05 10.745 0.39 ;
      RECT  3.265 0.05 3.385 0.41 ;
      RECT  3.785 0.05 3.905 0.41 ;
      RECT  4.305 0.05 4.425 0.41 ;
      RECT  0.065 0.05 0.185 0.48 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.225 7.885 0.445 ;
      RECT  7.75 0.445 10.535 0.51 ;
      RECT  4.515 0.31 6.91 0.49 ;
      RECT  4.515 0.49 4.685 0.5 ;
      RECT  6.74 0.49 6.91 0.51 ;
      RECT  3.54 0.31 3.65 0.5 ;
      RECT  3.54 0.5 4.685 0.51 ;
      RECT  4.06 0.335 4.15 0.5 ;
      RECT  1.94 0.31 2.05 0.355 ;
      RECT  1.94 0.355 3.125 0.405 ;
      RECT  2.95 0.31 3.125 0.355 ;
      RECT  0.82 0.405 3.125 0.445 ;
      RECT  0.325 0.31 0.45 0.445 ;
      RECT  0.325 0.445 3.125 0.51 ;
      RECT  0.325 0.51 4.685 0.535 ;
      RECT  6.74 0.51 10.535 0.535 ;
      RECT  7.245 0.22 7.365 0.51 ;
      RECT  2.95 0.535 4.685 0.69 ;
      RECT  6.74 0.535 9.25 0.69 ;
      RECT  8.95 0.69 9.25 1.11 ;
      RECT  8.02 1.11 10.45 1.2 ;
      RECT  8.02 1.2 10.745 1.29 ;
      RECT  10.625 1.29 10.745 1.62 ;
    END
    ANTENNADIFFAREA 1.885 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.72 1.03 5.025 1.11 ;
      RECT  1.68 1.11 6.06 1.18 ;
      RECT  0.065 1.18 7.69 1.28 ;
      RECT  0.065 1.28 0.185 1.43 ;
      RECT  3.975 1.4 10.51 1.52 ;
      RECT  5.63 1.52 9.445 1.56 ;
      RECT  6.67 1.56 9.445 1.59 ;
      RECT  6.67 1.59 8.405 1.63 ;
  END
END SEN_NR3_T_12
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_2
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_2
  CLASS CORE ;
  FOREIGN SEN_NR3_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.685 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1122 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.685 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1482 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.685 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1482 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.685 1.44 1.805 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  2.21 1.21 2.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.62 0.05 0.79 0.32 ;
      RECT  1.27 0.05 1.445 0.32 ;
      RECT  1.98 0.05 2.1 0.585 ;
      RECT  0.125 0.05 0.245 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.335 0.41 1.855 0.53 ;
      RECT  0.55 0.53 0.65 1.11 ;
      RECT  0.35 1.11 0.65 1.29 ;
    END
    ANTENNADIFFAREA 0.324 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.81 1.225 2.115 1.345 ;
      RECT  0.125 1.31 0.245 1.44 ;
      RECT  0.125 1.44 1.37 1.56 ;
  END
END SEN_NR3_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_3
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_3
  CLASS CORE ;
  FOREIGN SEN_NR3_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.925 ;
      RECT  0.35 0.925 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1656 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.96 ;
      RECT  1.35 0.96 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2181 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.65 3.05 0.75 ;
      RECT  2.95 0.75 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2181 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.4 1.44 2.54 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  2.92 1.44 3.055 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.84 0.05 0.98 0.36 ;
      RECT  1.38 0.05 1.52 0.36 ;
      RECT  2.13 0.05 2.27 0.36 ;
      RECT  2.66 0.05 2.8 0.36 ;
      RECT  0.28 0.05 0.42 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.295 2.53 0.45 ;
      RECT  0.535 0.45 3.05 0.56 ;
      RECT  2.93 0.295 3.05 0.45 ;
      RECT  0.75 0.56 0.85 1.22 ;
      RECT  0.07 1.22 0.85 1.345 ;
      RECT  0.07 1.345 0.19 1.475 ;
    END
    ANTENNADIFFAREA 0.523 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.04 1.24 3.31 1.35 ;
      RECT  3.19 1.35 3.31 1.48 ;
      RECT  0.28 1.44 2.08 1.56 ;
  END
END SEN_NR3_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_4
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_4
  CLASS CORE ;
  FOREIGN SEN_NR3_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.685 0.65 0.9 ;
      RECT  0.15 0.9 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2241 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.655 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2961 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.635 3.65 0.735 ;
      RECT  3.55 0.735 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2961 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.765 1.44 2.905 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  3.285 1.44 3.42 1.75 ;
      RECT  3.815 1.21 3.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.565 0.05 0.735 0.315 ;
      RECT  1.085 0.05 1.255 0.315 ;
      RECT  1.605 0.05 1.775 0.315 ;
      RECT  2.125 0.05 2.295 0.315 ;
      RECT  2.775 0.05 2.895 0.345 ;
      RECT  3.295 0.05 3.415 0.345 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  3.805 0.05 3.94 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.515 0.255 2.65 0.405 ;
      RECT  0.28 0.405 2.65 0.435 ;
      RECT  0.28 0.435 3.675 0.525 ;
      RECT  3.035 0.255 3.16 0.435 ;
      RECT  3.55 0.255 3.675 0.435 ;
      RECT  0.95 0.525 1.05 1.11 ;
      RECT  0.34 1.11 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.658 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.32 1.215 3.725 1.345 ;
      RECT  0.065 1.335 0.19 1.435 ;
      RECT  0.065 1.435 2.33 1.46 ;
      RECT  0.07 1.46 2.33 1.565 ;
  END
END SEN_NR3_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_5
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_5
  CLASS CORE ;
  FOREIGN SEN_NR3_T_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 4.85 0.71 ;
      RECT  3.95 0.71 4.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2796 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.7 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3516 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.68 ;
      RECT  0.15 0.68 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3516 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.35 1.44 0.47 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  0.87 1.44 0.99 1.75 ;
      RECT  1.39 1.44 1.51 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.59 0.05 0.71 0.36 ;
      RECT  1.12 0.05 1.24 0.36 ;
      RECT  1.735 0.05 1.855 0.36 ;
      RECT  2.43 0.05 2.55 0.36 ;
      RECT  2.95 0.05 3.07 0.36 ;
      RECT  3.47 0.05 3.59 0.36 ;
      RECT  3.99 0.05 4.11 0.36 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  4.53 0.05 4.65 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.25 0.45 0.45 ;
      RECT  0.34 0.45 4.42 0.54 ;
      RECT  0.85 0.255 0.97 0.45 ;
      RECT  1.405 0.255 1.51 0.45 ;
      RECT  2.15 0.25 2.275 0.45 ;
      RECT  2.69 0.25 2.795 0.45 ;
      RECT  3.21 0.25 3.33 0.45 ;
      RECT  3.745 0.54 4.42 0.56 ;
      RECT  3.745 0.56 3.855 1.105 ;
      RECT  3.745 1.105 4.89 1.29 ;
    END
    ANTENNADIFFAREA 0.83 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.18 3.385 1.33 ;
      RECT  0.07 1.33 0.19 1.42 ;
      RECT  1.855 1.425 4.685 1.575 ;
  END
END SEN_NR3_T_5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_6
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_6
  CLASS CORE ;
  FOREIGN SEN_NR3_T_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.23 0.71 5.45 0.895 ;
      RECT  5.35 0.895 5.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3312 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.635 3.65 0.735 ;
      RECT  3.55 0.735 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4392 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.61 0.63 1.65 0.74 ;
      RECT  1.55 0.74 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4392 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.61 1.44 0.73 1.75 ;
      RECT  1.13 1.44 1.25 1.75 ;
      RECT  1.65 1.44 1.77 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.59 0.05 0.71 0.36 ;
      RECT  1.11 0.05 1.23 0.36 ;
      RECT  1.65 0.05 1.77 0.36 ;
      RECT  2.17 0.05 2.29 0.36 ;
      RECT  2.69 0.05 2.81 0.36 ;
      RECT  3.21 0.05 3.33 0.36 ;
      RECT  3.76 0.05 3.88 0.36 ;
      RECT  4.22 0.05 4.34 0.36 ;
      RECT  4.77 0.05 4.89 0.36 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  5.32 0.05 5.44 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.33 0.255 0.45 0.45 ;
      RECT  0.33 0.45 5.2 0.54 ;
      RECT  0.85 0.26 0.97 0.45 ;
      RECT  1.405 0.26 1.51 0.45 ;
      RECT  1.91 0.255 2.05 0.45 ;
      RECT  2.41 0.255 2.535 0.45 ;
      RECT  2.95 0.255 3.055 0.45 ;
      RECT  3.47 0.255 3.59 0.45 ;
      RECT  3.95 0.54 5.2 0.56 ;
      RECT  3.95 0.56 4.08 1.105 ;
      RECT  3.95 1.105 5.25 1.29 ;
    END
    ANTENNADIFFAREA 0.942 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 1.18 3.65 1.33 ;
      RECT  2.145 1.425 5.415 1.575 ;
      RECT  5.29 1.575 5.415 1.645 ;
  END
END SEN_NR3_T_6
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_T_8
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_T_8
  CLASS CORE ;
  FOREIGN SEN_NR3_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.325 0.71 6.85 0.89 ;
      RECT  6.75 0.89 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.905 0.635 4.45 0.735 ;
      RECT  4.35 0.735 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5562 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.635 2.075 0.735 ;
      RECT  0.75 0.735 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5562 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  1.625 1.44 1.745 1.75 ;
      RECT  2.145 1.44 2.265 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  1.08 0.05 1.265 0.305 ;
      RECT  1.6 0.05 1.77 0.305 ;
      RECT  2.12 0.05 2.29 0.305 ;
      RECT  2.64 0.05 2.81 0.305 ;
      RECT  3.16 0.05 3.33 0.305 ;
      RECT  3.68 0.05 3.865 0.305 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.785 0.05 4.905 0.345 ;
      RECT  0.585 0.05 0.705 0.36 ;
      RECT  5.24 0.05 5.385 0.36 ;
      RECT  5.785 0.05 5.905 0.36 ;
      RECT  6.305 0.05 6.425 0.36 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  6.815 0.05 6.94 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.31 3.05 0.395 ;
      RECT  0.82 0.395 4.65 0.45 ;
      RECT  4.5 0.285 4.65 0.395 ;
      RECT  0.325 0.24 0.45 0.45 ;
      RECT  0.325 0.45 6.735 0.545 ;
      RECT  4.525 0.545 6.735 0.58 ;
      RECT  4.945 0.58 5.115 1.105 ;
      RECT  4.945 1.105 6.65 1.19 ;
      RECT  4.945 1.19 6.755 1.29 ;
    END
    ANTENNADIFFAREA 1.284 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.345 1.15 3.585 1.19 ;
      RECT  0.275 1.19 4.66 1.32 ;
      RECT  2.64 1.425 6.945 1.555 ;
      RECT  4.225 1.555 5.385 1.595 ;
      RECT  6.825 1.555 6.945 1.625 ;
  END
END SEN_NR3_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_G_1
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_G_1
  CLASS CORE ;
  FOREIGN SEN_NR3_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.91 1.21 1.03 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.63 0.05 0.77 0.365 ;
      RECT  0.06 0.05 0.195 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.19 0.46 0.455 ;
      RECT  0.35 0.455 1.05 0.545 ;
      RECT  0.95 0.3 1.05 0.455 ;
      RECT  0.35 0.545 0.45 1.31 ;
      RECT  0.065 1.31 0.45 1.49 ;
    END
    ANTENNADIFFAREA 0.279 ;
  END X
END SEN_NR3_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_G_2
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_G_2
  CLASS CORE ;
  FOREIGN SEN_NR3_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.93 ;
      RECT  0.15 0.93 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.925 ;
      RECT  0.75 0.925 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.05 0.925 ;
      RECT  1.95 0.925 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.455 1.24 1.575 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  2.01 1.21 2.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.635 0.05 0.775 0.36 ;
      RECT  1.295 0.05 1.435 0.36 ;
      RECT  0.11 0.05 0.23 0.59 ;
      RECT  2.01 0.05 2.13 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.335 0.455 1.895 0.545 ;
      RECT  0.55 0.545 0.65 1.11 ;
      RECT  0.35 1.11 0.65 1.29 ;
    END
    ANTENNADIFFAREA 0.438 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.945 1.04 1.845 1.15 ;
      RECT  0.945 1.15 1.065 1.26 ;
      RECT  1.73 1.15 1.845 1.26 ;
      RECT  0.125 1.32 0.245 1.44 ;
      RECT  0.125 1.44 1.365 1.56 ;
  END
END SEN_NR3_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_G_3
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_G_3
  CLASS CORE ;
  FOREIGN SEN_NR3_G_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.925 ;
      RECT  0.35 0.925 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.46 0.925 ;
      RECT  1.15 0.925 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.935 0.71 2.25 0.925 ;
      RECT  2.15 0.925 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.875 1.44 2.015 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  2.405 1.21 2.525 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.575 0.05 0.715 0.36 ;
      RECT  1.095 0.05 1.235 0.36 ;
      RECT  1.615 0.05 1.755 0.36 ;
      RECT  2.135 0.05 2.275 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.405 0.3 2.525 0.455 ;
      RECT  0.275 0.455 2.525 0.545 ;
      RECT  0.75 0.545 0.85 1.24 ;
      RECT  0.065 1.24 0.85 1.345 ;
      RECT  0.065 1.345 0.185 1.46 ;
    END
    ANTENNADIFFAREA 0.677 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.055 1.245 2.315 1.345 ;
      RECT  0.275 1.44 1.54 1.56 ;
  END
END SEN_NR3_G_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3_G_4
#      Description : "3-Input NOR"
#      Equation    : X=!(A1|A2|A3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3_G_4
  CLASS CORE ;
  FOREIGN SEN_NR3_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.685 0.9 ;
      RECT  0.15 0.9 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.885 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.375 1.44 2.505 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  2.885 1.44 3.025 1.75 ;
      RECT  3.415 1.21 3.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.565 0.05 0.705 0.36 ;
      RECT  1.085 0.05 1.225 0.36 ;
      RECT  1.605 0.05 1.745 0.36 ;
      RECT  2.245 0.05 2.385 0.36 ;
      RECT  2.885 0.05 3.025 0.36 ;
      RECT  0.055 0.05 0.185 0.39 ;
      RECT  3.415 0.05 3.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.26 0.45 3.325 0.56 ;
      RECT  0.95 0.56 1.05 1.11 ;
      RECT  0.35 1.11 1.05 1.2 ;
      RECT  0.26 1.2 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.816 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.3 1.23 3.325 1.34 ;
      RECT  0.055 1.43 2.28 1.55 ;
      RECT  0.055 1.55 0.175 1.625 ;
  END
END SEN_NR3_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3B_1
#      Description : "3-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3B_1
  CLASS CORE ;
  FOREIGN SEN_NR3B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.195 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0516 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.51 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0606 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.465 0.47 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.92 0.05 1.04 0.36 ;
      RECT  0.32 0.05 0.455 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.57 0.265 0.83 0.385 ;
      RECT  0.74 0.385 0.83 0.45 ;
      RECT  0.74 0.45 1.295 0.54 ;
      RECT  1.15 0.54 1.295 0.69 ;
      RECT  1.185 0.69 1.295 1.11 ;
      RECT  1.15 1.11 1.295 1.495 ;
    END
    ANTENNADIFFAREA 0.25 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.945 0.775 1.085 0.95 ;
      RECT  0.945 0.95 1.035 1.485 ;
      RECT  0.055 0.38 0.175 0.515 ;
      RECT  0.055 0.515 0.43 0.605 ;
      RECT  0.34 0.605 0.43 1.285 ;
      RECT  0.055 1.285 0.65 1.375 ;
      RECT  0.56 1.375 0.65 1.485 ;
      RECT  0.055 1.375 0.175 1.62 ;
      RECT  0.56 1.485 1.035 1.575 ;
  END
END SEN_NR3B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3B_2
#      Description : "3-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3B_2
  CLASS CORE ;
  FOREIGN SEN_NR3B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.65 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1032 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1212 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.05 1.41 0.18 1.75 ;
      RECT  0.0 1.75 2.8 1.85 ;
      RECT  0.57 1.42 0.7 1.75 ;
      RECT  2.07 1.42 2.2 1.75 ;
      RECT  2.6 1.215 2.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      RECT  1.875 0.05 2.005 0.385 ;
      RECT  0.05 0.05 0.18 0.39 ;
      RECT  0.625 0.05 0.755 0.39 ;
      RECT  1.27 0.05 1.4 0.39 ;
      RECT  2.53 0.05 2.65 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.29 0.5 1.76 0.59 ;
      RECT  1.35 0.59 1.45 1.11 ;
      RECT  1.35 1.11 1.855 1.29 ;
    END
    ANTENNADIFFAREA 0.366 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.195 0.36 2.315 0.5 ;
      RECT  1.945 0.5 2.315 0.59 ;
      RECT  1.945 0.59 2.05 0.75 ;
      RECT  1.55 0.75 2.05 0.855 ;
      RECT  1.945 0.855 2.05 1.21 ;
      RECT  1.945 1.21 2.485 1.33 ;
      RECT  0.26 1.21 1.21 1.33 ;
      RECT  0.805 1.42 1.965 1.54 ;
      RECT  1.845 1.54 1.965 1.62 ;
      RECT  0.805 1.54 0.925 1.63 ;
  END
END SEN_NR3B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3B_3
#      Description : "3-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3B_3
  CLASS CORE ;
  FOREIGN SEN_NR3B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1548 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1818 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1818 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.185 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.57 1.445 0.7 1.75 ;
      RECT  2.895 1.415 3.025 1.75 ;
      RECT  3.415 1.41 3.54 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  2.895 0.05 3.025 0.365 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  0.57 0.05 0.7 0.39 ;
      RECT  1.09 0.05 1.22 0.39 ;
      RECT  1.61 0.05 1.74 0.39 ;
      RECT  2.13 0.05 2.27 0.39 ;
      RECT  3.415 0.05 3.545 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.395 0.37 2.515 0.48 ;
      RECT  0.26 0.48 2.515 0.59 ;
      RECT  1.75 0.59 1.85 1.11 ;
      RECT  1.75 1.11 2.515 1.29 ;
    END
    ANTENNADIFFAREA 0.61 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.615 0.455 3.305 0.575 ;
      RECT  2.615 0.575 2.705 0.745 ;
      RECT  1.94 0.745 2.705 0.855 ;
      RECT  2.615 0.855 2.705 1.19 ;
      RECT  2.615 1.19 3.33 1.315 ;
      RECT  0.29 1.235 1.53 1.355 ;
      RECT  1.04 1.445 2.31 1.565 ;
  END
END SEN_NR3B_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3B_4
#      Description : "3-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3B_4
  CLASS CORE ;
  FOREIGN SEN_NR3B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.9 0.695 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2064 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2424 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.575 1.435 0.715 1.75 ;
      RECT  1.095 1.43 1.23 1.75 ;
      RECT  3.83 1.415 3.96 1.75 ;
      RECT  4.38 1.215 4.5 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  1.655 0.05 1.785 0.36 ;
      RECT  2.79 0.05 2.92 0.36 ;
      RECT  3.88 0.05 4.015 0.365 ;
      RECT  0.57 0.05 0.72 0.37 ;
      RECT  2.2 0.05 2.33 0.37 ;
      RECT  1.1 0.05 1.23 0.375 ;
      RECT  4.42 0.05 4.55 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.34 0.05 3.46 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.3 0.47 3.23 0.59 ;
      RECT  2.55 0.59 2.65 1.11 ;
      RECT  2.55 1.11 3.25 1.29 ;
    END
    ANTENNADIFFAREA 0.736 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.57 0.46 4.33 0.58 ;
      RECT  3.57 0.58 3.695 0.75 ;
      RECT  2.805 0.75 3.695 0.85 ;
      RECT  3.57 0.85 3.695 1.205 ;
      RECT  3.57 1.205 4.27 1.32 ;
      RECT  1.265 1.025 1.86 1.135 ;
      RECT  1.77 1.135 1.86 1.205 ;
      RECT  1.77 1.205 2.455 1.325 ;
      RECT  2.325 1.325 2.455 1.445 ;
      RECT  2.325 1.445 3.54 1.565 ;
      RECT  0.3 1.225 1.67 1.34 ;
      RECT  1.55 1.34 1.67 1.44 ;
      RECT  1.55 1.44 2.215 1.56 ;
  END
END SEN_NR3B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR3B_DG_8
#      Description : "3-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR3B_DG_8
  CLASS CORE ;
  FOREIGN SEN_NR3B_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.51 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.905 0.71 6.005 1.2 ;
      RECT  5.12 0.71 5.25 1.29 ;
      RECT  4.34 0.71 4.45 1.2 ;
      RECT  3.6 0.71 3.715 1.2 ;
      RECT  2.75 0.71 2.85 1.2 ;
      RECT  2.0 0.67 2.1 1.09 ;
      RECT  1.27 0.67 1.37 1.09 ;
      RECT  0.455 0.71 0.65 0.89 ;
      RECT  0.535 0.89 0.65 1.29 ;
      LAYER M2 ;
      RECT  0.51 0.95 6.045 1.05 ;
      LAYER V1 ;
      RECT  5.905 0.95 6.005 1.05 ;
      RECT  5.15 0.95 5.25 1.05 ;
      RECT  4.34 0.95 4.44 1.05 ;
      RECT  3.6 0.95 3.7 1.05 ;
      RECT  2.75 0.95 2.85 1.05 ;
      RECT  2.0 0.95 2.1 1.05 ;
      RECT  1.27 0.95 1.37 1.05 ;
      RECT  0.55 0.95 0.65 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.125 0.71 6.45 0.89 ;
      RECT  6.125 0.89 6.215 1.56 ;
      RECT  4.55 0.71 5.03 0.89 ;
      RECT  4.55 0.89 4.65 1.56 ;
      RECT  4.94 0.89 5.03 1.56 ;
      RECT  2.95 0.71 3.47 0.89 ;
      RECT  2.95 0.89 3.05 1.56 ;
      RECT  3.38 0.89 3.47 1.56 ;
      RECT  1.46 0.71 1.91 0.89 ;
      RECT  1.46 0.89 1.55 1.56 ;
      RECT  1.82 0.89 1.91 1.56 ;
      RECT  0.15 0.71 0.365 1.09 ;
      RECT  0.275 1.09 0.365 1.56 ;
      RECT  0.275 1.56 1.55 1.65 ;
      RECT  1.82 1.56 3.05 1.65 ;
      RECT  3.38 1.56 4.65 1.65 ;
      RECT  4.94 1.56 6.215 1.65 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  1.64 1.19 1.73 1.75 ;
      RECT  3.185 1.185 3.29 1.75 ;
      RECT  4.76 1.2 4.85 1.75 ;
      RECT  6.305 1.16 6.425 1.75 ;
      RECT  6.825 1.41 6.945 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  0.585 0.05 0.705 0.36 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  1.625 0.05 1.745 0.36 ;
      RECT  2.145 0.05 2.265 0.36 ;
      RECT  2.665 0.05 2.785 0.36 ;
      RECT  3.185 0.05 3.305 0.36 ;
      RECT  3.705 0.05 3.825 0.36 ;
      RECT  4.225 0.05 4.345 0.36 ;
      RECT  4.745 0.05 4.865 0.36 ;
      RECT  5.265 0.05 5.385 0.36 ;
      RECT  5.785 0.05 5.905 0.36 ;
      RECT  6.825 0.05 6.945 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.305 0.05 6.425 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.275 0.45 6.215 0.57 ;
      RECT  0.75 0.57 5.45 0.58 ;
      RECT  2.55 0.58 4.25 0.62 ;
      RECT  0.75 0.58 0.85 1.38 ;
      RECT  5.35 0.58 5.45 1.38 ;
      RECT  2.55 0.62 2.65 1.38 ;
      RECT  4.15 0.62 4.25 1.38 ;
      RECT  0.75 1.38 1.015 1.47 ;
      RECT  2.355 1.38 2.65 1.47 ;
      RECT  3.915 1.38 4.25 1.47 ;
      RECT  5.35 1.38 5.695 1.47 ;
    END
    ANTENNADIFFAREA 1.632 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.54 0.24 6.735 0.36 ;
      RECT  6.54 0.36 6.64 1.24 ;
      RECT  6.54 1.24 6.735 1.36 ;
      RECT  0.95 0.71 1.05 1.29 ;
      RECT  2.35 0.71 2.45 1.29 ;
      RECT  3.95 0.71 4.05 1.29 ;
      RECT  5.55 0.71 5.65 1.29 ;
      LAYER M2 ;
      RECT  0.91 1.15 6.68 1.25 ;
      LAYER V1 ;
      RECT  0.95 1.15 1.05 1.25 ;
      RECT  2.35 1.15 2.45 1.25 ;
      RECT  3.95 1.15 4.05 1.25 ;
      RECT  5.55 1.15 5.65 1.25 ;
      RECT  6.54 1.15 6.64 1.25 ;
  END
END SEN_NR3B_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4_0P5
#      Description : "4-Input NOR"
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4_0P5
  CLASS CORE ;
  FOREIGN SEN_NR4_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.41 0.21 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.59 0.05 0.73 0.38 ;
      RECT  0.07 0.05 0.21 0.39 ;
      RECT  1.12 0.05 1.26 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.18 0.46 0.47 ;
      RECT  0.35 0.47 0.98 0.475 ;
      RECT  0.86 0.175 0.98 0.47 ;
      RECT  0.35 0.475 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.31 ;
      RECT  0.95 1.31 1.25 1.49 ;
    END
    ANTENNADIFFAREA 0.12 ;
  END X
END SEN_NR4_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4_1
#      Description : "4-Input NOR"
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4_1
  CLASS CORE ;
  FOREIGN SEN_NR4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.655 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.695 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.085 1.21 0.2 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.6 0.05 0.72 0.38 ;
      RECT  0.07 0.05 0.21 0.39 ;
      RECT  1.12 0.05 1.26 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.23 0.46 0.47 ;
      RECT  0.35 0.47 0.98 0.475 ;
      RECT  0.86 0.23 0.98 0.47 ;
      RECT  0.35 0.475 1.05 0.56 ;
      RECT  0.95 0.56 1.05 1.31 ;
      RECT  0.95 1.31 1.25 1.49 ;
    END
    ANTENNADIFFAREA 0.204 ;
  END X
END SEN_NR4_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4_2
#      Description : "4-Input NOR"
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4_2
  CLASS CORE ;
  FOREIGN SEN_NR4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.685 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.685 1.85 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.685 2.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.14 1.4 2.26 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.59 0.05 0.71 0.38 ;
      RECT  1.225 0.05 1.385 0.38 ;
      RECT  1.88 0.05 2.0 0.38 ;
      RECT  0.065 0.05 0.2 0.39 ;
      RECT  2.41 0.05 2.535 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.345 0.21 0.45 0.47 ;
      RECT  0.345 0.47 2.255 0.56 ;
      RECT  0.855 0.185 0.975 0.47 ;
      RECT  1.62 0.18 1.74 0.47 ;
      RECT  2.145 0.18 2.255 0.47 ;
      RECT  0.345 0.56 0.45 1.48 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.85 1.2 1.74 1.29 ;
      RECT  0.85 1.29 0.97 1.48 ;
      RECT  1.62 1.29 1.74 1.48 ;
      RECT  1.88 1.2 2.52 1.29 ;
      RECT  2.4 1.29 2.52 1.485 ;
      RECT  1.88 1.29 2.0 1.57 ;
      RECT  1.36 1.38 1.48 1.57 ;
      RECT  1.36 1.57 2.0 1.66 ;
      RECT  0.07 1.4 0.185 1.57 ;
      RECT  0.07 1.57 1.23 1.66 ;
      RECT  0.59 1.37 0.71 1.57 ;
      RECT  1.11 1.38 1.23 1.57 ;
  END
END SEN_NR4_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4_3
#      Description : "4-Input NOR"
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4_3
  CLASS CORE ;
  FOREIGN SEN_NR4_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.505 3.25 0.71 ;
      RECT  2.94 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1578 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.895 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1578 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.055 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1578 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.505 0.25 0.71 ;
      RECT  0.15 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1578 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.585 1.4 0.705 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.845 0.05 0.965 0.38 ;
      RECT  1.625 0.05 1.745 0.38 ;
      RECT  2.405 0.05 2.525 0.38 ;
      RECT  0.34 0.05 0.47 0.59 ;
      RECT  2.945 0.05 3.055 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.585 0.36 0.705 0.47 ;
      RECT  0.585 0.47 2.85 0.585 ;
      RECT  2.75 0.31 2.85 0.47 ;
      RECT  2.75 0.585 2.85 1.11 ;
      RECT  2.67 1.11 3.305 1.29 ;
    END
    ANTENNADIFFAREA 0.76 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 1.2 0.965 1.29 ;
      RECT  0.34 1.29 0.43 1.5 ;
      RECT  0.845 1.29 0.965 1.57 ;
      RECT  0.845 1.57 1.485 1.66 ;
      RECT  1.365 1.38 1.485 1.57 ;
      RECT  1.105 1.2 1.745 1.29 ;
      RECT  1.105 1.29 1.225 1.48 ;
      RECT  1.625 1.29 1.745 1.57 ;
      RECT  1.625 1.57 2.265 1.66 ;
      RECT  2.145 1.38 2.265 1.57 ;
      RECT  1.9 1.2 2.525 1.29 ;
      RECT  1.9 1.29 1.99 1.48 ;
      RECT  2.405 1.29 2.525 1.525 ;
      RECT  2.405 1.525 3.045 1.615 ;
      RECT  2.925 1.4 3.045 1.525 ;
  END
END SEN_NR4_3
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4_4
#      Description : "4-Input NOR"
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4_4
  CLASS CORE ;
  FOREIGN SEN_NR4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.685 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.21 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.685 1.91 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.21 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.685 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.21 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.685 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.21 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  3.63 1.41 3.75 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  4.15 1.41 4.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.585 0.05 0.705 0.355 ;
      RECT  1.105 0.05 1.225 0.355 ;
      RECT  1.625 0.05 1.745 0.355 ;
      RECT  2.24 0.05 2.36 0.355 ;
      RECT  2.85 0.05 2.97 0.355 ;
      RECT  3.37 0.05 3.49 0.355 ;
      RECT  3.89 0.05 4.01 0.355 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  4.4 0.05 4.54 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.225 0.45 0.445 ;
      RECT  0.34 0.445 4.27 0.56 ;
      RECT  0.845 0.225 0.965 0.445 ;
      RECT  1.35 0.225 1.485 0.445 ;
      RECT  1.885 0.225 2.05 0.445 ;
      RECT  2.55 0.23 2.71 0.445 ;
      RECT  3.11 0.23 3.25 0.445 ;
      RECT  3.63 0.23 3.75 0.445 ;
      RECT  4.15 0.23 4.27 0.445 ;
      RECT  0.75 0.56 0.85 1.11 ;
      RECT  0.34 1.11 0.965 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.045 1.025 2.71 1.12 ;
      RECT  2.045 1.12 2.15 1.14 ;
      RECT  2.59 1.12 2.71 1.24 ;
      RECT  1.325 1.14 2.15 1.26 ;
      RECT  2.59 1.24 3.255 1.36 ;
      RECT  3.37 1.2 4.53 1.32 ;
      RECT  3.37 1.32 3.49 1.465 ;
      RECT  4.41 1.32 4.53 1.475 ;
      RECT  2.295 1.21 2.475 1.33 ;
      RECT  2.385 1.33 2.475 1.465 ;
      RECT  2.385 1.465 3.49 1.6 ;
      RECT  0.065 1.345 0.19 1.465 ;
      RECT  0.065 1.465 2.265 1.61 ;
      RECT  2.145 1.415 2.265 1.465 ;
  END
END SEN_NR4_4
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4_6
#      Description : "4-Input NOR"
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4_6
  CLASS CORE ;
  FOREIGN SEN_NR4_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.065 0.71 5.85 0.89 ;
      RECT  5.75 0.89 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3156 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.5 0.67 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3156 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.67 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3156 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.48 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3156 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.305 1.48 0.475 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.825 1.48 0.995 1.75 ;
      RECT  1.345 1.48 1.515 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  0.565 0.05 0.735 0.32 ;
      RECT  1.215 0.05 1.385 0.32 ;
      RECT  1.865 0.05 2.035 0.32 ;
      RECT  2.385 0.05 2.555 0.32 ;
      RECT  2.905 0.05 3.075 0.32 ;
      RECT  4.615 0.05 4.785 0.32 ;
      RECT  5.245 0.05 5.415 0.32 ;
      RECT  3.425 0.05 3.595 0.325 ;
      RECT  3.945 0.05 4.115 0.325 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  5.805 0.05 5.925 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.345 0.31 0.45 0.43 ;
      RECT  0.345 0.43 5.65 0.56 ;
      RECT  1.63 0.255 1.75 0.43 ;
      RECT  2.15 0.255 2.27 0.43 ;
      RECT  2.67 0.255 2.79 0.43 ;
      RECT  3.19 0.255 3.31 0.43 ;
      RECT  3.71 0.26 3.855 0.43 ;
      RECT  4.23 0.255 4.35 0.43 ;
      RECT  5.53 0.3 5.65 0.43 ;
      RECT  4.75 0.56 4.88 1.11 ;
      RECT  4.35 1.11 5.65 1.295 ;
    END
    ANTENNADIFFAREA 1.018 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.865 1.235 4.145 1.365 ;
      RECT  0.07 1.25 1.755 1.38 ;
      RECT  0.07 1.38 0.19 1.47 ;
      RECT  1.625 1.38 1.755 1.475 ;
      RECT  1.625 1.475 2.815 1.605 ;
      RECT  5.79 1.37 5.91 1.475 ;
      RECT  3.15 1.475 5.91 1.605 ;
  END
END SEN_NR4_6
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4_8
#      Description : "4-Input NOR"
#      Equation    : X=!(A1|A2|A3|A4)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4_8
  CLASS CORE ;
  FOREIGN SEN_NR4_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.62 0.71 8.05 0.905 ;
      RECT  7.95 0.905 8.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.885 0.68 5.85 0.89 ;
      RECT  5.75 0.89 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.68 3.65 0.89 ;
      RECT  3.55 0.89 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4215 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.425 0.45 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.85 1.425 0.97 1.75 ;
      RECT  1.37 1.425 1.49 1.75 ;
      RECT  1.89 1.425 2.01 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  1.085 0.05 1.255 0.32 ;
      RECT  1.735 0.05 1.905 0.32 ;
      RECT  2.385 0.05 2.555 0.32 ;
      RECT  2.905 0.05 3.075 0.32 ;
      RECT  3.425 0.05 3.6 0.32 ;
      RECT  3.945 0.05 4.12 0.32 ;
      RECT  4.465 0.05 4.64 0.32 ;
      RECT  6.175 0.05 6.345 0.32 ;
      RECT  6.805 0.05 6.975 0.32 ;
      RECT  7.325 0.05 7.495 0.32 ;
      RECT  4.985 0.05 5.155 0.325 ;
      RECT  5.505 0.05 5.675 0.325 ;
      RECT  0.565 0.05 0.735 0.335 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.79 0.26 6.05 0.415 ;
      RECT  5.79 0.415 7.79 0.43 ;
      RECT  0.345 0.31 0.45 0.43 ;
      RECT  0.345 0.43 7.79 0.57 ;
      RECT  2.15 0.255 2.27 0.43 ;
      RECT  2.67 0.255 2.79 0.43 ;
      RECT  3.19 0.255 3.31 0.43 ;
      RECT  3.71 0.26 3.85 0.43 ;
      RECT  4.23 0.26 4.35 0.43 ;
      RECT  4.75 0.26 4.87 0.43 ;
      RECT  5.27 0.26 5.415 0.43 ;
      RECT  6.35 0.57 7.79 0.58 ;
      RECT  6.35 0.58 6.52 1.11 ;
      RECT  5.95 1.11 7.85 1.29 ;
    END
    ANTENNADIFFAREA 1.424 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 1.185 2.285 1.325 ;
      RECT  0.07 1.325 0.19 1.45 ;
      RECT  2.145 1.325 2.285 1.475 ;
      RECT  2.145 1.475 3.87 1.615 ;
      RECT  2.38 1.225 5.675 1.365 ;
      RECT  4.205 1.475 8.04 1.615 ;
  END
END SEN_NR4_8
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4B_1
#      Description : "4-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4B_1
  CLASS CORE ;
  FOREIGN SEN_NR4B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.185 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0219 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.705 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.535 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0525 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.455 0.445 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.855 0.05 0.975 0.22 ;
      RECT  1.395 0.05 1.515 0.22 ;
      RECT  0.325 0.05 0.445 0.42 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.535 0.31 1.505 0.43 ;
      RECT  1.35 0.43 1.505 0.57 ;
      RECT  1.4 0.57 1.505 1.11 ;
      RECT  1.35 1.11 1.505 1.49 ;
    END
    ANTENNADIFFAREA 0.204 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.185 0.185 0.525 ;
      RECT  0.065 0.525 1.25 0.615 ;
      RECT  1.15 0.615 1.25 0.665 ;
      RECT  1.15 0.665 1.305 0.835 ;
      RECT  1.15 0.835 1.25 1.455 ;
      RECT  0.065 1.275 0.645 1.365 ;
      RECT  0.555 1.365 0.645 1.455 ;
      RECT  0.065 1.365 0.185 1.62 ;
      RECT  0.555 1.455 1.25 1.545 ;
  END
END SEN_NR4B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4B_2
#      Description : "4-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4B_2
  CLASS CORE ;
  FOREIGN SEN_NR4B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.042 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.685 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.685 2.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.685 2.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.105 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  2.56 1.38 2.68 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  1.075 0.05 1.195 0.38 ;
      RECT  1.685 0.05 1.815 0.38 ;
      RECT  2.3 0.05 2.42 0.38 ;
      RECT  0.06 0.05 0.195 0.39 ;
      RECT  2.81 0.05 2.94 0.39 ;
      RECT  0.555 0.05 0.675 0.415 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.815 0.215 0.935 0.47 ;
      RECT  0.815 0.47 2.675 0.56 ;
      RECT  1.33 0.185 1.455 0.47 ;
      RECT  2.04 0.185 2.165 0.47 ;
      RECT  2.55 0.185 2.675 0.47 ;
      RECT  0.95 0.56 1.05 1.11 ;
      RECT  0.73 1.11 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.28 0.445 0.685 ;
      RECT  0.34 0.685 0.84 0.795 ;
      RECT  0.34 0.795 0.445 1.42 ;
      RECT  1.14 1.045 1.74 1.165 ;
      RECT  1.14 1.165 1.23 1.45 ;
      RECT  0.53 1.45 1.23 1.57 ;
      RECT  2.3 1.2 2.94 1.29 ;
      RECT  2.3 1.29 2.42 1.465 ;
      RECT  2.82 1.29 2.94 1.62 ;
      RECT  1.725 1.465 2.42 1.585 ;
      RECT  1.335 1.255 2.21 1.375 ;
      RECT  1.335 1.375 1.455 1.515 ;
  END
END SEN_NR4B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_NR4B_4
#      Description : "4-Input NOR (A inverted input)"
#      Equation    : X=!(!A|B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_NR4B_4
  CLASS CORE ;
  FOREIGN SEN_NR4B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0792 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.03 0.635 2.65 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.83 0.635 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2106 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.585 1.395 0.695 1.75 ;
      RECT  3.63 1.41 3.75 1.75 ;
      RECT  4.15 1.41 4.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  1.29 0.05 1.41 0.345 ;
      RECT  1.81 0.05 1.93 0.345 ;
      RECT  2.33 0.05 2.45 0.345 ;
      RECT  2.85 0.05 2.97 0.345 ;
      RECT  3.37 0.05 3.49 0.345 ;
      RECT  3.89 0.05 4.01 0.345 ;
      RECT  0.77 0.05 0.89 0.37 ;
      RECT  0.19 0.05 0.33 0.39 ;
      RECT  4.41 0.05 4.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.03 0.18 1.15 0.435 ;
      RECT  1.03 0.435 4.27 0.525 ;
      RECT  1.55 0.175 1.67 0.435 ;
      RECT  2.07 0.175 2.19 0.435 ;
      RECT  2.55 0.185 2.71 0.435 ;
      RECT  3.11 0.185 3.25 0.435 ;
      RECT  3.63 0.18 3.75 0.435 ;
      RECT  4.15 0.18 4.27 0.435 ;
      RECT  1.75 0.525 1.85 1.11 ;
      RECT  1.005 1.11 1.85 1.29 ;
    END
    ANTENNADIFFAREA 0.684 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.51 0.175 0.63 0.47 ;
      RECT  0.51 0.47 0.83 0.56 ;
      RECT  0.74 0.56 0.83 0.755 ;
      RECT  0.74 0.755 1.45 0.865 ;
      RECT  0.74 0.865 0.83 1.005 ;
      RECT  0.325 1.005 0.83 1.095 ;
      RECT  0.325 1.095 0.445 1.555 ;
      RECT  3.37 1.2 4.53 1.32 ;
      RECT  3.37 1.32 3.49 1.43 ;
      RECT  4.41 1.32 4.53 1.45 ;
      RECT  2.8 1.43 3.49 1.55 ;
      RECT  2.015 1.22 3.28 1.34 ;
      RECT  0.785 1.185 0.89 1.44 ;
      RECT  0.785 1.44 2.515 1.56 ;
  END
END SEN_NR4B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21_1
#      Description : "One 2-input OR into 2-input AND"
#      Equation    : X=(A1|A2)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21_1
  CLASS CORE ;
  FOREIGN SEN_OA21_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0486 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.075 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.83 1.43 0.95 1.75 ;
      RECT  1.08 1.43 1.2 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  1.13 0.05 1.25 0.385 ;
      RECT  0.35 0.05 0.47 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.3 1.5 0.5 ;
      RECT  1.35 0.5 1.45 1.29 ;
    END
    ANTENNADIFFAREA 0.185 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.37 0.195 0.49 ;
      RECT  0.075 0.49 0.74 0.59 ;
      RECT  0.62 0.37 0.74 0.49 ;
      RECT  0.84 0.49 1.245 0.59 ;
      RECT  1.155 0.59 1.245 1.22 ;
      RECT  0.555 1.22 1.245 1.34 ;
      RECT  0.555 1.34 0.675 1.44 ;
  END
END SEN_OA21_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21_2
#      Description : "One 2-input OR into 2-input AND"
#      Equation    : X=(A1|A2)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21_2
  CLASS CORE ;
  FOREIGN SEN_OA21_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0972 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.41 0.445 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.355 1.43 1.475 1.75 ;
      RECT  1.88 1.43 2.0 1.75 ;
      RECT  2.415 1.21 2.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.88 0.05 2.0 0.385 ;
      RECT  0.325 0.05 0.445 0.39 ;
      RECT  0.845 0.05 0.965 0.39 ;
      RECT  2.415 0.05 2.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.3 2.25 1.3 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.24 1.77 0.36 ;
      RECT  1.105 0.36 1.225 0.49 ;
      RECT  0.065 0.37 0.185 0.49 ;
      RECT  0.065 0.49 1.225 0.59 ;
      RECT  1.335 0.49 2.06 0.59 ;
      RECT  1.97 0.59 2.06 0.755 ;
      RECT  1.965 0.755 2.06 0.925 ;
      RECT  1.97 0.925 2.06 1.22 ;
      RECT  0.82 1.22 2.06 1.34 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.585 1.3 0.705 1.44 ;
      RECT  0.585 1.44 1.25 1.56 ;
  END
END SEN_OA21_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21_4
#      Description : "One 2-input OR into 2-input AND"
#      Equation    : X=(A1|A2)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21_4
  CLASS CORE ;
  FOREIGN SEN_OA21_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1941 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.41 0.455 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.855 1.41 0.975 1.75 ;
      RECT  2.67 1.41 2.79 1.75 ;
      RECT  3.195 1.41 3.315 1.75 ;
      RECT  3.46 1.21 3.58 1.75 ;
      RECT  4.04 1.21 4.16 1.75 ;
      RECT  4.6 1.21 4.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.335 0.05 0.455 0.385 ;
      RECT  0.855 0.05 0.975 0.39 ;
      RECT  1.375 0.05 1.495 0.39 ;
      RECT  1.895 0.05 2.015 0.39 ;
      RECT  4.015 0.05 4.185 0.515 ;
      RECT  3.46 0.05 3.58 0.59 ;
      RECT  4.6 0.05 4.72 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.74 0.31 3.86 0.605 ;
      RECT  3.74 0.605 4.46 0.695 ;
      RECT  4.34 0.31 4.46 0.605 ;
      RECT  4.35 0.695 4.46 1.005 ;
      RECT  3.74 1.005 4.46 1.105 ;
      RECT  3.74 1.105 3.86 1.3 ;
      RECT  4.34 1.105 4.46 1.3 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.155 0.24 3.34 0.36 ;
      RECT  2.155 0.36 2.275 0.48 ;
      RECT  0.075 0.37 0.195 0.48 ;
      RECT  0.075 0.48 2.275 0.59 ;
      RECT  2.385 0.46 3.33 0.58 ;
      RECT  3.23 0.58 3.33 0.785 ;
      RECT  3.23 0.785 4.25 0.895 ;
      RECT  3.23 0.895 3.33 1.21 ;
      RECT  1.345 1.21 3.33 1.32 ;
      RECT  0.075 1.21 1.235 1.31 ;
      RECT  0.075 1.31 0.195 1.43 ;
      RECT  1.115 1.31 1.235 1.44 ;
      RECT  1.115 1.44 2.33 1.56 ;
  END
END SEN_OA21_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21_8
#      Description : "One 2-input OR into 2-input AND"
#      Equation    : X=(A1|A2)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21_8
  CLASS CORE ;
  FOREIGN SEN_OA21_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.45 0.92 ;
      RECT  0.35 0.92 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4752 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.51 6.45 0.71 ;
      RECT  4.95 0.71 6.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4752 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.26 0.835 ;
      RECT  1.55 0.835 3.555 0.955 ;
      RECT  1.55 0.955 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.395 1.575 2.515 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  3.005 1.575 3.125 1.75 ;
      RECT  3.61 1.575 3.73 1.75 ;
      RECT  4.225 1.575 4.345 1.75 ;
      RECT  4.75 1.46 4.92 1.75 ;
      RECT  5.27 1.46 5.44 1.75 ;
      RECT  5.79 1.46 5.96 1.75 ;
      RECT  6.335 1.38 6.455 1.75 ;
      RECT  6.855 1.42 6.975 1.75 ;
      RECT  7.375 1.415 7.495 1.75 ;
      RECT  7.895 1.415 8.015 1.75 ;
      RECT  8.415 1.21 8.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  4.19 0.05 4.36 0.19 ;
      RECT  0.325 0.05 0.445 0.385 ;
      RECT  0.845 0.05 0.965 0.385 ;
      RECT  1.365 0.05 1.485 0.385 ;
      RECT  1.885 0.05 2.005 0.385 ;
      RECT  4.775 0.05 4.895 0.385 ;
      RECT  5.295 0.05 5.415 0.385 ;
      RECT  5.815 0.05 5.935 0.385 ;
      RECT  6.335 0.05 6.455 0.385 ;
      RECT  6.855 0.05 6.975 0.385 ;
      RECT  7.375 0.05 7.495 0.385 ;
      RECT  7.895 0.05 8.015 0.385 ;
      RECT  8.415 0.05 8.535 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.545 0.475 8.325 0.595 ;
      RECT  6.545 0.595 8.05 0.605 ;
      RECT  7.88 0.605 8.05 1.11 ;
      RECT  6.95 1.11 8.275 1.24 ;
      RECT  6.55 1.24 8.275 1.29 ;
      RECT  6.55 1.29 7.05 1.33 ;
      RECT  6.55 1.33 6.715 1.53 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.12 0.28 4.66 0.45 ;
      RECT  2.12 0.45 2.29 0.475 ;
      RECT  4.49 0.45 4.66 0.48 ;
      RECT  0.065 0.38 0.185 0.475 ;
      RECT  0.065 0.475 2.29 0.6 ;
      RECT  4.49 0.48 6.245 0.61 ;
      RECT  6.6 0.715 7.775 0.885 ;
      RECT  6.6 0.885 6.77 1.025 ;
      RECT  2.38 0.54 4.11 0.67 ;
      RECT  3.94 0.67 4.11 1.025 ;
      RECT  3.94 1.025 6.77 1.065 ;
      RECT  1.86 1.065 6.77 1.15 ;
      RECT  1.86 1.15 4.11 1.21 ;
      RECT  0.275 1.21 4.11 1.225 ;
      RECT  0.275 1.225 2.03 1.34 ;
      RECT  4.48 1.24 6.245 1.315 ;
      RECT  2.12 1.315 6.245 1.37 ;
      RECT  2.12 1.37 4.65 1.45 ;
      RECT  0.065 1.365 0.185 1.45 ;
      RECT  0.065 1.45 4.65 1.485 ;
      RECT  0.065 1.485 2.29 1.59 ;
  END
END SEN_OA21_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21B_0P5
#      Description : "One 2-input OR into 2-input AND (1 inverted input)"
#      Equation    : X=(A1|A2)&!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21B_0P5
  CLASS CORE ;
  FOREIGN SEN_OA21B_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.51 0.255 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.6 1.615 0.78 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.195 0.05 1.315 0.25 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  0.61 0.05 0.73 0.42 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.875 0.18 0.995 0.34 ;
      RECT  0.875 0.34 1.25 0.435 ;
      RECT  1.15 0.435 1.25 1.535 ;
    END
    ANTENNADIFFAREA 0.106 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.345 0.185 0.46 0.53 ;
      RECT  0.345 0.53 1.06 0.62 ;
      RECT  0.95 0.62 1.06 1.405 ;
      RECT  0.08 1.405 1.06 1.525 ;
      RECT  0.08 1.525 0.2 1.62 ;
  END
END SEN_OA21B_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21B_1
#      Description : "One 2-input OR into 2-input AND (1 inverted input)"
#      Equation    : X=(A1|A2)&!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21B_1
  CLASS CORE ;
  FOREIGN SEN_OA21B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.175 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.205 1.21 1.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.055 0.05 0.175 0.39 ;
      RECT  0.64 0.05 0.76 0.39 ;
      RECT  1.205 0.05 1.325 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.31 1.05 1.31 ;
      RECT  0.75 1.31 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.192 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.27 0.46 0.5 ;
      RECT  0.34 0.5 0.85 0.59 ;
      RECT  0.75 0.59 0.85 1.1 ;
      RECT  0.57 1.1 0.85 1.19 ;
      RECT  0.57 1.19 0.66 1.455 ;
      RECT  0.46 1.455 0.66 1.575 ;
  END
END SEN_OA21B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21B_2
#      Description : "One 2-input OR into 2-input AND (1 inverted input)"
#      Equation    : X=(A1|A2)&!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21B_2
  CLASS CORE ;
  FOREIGN SEN_OA21B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  2.15 1.41 2.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.07 0.05 0.19 0.39 ;
      RECT  0.59 0.05 0.71 0.39 ;
      RECT  1.11 0.05 1.23 0.39 ;
      RECT  1.37 0.05 1.49 0.39 ;
      RECT  1.89 0.05 2.01 0.39 ;
      RECT  2.41 0.05 2.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.54 0.495 2.3 0.615 ;
      RECT  1.54 0.615 2.05 0.69 ;
      RECT  1.95 0.69 2.05 1.0 ;
      RECT  1.55 1.0 2.05 1.12 ;
      RECT  1.55 1.12 1.655 1.3 ;
    END
    ANTENNADIFFAREA 0.308 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.33 0.27 0.45 0.5 ;
      RECT  0.33 0.5 1.245 0.59 ;
      RECT  0.85 0.27 0.97 0.5 ;
      RECT  1.155 0.59 1.245 0.785 ;
      RECT  1.155 0.785 1.77 0.895 ;
      RECT  1.155 0.895 1.245 1.21 ;
      RECT  0.825 1.21 1.245 1.33 ;
      RECT  0.07 1.21 0.715 1.32 ;
      RECT  0.07 1.32 0.19 1.43 ;
      RECT  0.585 1.32 0.715 1.44 ;
      RECT  0.585 1.44 1.255 1.56 ;
      RECT  1.89 1.21 2.53 1.32 ;
      RECT  2.41 1.32 2.53 1.43 ;
      RECT  1.89 1.32 2.01 1.44 ;
      RECT  1.345 1.44 2.01 1.56 ;
  END
END SEN_OA21B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21B_3
#      Description : "One 2-input OR into 2-input AND (1 inverted input)"
#      Equation    : X=(A1|A2)&!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21B_3
  CLASS CORE ;
  FOREIGN SEN_OA21B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.14 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.144 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.144 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.45 0.89 ;
      RECT  2.95 0.89 3.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.585 1.415 0.705 1.75 ;
      RECT  2.895 1.415 3.015 1.75 ;
      RECT  3.415 1.21 3.535 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.845 0.05 0.965 0.385 ;
      RECT  1.44 0.05 1.56 0.385 ;
      RECT  2.115 0.05 2.235 0.385 ;
      RECT  2.635 0.05 2.755 0.385 ;
      RECT  3.155 0.05 3.275 0.385 ;
      RECT  0.24 0.05 0.36 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.415 0.39 3.535 0.495 ;
      RECT  1.855 0.495 3.535 0.615 ;
      RECT  1.855 0.615 2.86 0.69 ;
      RECT  2.35 0.69 2.45 1.11 ;
      RECT  1.855 1.11 2.51 1.29 ;
    END
    ANTENNADIFFAREA 0.561 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.53 0.485 1.725 0.605 ;
      RECT  1.625 0.605 1.725 0.78 ;
      RECT  1.625 0.78 2.25 0.89 ;
      RECT  1.625 0.89 1.745 1.21 ;
      RECT  1.08 1.21 1.745 1.33 ;
      RECT  0.3 1.195 0.965 1.315 ;
      RECT  0.845 1.315 0.965 1.44 ;
      RECT  0.845 1.44 1.54 1.56 ;
      RECT  2.635 1.195 3.3 1.315 ;
      RECT  2.635 1.315 2.755 1.44 ;
      RECT  2.06 1.44 2.755 1.56 ;
  END
END SEN_OA21B_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21B_4
#      Description : "One 2-input OR into 2-input AND (1 inverted input)"
#      Equation    : X=(A1|A2)&!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21B_4
  CLASS CORE ;
  FOREIGN SEN_OA21B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.192 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.192 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.45 0.89 ;
      RECT  3.95 0.89 4.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.41 0.45 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.85 1.41 0.97 1.75 ;
      RECT  3.83 1.41 3.95 1.75 ;
      RECT  4.35 1.41 4.47 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.615 0.05 0.735 0.385 ;
      RECT  1.605 0.05 1.725 0.385 ;
      RECT  2.175 0.05 2.295 0.385 ;
      RECT  3.025 0.05 3.145 0.385 ;
      RECT  3.57 0.05 3.69 0.385 ;
      RECT  4.09 0.05 4.21 0.385 ;
      RECT  0.07 0.05 0.19 0.585 ;
      RECT  2.455 0.05 2.575 0.585 ;
      RECT  4.61 0.05 4.73 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.74 0.485 4.495 0.51 ;
      RECT  2.74 0.51 4.495 0.605 ;
      RECT  2.74 0.605 3.86 0.69 ;
      RECT  3.35 0.69 3.45 1.11 ;
      RECT  2.74 1.11 3.45 1.29 ;
    END
    ANTENNADIFFAREA 0.616 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.305 0.475 2.245 0.595 ;
      RECT  2.155 0.595 2.245 0.785 ;
      RECT  2.155 0.785 3.25 0.895 ;
      RECT  2.155 0.895 2.245 1.21 ;
      RECT  1.345 1.21 2.245 1.33 ;
      RECT  3.57 1.21 4.73 1.31 ;
      RECT  4.61 1.31 4.73 1.43 ;
      RECT  3.57 1.31 3.69 1.44 ;
      RECT  2.43 1.44 3.69 1.56 ;
      RECT  0.07 1.21 1.23 1.32 ;
      RECT  0.07 1.32 0.19 1.43 ;
      RECT  1.11 1.32 1.23 1.44 ;
      RECT  1.11 1.44 2.32 1.56 ;
  END
END SEN_OA21B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA21B_8
#      Description : "One 2-input OR into 2-input AND (1 inverted input)"
#      Equation    : X=(A1|A2)&!B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA21B_8
  CLASS CORE ;
  FOREIGN SEN_OA21B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.665 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2556 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2556 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  4.985 1.44 5.13 1.75 ;
      RECT  5.5 1.44 5.65 1.75 ;
      RECT  6.02 1.44 6.17 1.75 ;
      RECT  6.54 1.44 6.685 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  2.405 0.05 2.525 0.36 ;
      RECT  4.735 0.05 4.855 0.36 ;
      RECT  5.255 0.05 5.375 0.36 ;
      RECT  5.775 0.05 5.895 0.36 ;
      RECT  6.295 0.05 6.415 0.36 ;
      RECT  1.365 0.05 1.485 0.375 ;
      RECT  1.885 0.05 2.005 0.375 ;
      RECT  2.655 0.05 2.775 0.39 ;
      RECT  3.175 0.05 3.295 0.4 ;
      RECT  3.695 0.05 3.815 0.4 ;
      RECT  4.215 0.05 4.335 0.4 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  6.815 0.05 6.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.84 0.45 6.725 0.51 ;
      RECT  2.75 0.51 6.725 0.57 ;
      RECT  2.75 0.57 5.665 0.62 ;
      RECT  2.75 0.62 5.05 0.69 ;
      RECT  4.465 0.69 4.65 1.11 ;
      RECT  2.75 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.145 0.22 2.265 0.46 ;
      RECT  2.145 0.46 2.545 0.465 ;
      RECT  1.105 0.24 1.225 0.445 ;
      RECT  0.275 0.445 1.225 0.465 ;
      RECT  0.275 0.465 2.545 0.555 ;
      RECT  1.625 0.24 1.745 0.465 ;
      RECT  2.445 0.555 2.545 0.795 ;
      RECT  2.445 0.795 4.345 0.905 ;
      RECT  2.445 0.905 2.565 1.25 ;
      RECT  1.575 1.25 2.565 1.375 ;
      RECT  4.74 1.2 5.405 1.22 ;
      RECT  4.74 1.22 6.935 1.35 ;
      RECT  4.74 1.35 4.89 1.455 ;
      RECT  6.815 1.35 6.935 1.48 ;
      RECT  2.655 1.39 2.78 1.455 ;
      RECT  2.655 1.455 4.89 1.585 ;
      RECT  4.195 1.585 4.89 1.605 ;
      RECT  0.275 1.23 1.485 1.35 ;
      RECT  1.365 1.35 1.485 1.465 ;
      RECT  1.365 1.465 2.56 1.585 ;
  END
END SEN_OA21B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OA222_0P5
#      Description : "Three 2-input ORs into a 3-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)&(C1|C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA222_0P5
  CLASS CORE ;
  FOREIGN SEN_OA222_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.91 0.65 1.09 ;
      RECT  0.35 1.09 0.45 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.905 0.855 1.33 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  0.95 0.91 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.74 0.71 1.87 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0231 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.125 1.43 1.24 1.75 ;
      RECT  1.875 1.465 2.045 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  1.9 0.05 2.02 0.39 ;
      RECT  0.59 0.05 0.71 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.2 2.28 1.53 ;
    END
    ANTENNADIFFAREA 0.097 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.835 0.14 1.795 0.23 ;
      RECT  0.835 0.23 1.005 0.325 ;
      RECT  1.625 0.23 1.795 0.43 ;
      RECT  1.13 0.23 1.25 0.47 ;
      RECT  1.39 0.325 1.51 0.53 ;
      RECT  1.39 0.53 2.06 0.62 ;
      RECT  1.965 0.62 2.06 1.25 ;
      RECT  0.945 1.25 2.06 1.34 ;
      RECT  0.945 1.34 1.035 1.48 ;
      RECT  1.38 1.34 1.5 1.615 ;
      RECT  0.54 1.48 1.035 1.6 ;
      RECT  0.34 0.17 0.45 0.655 ;
      RECT  0.34 0.655 1.24 0.775 ;
      RECT  1.12 0.58 1.24 0.655 ;
  END
END SEN_OA222_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OA222_1
#      Description : "Three 2-input ORs into a 3-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)&(C1|C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA222_1
  CLASS CORE ;
  FOREIGN SEN_OA222_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.91 0.65 1.09 ;
      RECT  0.35 1.09 0.45 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.91 0.85 1.34 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 0.91 ;
      RECT  0.95 0.91 1.45 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.16 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.74 0.71 1.87 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0405 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.125 1.43 1.24 1.75 ;
      RECT  1.875 1.465 2.045 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.33 0.05 0.45 0.36 ;
      RECT  1.9 0.05 2.02 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.31 2.275 1.49 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.81 0.14 1.51 0.23 ;
      RECT  0.81 0.23 0.98 0.32 ;
      RECT  1.39 0.23 1.51 0.36 ;
      RECT  0.07 0.26 0.19 0.45 ;
      RECT  0.07 0.45 0.71 0.54 ;
      RECT  0.59 0.26 0.71 0.45 ;
      RECT  0.6 0.54 0.71 0.7 ;
      RECT  0.6 0.7 1.24 0.82 ;
      RECT  1.12 0.63 1.24 0.7 ;
      RECT  1.13 0.325 1.25 0.45 ;
      RECT  1.13 0.45 2.06 0.54 ;
      RECT  1.65 0.26 1.77 0.45 ;
      RECT  1.965 0.54 2.06 1.25 ;
      RECT  0.945 1.25 2.06 1.34 ;
      RECT  1.33 1.34 2.06 1.365 ;
      RECT  0.945 1.34 1.035 1.48 ;
      RECT  0.54 1.48 1.035 1.6 ;
  END
END SEN_OA222_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA222_2
#      Description : "Three 2-input ORs into a 3-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)&(C1|C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA222_2
  CLASS CORE ;
  FOREIGN SEN_OA222_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.655 0.89 ;
      RECT  0.55 0.89 0.655 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.695 1.25 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 0.71 ;
      RECT  1.35 0.71 1.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 0.71 ;
      RECT  1.75 0.71 2.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.34 0.695 2.655 0.89 ;
      RECT  2.55 0.89 2.655 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.44 0.45 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  1.405 1.48 1.575 1.75 ;
      RECT  2.715 1.465 2.885 1.75 ;
      RECT  3.07 1.175 3.19 1.75 ;
      RECT  3.6 1.41 3.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.56 0.05 0.73 0.32 ;
      RECT  2.81 0.05 2.98 0.335 ;
      RECT  3.355 0.05 3.475 0.38 ;
      RECT  0.06 0.05 0.2 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.095 0.3 3.25 0.5 ;
      RECT  3.095 0.5 3.74 0.535 ;
      RECT  3.565 0.34 3.74 0.5 ;
      RECT  3.095 0.535 3.65 0.69 ;
      RECT  3.55 0.69 3.65 1.11 ;
      RECT  3.35 1.11 3.65 1.29 ;
    END
    ANTENNADIFFAREA 0.228 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.08 0.14 2.42 0.23 ;
      RECT  1.08 0.23 1.25 0.32 ;
      RECT  2.25 0.23 2.42 0.32 ;
      RECT  1.75 0.23 1.87 0.375 ;
      RECT  0.325 0.175 0.445 0.41 ;
      RECT  0.325 0.41 1.51 0.425 ;
      RECT  0.845 0.175 0.965 0.41 ;
      RECT  1.34 0.32 1.51 0.41 ;
      RECT  0.355 0.425 1.43 0.515 ;
      RECT  1.985 0.32 2.16 0.41 ;
      RECT  1.985 0.41 2.65 0.43 ;
      RECT  2.53 0.21 2.65 0.41 ;
      RECT  1.985 0.43 2.925 0.52 ;
      RECT  2.835 0.52 2.925 0.78 ;
      RECT  2.835 0.78 3.45 0.89 ;
      RECT  2.835 0.89 2.925 1.255 ;
      RECT  0.94 1.12 2.02 1.21 ;
      RECT  0.94 1.21 1.03 1.255 ;
      RECT  1.93 1.21 2.02 1.255 ;
      RECT  0.91 1.255 1.03 1.465 ;
      RECT  1.93 1.255 2.925 1.375 ;
      RECT  0.065 1.26 0.705 1.35 ;
      RECT  0.585 1.35 0.705 1.515 ;
      RECT  0.065 1.35 0.185 1.525 ;
      RECT  1.17 1.3 1.805 1.39 ;
      RECT  1.17 1.39 1.29 1.52 ;
      RECT  1.69 1.39 1.805 1.61 ;
      RECT  1.895 1.465 2.61 1.585 ;
  END
END SEN_OA222_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA222_3
#      Description : "Three 2-input ORs into a 3-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)&(C1|C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA222_3
  CLASS CORE ;
  FOREIGN SEN_OA222_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.9 ;
      RECT  0.75 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.85 0.895 ;
      RECT  1.35 0.895 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.71 ;
      RECT  2.15 0.71 2.45 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.05 0.895 ;
      RECT  2.95 0.895 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.45 0.895 ;
      RECT  3.35 0.895 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.44 0.45 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  2.125 1.4 2.245 1.75 ;
      RECT  3.37 1.4 3.49 1.75 ;
      RECT  3.835 1.4 3.955 1.75 ;
      RECT  4.355 1.4 4.475 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  4.34 0.05 4.49 0.4 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  3.84 0.05 3.955 0.69 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.055 0.51 4.735 0.69 ;
      RECT  4.55 0.69 4.65 1.11 ;
      RECT  3.95 1.11 4.735 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.9 0.16 2.53 0.19 ;
      RECT  1.355 0.19 3.75 0.26 ;
      RECT  1.355 0.26 2.03 0.32 ;
      RECT  2.43 0.26 3.75 0.32 ;
      RECT  1.355 0.32 1.475 0.36 ;
      RECT  3.63 0.32 3.75 0.36 ;
      RECT  2.135 0.375 2.255 0.45 ;
      RECT  0.275 0.45 2.255 0.57 ;
      RECT  2.54 0.45 3.75 0.57 ;
      RECT  3.645 0.57 3.75 0.785 ;
      RECT  2.54 0.57 2.65 0.99 ;
      RECT  3.645 0.785 4.46 0.895 ;
      RECT  1.615 0.99 2.835 1.08 ;
      RECT  1.615 1.08 1.735 1.18 ;
      RECT  2.72 1.08 2.835 1.22 ;
      RECT  0.795 1.18 1.735 1.3 ;
      RECT  2.72 1.22 3.02 1.34 ;
      RECT  3.63 1.08 3.75 1.22 ;
      RECT  3.11 1.22 3.75 1.31 ;
      RECT  3.11 1.31 3.23 1.465 ;
      RECT  2.545 1.465 3.23 1.585 ;
      RECT  1.875 1.17 2.565 1.29 ;
      RECT  1.875 1.29 2.0 1.525 ;
      RECT  1.355 1.4 1.475 1.525 ;
      RECT  1.355 1.525 2.0 1.615 ;
      RECT  0.065 1.26 0.705 1.35 ;
      RECT  0.585 1.35 0.705 1.465 ;
      RECT  0.065 1.35 0.185 1.485 ;
      RECT  0.585 1.465 1.26 1.585 ;
  END
END SEN_OA222_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OA222_4
#      Description : "Three 2-input ORs into a 3-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)&(C1|C2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA222_4
  CLASS CORE ;
  FOREIGN SEN_OA222_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.895 ;
      RECT  0.15 0.895 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.895 ;
      RECT  1.35 0.895 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.71 ;
      RECT  1.95 0.71 2.45 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 2.65 0.71 ;
      RECT  2.55 0.71 3.05 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.85 0.895 ;
      RECT  3.75 0.895 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.4 0.445 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  2.135 1.44 2.255 1.75 ;
      RECT  3.43 1.435 3.55 1.75 ;
      RECT  3.94 1.215 4.06 1.75 ;
      RECT  4.46 1.4 4.58 1.75 ;
      RECT  4.99 1.21 5.11 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  3.94 0.05 4.07 0.36 ;
      RECT  1.105 0.05 1.225 0.4 ;
      RECT  4.46 0.05 4.58 0.4 ;
      RECT  0.585 0.05 0.705 0.41 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  4.99 0.05 5.11 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.51 4.85 0.69 ;
      RECT  4.75 0.69 4.85 1.11 ;
      RECT  4.15 1.11 4.85 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.33 0.215 3.835 0.335 ;
      RECT  2.135 0.435 2.255 0.5 ;
      RECT  0.275 0.5 2.255 0.62 ;
      RECT  2.86 0.455 4.06 0.575 ;
      RECT  3.94 0.575 4.06 0.785 ;
      RECT  3.165 0.575 3.255 1.0 ;
      RECT  3.94 0.785 4.64 0.895 ;
      RECT  1.615 1.0 3.255 1.12 ;
      RECT  1.615 1.12 1.735 1.22 ;
      RECT  0.795 1.22 1.735 1.34 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.585 1.3 0.705 1.455 ;
      RECT  0.065 1.3 0.185 1.5 ;
      RECT  0.585 1.455 1.25 1.575 ;
      RECT  1.875 1.21 2.57 1.33 ;
      RECT  1.875 1.33 1.995 1.48 ;
      RECT  1.355 1.43 1.475 1.48 ;
      RECT  1.355 1.48 1.995 1.6 ;
      RECT  3.17 1.21 3.84 1.33 ;
      RECT  3.17 1.33 3.29 1.44 ;
      RECT  2.59 1.44 3.29 1.56 ;
  END
END SEN_OA222_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_1
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_1
  CLASS CORE ;
  FOREIGN SEN_OA22_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.7 1.25 0.9 ;
      RECT  0.95 0.9 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.65 0.9 ;
      RECT  0.35 0.9 0.45 1.295 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0624 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.32 1.41 1.45 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.335 0.05 1.46 0.37 ;
      RECT  0.32 0.05 0.45 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.415 1.735 0.585 ;
      RECT  1.55 0.585 1.65 1.215 ;
      RECT  1.55 1.215 1.735 1.385 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.59 0.16 1.225 0.25 ;
      RECT  1.11 0.25 1.225 0.375 ;
      RECT  0.59 0.25 0.7 0.5 ;
      RECT  0.065 0.37 0.185 0.5 ;
      RECT  0.065 0.5 0.7 0.59 ;
      RECT  0.82 0.47 1.46 0.59 ;
      RECT  1.34 0.59 1.46 1.21 ;
      RECT  1.14 1.21 1.46 1.3 ;
      RECT  1.14 1.3 1.23 1.41 ;
      RECT  0.62 1.41 1.23 1.5 ;
      RECT  0.62 1.5 0.74 1.63 ;
  END
END SEN_OA22_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_2
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_2
  CLASS CORE ;
  FOREIGN SEN_OA22_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1248 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.42 0.44 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.96 1.47 2.13 1.75 ;
      RECT  2.5 1.41 2.63 1.75 ;
      RECT  3.02 1.41 3.15 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  2.5 0.05 2.63 0.36 ;
      RECT  3.02 0.05 3.145 0.38 ;
      RECT  0.31 0.05 0.44 0.39 ;
      RECT  0.83 0.05 0.96 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.74 0.51 3.05 0.69 ;
      RECT  2.95 0.69 3.05 1.11 ;
      RECT  2.735 1.11 3.05 1.295 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.13 0.2 2.39 0.32 ;
      RECT  1.13 0.32 1.25 0.49 ;
      RECT  0.06 0.17 0.175 0.49 ;
      RECT  0.06 0.49 1.25 0.595 ;
      RECT  1.36 0.47 2.65 0.575 ;
      RECT  1.36 0.575 1.91 0.58 ;
      RECT  2.56 0.575 2.65 0.79 ;
      RECT  1.81 0.58 1.91 1.075 ;
      RECT  2.56 0.79 2.84 0.89 ;
      RECT  1.365 1.075 1.91 1.17 ;
      RECT  1.365 1.17 1.46 1.475 ;
      RECT  0.78 1.475 1.46 1.575 ;
      RECT  0.055 1.22 1.255 1.33 ;
      RECT  0.055 1.33 0.18 1.63 ;
      RECT  1.55 1.275 2.41 1.38 ;
      RECT  1.55 1.38 1.65 1.5 ;
  END
END SEN_OA22_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_4
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_4
  CLASS CORE ;
  FOREIGN SEN_OA22_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2496 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.42 0.45 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.84 1.42 0.97 1.75 ;
      RECT  3.64 1.47 3.83 1.75 ;
      RECT  4.185 1.47 4.355 1.75 ;
      RECT  4.73 1.21 4.85 1.75 ;
      RECT  5.275 1.41 5.405 1.75 ;
      RECT  5.8 1.21 5.925 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.455 0.05 1.585 0.39 ;
      RECT  2.015 0.05 2.145 0.39 ;
      RECT  5.275 0.05 5.405 0.39 ;
      RECT  5.805 0.05 5.925 0.59 ;
      RECT  4.71 0.05 4.83 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.51 5.655 0.69 ;
      RECT  5.55 0.69 5.655 1.11 ;
      RECT  4.95 1.11 5.655 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.3 0.2 4.57 0.32 ;
      RECT  2.3 0.32 2.43 0.49 ;
      RECT  0.065 0.37 0.185 0.49 ;
      RECT  0.065 0.49 2.43 0.59 ;
      RECT  2.545 0.47 4.45 0.59 ;
      RECT  4.35 0.59 4.45 0.79 ;
      RECT  3.15 0.59 3.25 1.025 ;
      RECT  4.35 0.79 5.44 0.89 ;
      RECT  2.95 1.025 3.59 1.14 ;
      RECT  2.95 1.14 3.04 1.215 ;
      RECT  2.385 1.215 3.04 1.33 ;
      RECT  2.385 1.33 2.5 1.455 ;
      RECT  1.31 1.455 2.5 1.58 ;
      RECT  0.065 1.21 2.29 1.33 ;
      RECT  0.065 1.33 0.185 1.43 ;
      RECT  3.155 1.245 4.615 1.37 ;
      RECT  3.155 1.37 3.27 1.455 ;
      RECT  2.61 1.455 3.27 1.59 ;
  END
END SEN_OA22_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_6
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_6
  CLASS CORE ;
  FOREIGN SEN_OA22_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.05 0.89 ;
      RECT  5.95 0.89 6.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.85 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.25 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.415 0.44 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  0.83 1.415 0.96 1.75 ;
      RECT  1.35 1.44 1.48 1.75 ;
      RECT  5.08 1.48 5.25 1.75 ;
      RECT  5.62 1.42 5.75 1.75 ;
      RECT  6.14 1.42 6.27 1.75 ;
      RECT  6.665 1.21 6.785 1.75 ;
      RECT  7.18 1.41 7.31 1.75 ;
      RECT  7.7 1.41 7.83 1.75 ;
      RECT  8.22 1.41 8.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  0.31 0.05 0.44 0.39 ;
      RECT  0.83 0.05 0.96 0.39 ;
      RECT  1.35 0.05 1.48 0.39 ;
      RECT  1.87 0.05 2.0 0.39 ;
      RECT  2.39 0.05 2.52 0.39 ;
      RECT  2.91 0.05 3.04 0.39 ;
      RECT  7.18 0.05 7.31 0.39 ;
      RECT  7.7 0.05 7.83 0.39 ;
      RECT  8.225 0.05 8.345 0.39 ;
      RECT  6.68 0.05 6.785 0.69 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.9 0.51 8.08 0.69 ;
      RECT  7.95 0.69 8.08 1.11 ;
      RECT  6.925 1.11 8.08 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.25 0.19 6.585 0.32 ;
      RECT  6.495 0.32 6.585 0.36 ;
      RECT  3.25 0.32 3.42 0.48 ;
      RECT  0.055 0.17 0.175 0.48 ;
      RECT  0.055 0.48 3.42 0.59 ;
      RECT  3.57 0.41 6.37 0.54 ;
      RECT  6.245 0.54 6.37 0.79 ;
      RECT  4.62 0.54 4.755 1.03 ;
      RECT  6.245 0.79 7.81 0.89 ;
      RECT  4.62 1.03 5.09 1.16 ;
      RECT  4.62 1.16 4.755 1.185 ;
      RECT  3.37 1.185 4.755 1.315 ;
      RECT  3.37 1.315 3.5 1.44 ;
      RECT  1.82 1.44 3.5 1.58 ;
      RECT  3.37 1.58 3.5 1.63 ;
      RECT  3.175 1.155 3.28 1.195 ;
      RECT  0.055 1.195 3.28 1.325 ;
      RECT  0.055 1.325 0.175 1.62 ;
      RECT  5.36 1.2 6.55 1.26 ;
      RECT  4.845 1.26 6.55 1.33 ;
      RECT  4.845 1.33 5.49 1.385 ;
      RECT  4.845 1.385 4.975 1.46 ;
      RECT  3.595 1.46 4.975 1.595 ;
  END
END SEN_OA22_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_DG_1
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_DG_1
  CLASS CORE ;
  FOREIGN SEN_OA22_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.815 ;
      RECT  0.675 0.815 0.85 0.985 ;
      RECT  0.75 0.985 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.815 0.525 1.09 ;
      RECT  0.35 1.09 0.45 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.32 1.19 1.44 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.325 0.05 0.445 0.405 ;
      RECT  1.355 0.05 1.475 0.435 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.615 0.335 1.735 0.51 ;
      RECT  1.55 0.51 1.735 0.6 ;
      RECT  1.55 0.6 1.65 1.31 ;
      RECT  1.55 1.31 1.735 1.49 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.14 1.225 0.23 ;
      RECT  1.105 0.23 1.225 0.415 ;
      RECT  0.585 0.23 0.705 0.5 ;
      RECT  0.065 0.195 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.59 ;
      RECT  0.82 0.32 0.99 0.505 ;
      RECT  0.82 0.505 1.23 0.595 ;
      RECT  1.14 0.595 1.23 0.785 ;
      RECT  1.14 0.785 1.43 0.895 ;
      RECT  1.14 0.895 1.23 1.495 ;
      RECT  0.54 1.495 1.23 1.585 ;
  END
END SEN_OA22_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_DG_2
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_DG_2
  CLASS CORE ;
  FOREIGN SEN_OA22_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.8 ;
      RECT  0.69 0.8 0.85 0.99 ;
      RECT  0.75 0.99 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.525 0.98 ;
      RECT  0.35 0.98 0.45 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.32 1.2 1.425 1.75 ;
      RECT  1.81 1.41 1.945 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  1.81 0.05 1.945 0.39 ;
      RECT  0.325 0.05 0.445 0.405 ;
      RECT  1.32 0.05 1.425 0.68 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.31 1.685 1.49 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.14 1.23 0.23 ;
      RECT  1.11 0.23 1.23 0.415 ;
      RECT  0.585 0.23 0.705 0.5 ;
      RECT  0.065 0.225 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.59 ;
      RECT  0.82 0.32 0.99 0.505 ;
      RECT  0.82 0.505 1.23 0.595 ;
      RECT  1.14 0.595 1.23 0.785 ;
      RECT  1.14 0.785 1.46 0.895 ;
      RECT  1.14 0.895 1.23 1.48 ;
      RECT  0.54 1.48 1.23 1.6 ;
  END
END SEN_OA22_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_DG_4
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_DG_4
  CLASS CORE ;
  FOREIGN SEN_OA22_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.705 0.71 0.85 0.93 ;
      RECT  0.75 0.93 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.575 0.89 ;
      RECT  0.35 0.89 0.45 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.32 1.195 1.44 1.75 ;
      RECT  1.875 1.4 1.995 1.75 ;
      RECT  2.4 1.21 2.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.875 0.05 1.995 0.4 ;
      RECT  0.325 0.05 0.445 0.405 ;
      RECT  2.4 0.05 2.52 0.59 ;
      RECT  1.355 0.05 1.475 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.615 0.51 2.25 0.69 ;
      RECT  2.15 0.69 2.25 1.11 ;
      RECT  1.615 1.11 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.14 1.225 0.23 ;
      RECT  1.105 0.23 1.225 0.415 ;
      RECT  0.585 0.23 0.705 0.5 ;
      RECT  0.065 0.35 0.185 0.5 ;
      RECT  0.065 0.5 0.705 0.59 ;
      RECT  0.845 0.35 0.965 0.505 ;
      RECT  0.845 0.505 1.23 0.595 ;
      RECT  1.14 0.595 1.23 0.785 ;
      RECT  1.14 0.785 2.055 0.895 ;
      RECT  1.14 0.895 1.23 1.48 ;
      RECT  0.54 1.48 1.23 1.6 ;
  END
END SEN_OA22_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_DG_8
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_DG_8
  CLASS CORE ;
  FOREIGN SEN_OA22_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.42 0.445 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  2.155 1.4 2.275 1.75 ;
      RECT  2.665 1.185 2.785 1.75 ;
      RECT  3.185 1.4 3.305 1.75 ;
      RECT  3.705 1.4 3.825 1.75 ;
      RECT  4.225 1.4 4.345 1.75 ;
      RECT  4.76 1.21 4.88 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.325 0.05 0.445 0.395 ;
      RECT  0.84 0.05 0.965 0.395 ;
      RECT  3.185 0.05 3.305 0.4 ;
      RECT  3.705 0.05 3.825 0.4 ;
      RECT  4.225 0.05 4.345 0.4 ;
      RECT  4.76 0.05 4.88 0.59 ;
      RECT  2.665 0.05 2.785 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.925 0.51 4.65 0.69 ;
      RECT  4.48 0.69 4.65 1.11 ;
      RECT  2.925 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.215 2.325 0.335 ;
      RECT  1.105 0.335 1.225 0.485 ;
      RECT  0.065 0.36 0.185 0.485 ;
      RECT  0.065 0.485 1.225 0.605 ;
      RECT  1.35 0.49 2.56 0.61 ;
      RECT  2.47 0.61 2.56 0.795 ;
      RECT  1.35 0.61 1.45 1.19 ;
      RECT  2.47 0.795 4.255 0.885 ;
      RECT  0.82 1.19 1.805 1.315 ;
      RECT  0.065 1.18 0.73 1.3 ;
      RECT  0.065 1.3 0.185 1.42 ;
      RECT  0.61 1.3 0.73 1.455 ;
      RECT  0.61 1.455 1.25 1.575 ;
      RECT  1.895 1.185 2.56 1.305 ;
      RECT  1.895 1.305 2.015 1.48 ;
      RECT  1.345 1.48 2.015 1.6 ;
  END
END SEN_OA22_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OA22_8
#      Description : "Two 2-input ORs into 2-input AND"
#      Equation    : X=(A1|A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA22_8
  CLASS CORE ;
  FOREIGN SEN_OA22_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 5.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4536 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.71 7.05 0.89 ;
      RECT  5.95 0.89 6.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4536 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 3.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4536 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.65 0.9 ;
      RECT  0.55 0.9 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4536 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.2 0.185 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  0.585 1.44 0.705 1.75 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  1.625 1.44 1.745 1.75 ;
      RECT  5.785 1.44 5.905 1.75 ;
      RECT  6.305 1.44 6.425 1.75 ;
      RECT  6.825 1.44 6.945 1.75 ;
      RECT  7.44 1.2 7.56 1.75 ;
      RECT  8.05 1.4 8.17 1.75 ;
      RECT  8.57 1.4 8.69 1.75 ;
      RECT  9.09 1.4 9.21 1.75 ;
      RECT  9.61 1.205 9.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  1.885 0.05 2.005 0.36 ;
      RECT  2.405 0.05 2.525 0.36 ;
      RECT  2.925 0.05 3.045 0.36 ;
      RECT  3.445 0.05 3.565 0.36 ;
      RECT  8.05 0.05 8.17 0.38 ;
      RECT  8.57 0.05 8.69 0.38 ;
      RECT  9.09 0.05 9.21 0.38 ;
      RECT  9.61 0.05 9.73 0.595 ;
      RECT  7.545 0.05 7.65 0.695 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.51 9.48 0.69 ;
      RECT  9.31 0.69 9.48 1.11 ;
      RECT  7.75 1.11 9.48 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.66 0.19 7.455 0.36 ;
      RECT  3.66 0.36 3.83 0.45 ;
      RECT  0.065 0.45 3.83 0.62 ;
      RECT  3.965 0.45 7.42 0.62 ;
      RECT  7.25 0.62 7.42 0.815 ;
      RECT  5.215 0.62 5.385 1.18 ;
      RECT  7.25 0.815 9.145 0.95 ;
      RECT  2.145 1.18 5.385 1.35 ;
      RECT  0.325 1.18 2.025 1.35 ;
      RECT  1.855 1.35 2.025 1.455 ;
      RECT  1.855 1.455 3.565 1.625 ;
      RECT  5.52 1.18 7.205 1.35 ;
      RECT  5.52 1.35 5.69 1.455 ;
      RECT  3.965 1.455 5.69 1.625 ;
  END
END SEN_OA22_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_0P5
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_0P5
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.085 0.97 ;
      RECT  0.95 0.97 1.05 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.71 0.65 0.965 ;
      RECT  0.55 0.965 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.024 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.57 1.41 0.72 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.105 1.44 1.225 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.585 0.05 0.705 0.385 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  1.54 0.05 1.66 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.045 0.24 1.45 0.36 ;
      RECT  1.355 0.36 1.45 0.48 ;
      RECT  1.355 0.48 1.65 0.57 ;
      RECT  1.55 0.57 1.65 1.31 ;
      RECT  1.55 1.31 1.725 1.49 ;
    END
    ANTENNADIFFAREA 0.096 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.17 0.445 0.475 ;
      RECT  0.34 0.475 1.265 0.565 ;
      RECT  1.175 0.565 1.265 0.785 ;
      RECT  0.34 0.565 0.43 1.41 ;
      RECT  1.175 0.785 1.45 0.895 ;
      RECT  0.07 1.41 0.43 1.5 ;
      RECT  0.07 1.5 0.185 1.63 ;
      RECT  0.845 1.24 1.46 1.35 ;
      RECT  0.845 1.35 0.96 1.53 ;
      RECT  1.355 1.35 1.46 1.53 ;
  END
END SEN_OA2BB2_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_1
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_1
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.14 0.71 1.255 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.86 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.525 0.71 0.65 1.335 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.56 1.495 0.73 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.1 1.44 1.23 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  1.52 0.05 1.73 0.19 ;
      RECT  0.58 0.05 0.71 0.38 ;
      RECT  0.065 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.28 1.65 0.38 ;
      RECT  1.55 0.38 1.65 1.215 ;
      RECT  1.55 1.215 1.73 1.385 ;
    END
    ANTENNADIFFAREA 0.238 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.395 0.43 0.47 ;
      RECT  0.34 0.47 1.46 0.56 ;
      RECT  1.345 0.56 1.46 0.935 ;
      RECT  0.34 0.56 0.43 1.41 ;
      RECT  0.065 1.41 0.43 1.5 ;
      RECT  0.065 1.5 0.185 1.63 ;
      RECT  0.79 1.25 1.46 1.35 ;
      RECT  1.355 1.35 1.46 1.47 ;
  END
END SEN_OA2BB2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_2
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_2
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.05 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.415 0.465 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  2.215 1.415 2.35 1.75 ;
      RECT  2.75 1.415 2.88 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.635 0.05 0.765 0.345 ;
      RECT  1.18 0.05 1.31 0.345 ;
      RECT  0.065 0.05 0.19 0.39 ;
      RECT  1.705 0.05 1.835 0.39 ;
      RECT  2.75 0.05 2.88 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.42 0.48 2.39 0.585 ;
      RECT  1.42 0.585 1.85 0.69 ;
      RECT  1.75 0.69 1.85 1.11 ;
      RECT  1.55 1.11 1.85 1.295 ;
    END
    ANTENNADIFFAREA 0.322 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.955 0.185 2.61 0.275 ;
      RECT  1.955 0.275 2.07 0.39 ;
      RECT  2.5 0.275 2.61 0.5 ;
      RECT  2.5 0.5 3.135 0.59 ;
      RECT  3.015 0.37 3.135 0.5 ;
      RECT  0.29 0.435 1.29 0.54 ;
      RECT  1.2 0.54 1.29 0.785 ;
      RECT  1.2 0.785 1.64 0.895 ;
      RECT  1.2 0.895 1.29 1.035 ;
      RECT  0.94 1.035 1.29 1.125 ;
      RECT  0.94 1.125 1.05 1.285 ;
      RECT  0.065 1.21 0.765 1.3 ;
      RECT  0.635 1.3 0.765 1.415 ;
      RECT  0.065 1.3 0.19 1.43 ;
      RECT  0.635 1.415 1.31 1.505 ;
      RECT  1.185 1.28 1.31 1.415 ;
      RECT  1.95 1.21 3.135 1.315 ;
      RECT  3.015 1.315 3.135 1.43 ;
      RECT  1.95 1.315 2.08 1.46 ;
      RECT  1.41 1.46 2.08 1.58 ;
  END
END SEN_OA2BB2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_3
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_3
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.895 ;
      RECT  2.75 0.895 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 4.05 0.9 ;
      RECT  3.55 0.9 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.465 0.905 ;
      RECT  0.95 0.905 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1221 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.65 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1221 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.055 1.41 0.19 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  0.575 1.4 0.695 1.75 ;
      RECT  2.905 1.45 3.025 1.75 ;
      RECT  3.425 1.45 3.545 1.75 ;
      RECT  3.945 1.45 4.065 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.905 0.05 1.09 0.32 ;
      RECT  1.71 0.05 1.88 0.32 ;
      RECT  3.685 0.05 3.805 0.35 ;
      RECT  2.385 0.05 2.505 0.385 ;
      RECT  0.27 0.05 0.41 0.39 ;
      RECT  4.21 0.05 4.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.03 0.51 3.335 0.62 ;
      RECT  2.03 0.62 2.65 0.69 ;
      RECT  2.35 0.69 2.45 1.11 ;
      RECT  1.865 1.11 2.505 1.29 ;
    END
    ANTENNADIFFAREA 0.504 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.85 0.24 3.57 0.36 ;
      RECT  3.45 0.36 3.57 0.44 ;
      RECT  3.45 0.44 4.115 0.56 ;
      RECT  0.525 0.42 1.735 0.53 ;
      RECT  1.615 0.53 1.735 0.78 ;
      RECT  1.615 0.78 2.245 0.89 ;
      RECT  1.615 0.89 1.735 1.22 ;
      RECT  1.07 1.22 1.735 1.33 ;
      RECT  0.315 1.205 0.955 1.295 ;
      RECT  0.835 1.295 0.955 1.465 ;
      RECT  0.315 1.295 0.435 1.57 ;
      RECT  0.835 1.465 1.54 1.585 ;
      RECT  2.64 1.245 4.33 1.355 ;
      RECT  2.64 1.355 2.76 1.445 ;
      RECT  4.21 1.355 4.33 1.51 ;
      RECT  2.05 1.445 2.76 1.555 ;
  END
END SEN_OA2BB2_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_4
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_4
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.45 0.89 ;
      RECT  5.35 0.89 5.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2253 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2253 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.42 0.45 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.84 1.42 0.97 1.75 ;
      RECT  3.735 1.42 3.865 1.75 ;
      RECT  4.275 1.42 4.405 1.75 ;
      RECT  4.795 1.44 4.925 1.75 ;
      RECT  5.335 1.42 5.465 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  0.58 0.05 0.71 0.345 ;
      RECT  1.1 0.05 1.23 0.345 ;
      RECT  1.65 0.05 1.78 0.345 ;
      RECT  4.795 0.05 4.925 0.36 ;
      RECT  5.335 0.05 5.465 0.36 ;
      RECT  2.69 0.05 2.82 0.38 ;
      RECT  3.21 0.05 3.34 0.38 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  2.175 0.05 2.295 0.565 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.47 4.425 0.57 ;
      RECT  3.15 0.57 3.25 1.11 ;
      RECT  2.685 1.11 3.325 1.29 ;
    END
    ANTENNADIFFAREA 0.632 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.43 0.22 4.665 0.325 ;
      RECT  4.54 0.325 4.665 0.46 ;
      RECT  4.54 0.46 5.735 0.58 ;
      RECT  5.615 0.36 5.735 0.46 ;
      RECT  0.29 0.435 2.08 0.535 ;
      RECT  1.96 0.535 2.08 0.78 ;
      RECT  1.96 0.78 3.04 0.895 ;
      RECT  1.96 0.895 2.08 1.21 ;
      RECT  1.37 1.21 2.08 1.31 ;
      RECT  0.06 1.21 1.235 1.33 ;
      RECT  0.06 1.33 0.19 1.43 ;
      RECT  1.125 1.33 1.235 1.45 ;
      RECT  1.125 1.45 2.32 1.56 ;
      RECT  3.46 1.21 5.735 1.33 ;
      RECT  5.615 1.33 5.735 1.43 ;
      RECT  3.46 1.33 3.59 1.465 ;
      RECT  2.425 1.35 2.545 1.465 ;
      RECT  2.425 1.465 3.59 1.575 ;
  END
END SEN_OA2BB2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_8
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_8
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.71 7.485 0.92 ;
      RECT  6.55 0.92 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.41 0.71 9.45 0.925 ;
      RECT  9.35 0.925 9.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.705 2.575 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3258 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.25 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3258 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.48 0.47 1.75 ;
      RECT  0.0 1.75 9.8 1.85 ;
      RECT  0.82 1.48 0.99 1.75 ;
      RECT  1.34 1.48 1.51 1.75 ;
      RECT  5.685 1.48 5.855 1.75 ;
      RECT  6.205 1.48 6.385 1.75 ;
      RECT  6.725 1.48 6.895 1.75 ;
      RECT  7.245 1.48 7.415 1.75 ;
      RECT  7.765 1.48 7.935 1.75 ;
      RECT  8.285 1.48 8.455 1.75 ;
      RECT  8.81 1.46 8.98 1.75 ;
      RECT  9.33 1.49 9.5 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      RECT  0.82 0.05 0.99 0.31 ;
      RECT  1.34 0.05 1.51 0.31 ;
      RECT  1.86 0.05 2.03 0.31 ;
      RECT  2.38 0.05 2.55 0.31 ;
      RECT  4.14 0.05 4.31 0.315 ;
      RECT  3.62 0.05 3.79 0.32 ;
      RECT  4.675 0.05 4.845 0.32 ;
      RECT  7.765 0.05 7.935 0.32 ;
      RECT  8.285 0.05 8.46 0.32 ;
      RECT  8.81 0.05 8.98 0.32 ;
      RECT  9.33 0.05 9.5 0.32 ;
      RECT  5.215 0.05 5.335 0.4 ;
      RECT  0.24 0.05 0.36 0.59 ;
      RECT  3.025 0.05 3.145 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.31 3.505 0.415 ;
      RECT  3.35 0.415 5.11 0.51 ;
      RECT  3.35 0.51 7.395 0.585 ;
      RECT  5.675 0.42 7.395 0.51 ;
      RECT  4.95 0.585 7.395 0.59 ;
      RECT  4.35 0.585 4.65 1.11 ;
      RECT  4.95 0.59 5.85 0.69 ;
      RECT  3.63 1.11 5.31 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.45 0.16 7.675 0.33 ;
      RECT  5.45 0.33 5.57 0.4 ;
      RECT  7.505 0.33 7.675 0.42 ;
      RECT  7.505 0.42 9.735 0.59 ;
      RECT  0.545 0.4 2.875 0.575 ;
      RECT  2.7 0.575 2.875 0.775 ;
      RECT  2.7 0.775 4.25 0.89 ;
      RECT  2.7 0.89 2.87 1.21 ;
      RECT  1.885 1.21 3.045 1.38 ;
      RECT  5.425 1.2 9.735 1.37 ;
      RECT  5.425 1.37 5.595 1.47 ;
      RECT  3.385 0.99 3.49 1.47 ;
      RECT  3.385 1.47 5.595 1.64 ;
      RECT  0.065 1.22 1.77 1.39 ;
      RECT  1.6 1.39 1.77 1.47 ;
      RECT  1.6 1.47 3.29 1.64 ;
      RECT  3.185 1.38 3.29 1.47 ;
  END
END SEN_OA2BB2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_DG_1
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_DG_1
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.085 0.925 ;
      RECT  0.95 0.925 1.05 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.71 0.65 0.955 ;
      RECT  0.55 0.955 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.105 1.44 1.225 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.06 0.05 0.2 0.39 ;
      RECT  0.585 0.05 0.705 0.39 ;
      RECT  1.54 0.05 1.66 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.185 0.24 1.45 0.36 ;
      RECT  1.355 0.36 1.45 0.5 ;
      RECT  1.355 0.5 1.65 0.59 ;
      RECT  1.55 0.59 1.65 1.11 ;
      RECT  1.55 1.11 1.735 1.29 ;
    END
    ANTENNADIFFAREA 0.276 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.2 0.445 0.485 ;
      RECT  0.34 0.485 1.265 0.575 ;
      RECT  1.175 0.575 1.265 0.785 ;
      RECT  0.34 0.575 0.43 1.41 ;
      RECT  1.175 0.785 1.45 0.895 ;
      RECT  0.065 1.41 0.43 1.5 ;
      RECT  0.065 1.5 0.185 1.63 ;
      RECT  0.79 1.24 1.46 1.35 ;
      RECT  1.355 1.35 1.46 1.46 ;
  END
END SEN_OA2BB2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_DG_2
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_DG_2
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.9 ;
      RECT  1.55 0.9 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.9 ;
      RECT  1.95 0.9 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.95 ;
      RECT  0.35 0.95 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.63 1.45 1.75 1.75 ;
      RECT  2.15 1.45 2.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.585 0.05 0.705 0.355 ;
      RECT  1.13 0.05 1.24 0.385 ;
      RECT  2.15 0.05 2.27 0.385 ;
      RECT  0.06 0.05 0.2 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.795 0.215 1.04 0.335 ;
      RECT  0.95 0.335 1.04 0.48 ;
      RECT  0.95 0.48 1.8 0.59 ;
      RECT  0.95 0.59 1.05 1.11 ;
      RECT  0.95 1.11 1.265 1.29 ;
    END
    ANTENNADIFFAREA 0.32 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.345 0.215 2.035 0.34 ;
      RECT  1.915 0.34 2.035 0.475 ;
      RECT  1.915 0.475 2.53 0.595 ;
      RECT  2.41 0.335 2.53 0.475 ;
      RECT  0.325 0.205 0.445 0.445 ;
      RECT  0.325 0.445 0.855 0.555 ;
      RECT  0.745 0.555 0.855 1.25 ;
      RECT  0.585 1.25 0.855 1.34 ;
      RECT  0.585 1.34 0.705 1.53 ;
      RECT  1.37 1.24 2.53 1.36 ;
      RECT  1.37 1.36 1.49 1.44 ;
      RECT  2.405 1.36 2.53 1.48 ;
      RECT  0.81 1.44 1.49 1.56 ;
  END
END SEN_OA2BB2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_DG_3
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_DG_3
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.15 0.895 ;
      RECT  1.75 0.895 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.95 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.535 1.41 0.665 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  1.825 1.42 1.945 1.75 ;
      RECT  2.345 1.42 2.465 1.75 ;
      RECT  2.865 1.42 2.985 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.785 0.05 0.905 0.345 ;
      RECT  2.605 0.05 2.725 0.375 ;
      RECT  0.11 0.05 0.25 0.39 ;
      RECT  1.305 0.05 1.425 0.4 ;
      RECT  3.14 0.05 3.26 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 2.255 0.62 ;
      RECT  0.95 0.62 1.65 0.69 ;
      RECT  1.35 0.69 1.45 1.11 ;
      RECT  0.75 1.11 1.45 1.29 ;
    END
    ANTENNADIFFAREA 0.504 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.765 0.24 2.49 0.36 ;
      RECT  2.37 0.36 2.49 0.465 ;
      RECT  2.37 0.465 3.035 0.585 ;
      RECT  0.35 0.435 0.86 0.555 ;
      RECT  0.75 0.555 0.86 0.785 ;
      RECT  0.35 0.555 0.45 1.25 ;
      RECT  0.75 0.785 1.26 0.895 ;
      RECT  0.065 1.25 0.45 1.35 ;
      RECT  0.065 1.35 0.185 1.47 ;
      RECT  1.57 1.215 3.245 1.325 ;
      RECT  1.57 1.325 1.68 1.445 ;
      RECT  3.125 1.325 3.245 1.51 ;
      RECT  0.99 1.445 1.68 1.555 ;
  END
END SEN_OA2BB2_DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_DG_4
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_DG_4
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.65 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.65 0.89 ;
      RECT  3.55 0.89 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.505 0.925 ;
      RECT  0.35 0.925 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.675 0.25 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.215 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  2.135 1.41 2.255 1.75 ;
      RECT  2.655 1.41 2.775 1.75 ;
      RECT  3.175 1.41 3.295 1.75 ;
      RECT  3.695 1.41 3.815 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  3.175 0.05 3.295 0.35 ;
      RECT  3.695 0.05 3.815 0.35 ;
      RECT  1.105 0.05 1.225 0.36 ;
      RECT  1.625 0.05 1.745 0.4 ;
      RECT  0.065 0.05 0.185 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.45 2.825 0.51 ;
      RECT  0.795 0.51 2.825 0.55 ;
      RECT  0.795 0.55 2.05 0.69 ;
      RECT  1.55 0.69 1.65 1.11 ;
      RECT  1.055 1.11 1.65 1.115 ;
      RECT  1.055 1.115 1.735 1.29 ;
    END
    ANTENNADIFFAREA 0.624 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.835 0.24 3.035 0.36 ;
      RECT  2.915 0.36 3.035 0.44 ;
      RECT  2.915 0.44 4.075 0.56 ;
      RECT  3.955 0.32 4.075 0.44 ;
      RECT  0.275 0.445 0.685 0.555 ;
      RECT  0.595 0.555 0.685 0.78 ;
      RECT  0.595 0.78 1.4 0.89 ;
      RECT  0.595 0.89 0.695 1.37 ;
      RECT  1.875 1.2 4.075 1.32 ;
      RECT  1.875 1.32 1.995 1.44 ;
      RECT  3.955 1.32 4.075 1.475 ;
      RECT  0.785 1.44 1.995 1.56 ;
  END
END SEN_OA2BB2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA2BB2_DG_8
#      Description : "One 2-input OR with inverted inputs + 2-input OR into 2-input AND"
#      Equation    : X=(!A1|!A2)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA2BB2_DG_8
  CLASS CORE ;
  FOREIGN SEN_OA2BB2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 5.45 0.895 ;
      RECT  5.35 0.895 5.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 7.25 0.895 ;
      RECT  7.15 0.895 7.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.9 ;
      RECT  0.75 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.45 0.445 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  3.695 1.44 3.815 1.75 ;
      RECT  4.215 1.44 4.335 1.75 ;
      RECT  4.735 1.44 4.855 1.75 ;
      RECT  5.255 1.44 5.375 1.75 ;
      RECT  5.775 1.44 5.895 1.75 ;
      RECT  6.295 1.44 6.415 1.75 ;
      RECT  6.815 1.44 6.935 1.75 ;
      RECT  7.335 1.44 7.455 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  5.75 0.05 5.92 0.34 ;
      RECT  6.27 0.05 6.44 0.34 ;
      RECT  6.79 0.05 6.96 0.34 ;
      RECT  7.31 0.05 7.48 0.34 ;
      RECT  0.585 0.05 0.705 0.35 ;
      RECT  1.105 0.05 1.225 0.35 ;
      RECT  1.625 0.05 1.745 0.4 ;
      RECT  2.145 0.05 2.265 0.4 ;
      RECT  2.665 0.05 2.785 0.4 ;
      RECT  3.185 0.05 3.305 0.4 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.49 5.4 0.51 ;
      RECT  1.35 0.51 5.4 0.6 ;
      RECT  1.35 0.6 4.25 0.69 ;
      RECT  3.15 0.69 3.32 1.11 ;
      RECT  1.55 1.11 3.32 1.29 ;
    END
    ANTENNADIFFAREA 1.248 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.45 0.21 5.66 0.38 ;
      RECT  5.49 0.38 5.66 0.43 ;
      RECT  5.49 0.43 7.715 0.6 ;
      RECT  0.275 0.44 1.26 0.56 ;
      RECT  1.14 0.56 1.26 0.785 ;
      RECT  1.14 0.785 2.885 0.895 ;
      RECT  1.14 0.895 1.26 1.245 ;
      RECT  0.795 1.245 1.26 1.355 ;
      RECT  3.41 1.18 7.715 1.35 ;
      RECT  3.41 1.35 3.58 1.415 ;
      RECT  1.355 1.415 3.58 1.585 ;
      RECT  0.065 1.245 0.705 1.355 ;
      RECT  0.585 1.355 0.705 1.445 ;
      RECT  0.065 1.355 0.185 1.47 ;
      RECT  0.585 1.445 1.25 1.555 ;
  END
END SEN_OA2BB2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OA31_0P5
#      Description : "One 3-input OR into 2-input AND"
#      Equation    : X=(A1|A2|A3)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA31_0P5
  CLASS CORE ;
  FOREIGN SEN_OA31_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.05 0.71 1.25 0.95 ;
      RECT  1.15 0.95 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0258 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.875 1.105 ;
      RECT  0.75 1.105 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0258 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.545 0.7 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0258 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0201 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.615 0.495 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.42 1.41 1.54 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.85 0.05 1.02 0.195 ;
      RECT  0.345 0.05 0.465 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.075 0.185 0.25 0.69 ;
      RECT  0.075 0.69 0.175 1.11 ;
      RECT  0.075 1.11 0.25 1.515 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.555 0.285 1.32 0.39 ;
      RECT  1.41 0.185 1.53 0.485 ;
      RECT  0.355 0.485 1.53 0.575 ;
      RECT  0.355 0.575 0.445 0.775 ;
      RECT  0.285 0.775 0.445 0.945 ;
      RECT  0.355 0.945 0.445 1.435 ;
      RECT  0.355 1.435 1.32 1.525 ;
      RECT  1.125 1.525 1.32 1.56 ;
  END
END SEN_OA31_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OA31_1
#      Description : "One 3-input OR into 2-input AND"
#      Equation    : X=(A1|A2|A3)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA31_1
  CLASS CORE ;
  FOREIGN SEN_OA31_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.54 0.71 0.65 1.5 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.86 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.09 0.925 ;
      RECT  0.95 0.925 1.05 1.5 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0516 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.14 1.455 1.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.59 0.05 0.72 0.225 ;
      RECT  1.135 0.05 1.26 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.42 0.45 1.535 1.11 ;
      RECT  1.15 1.11 1.535 1.29 ;
      RECT  1.35 1.29 1.45 1.5 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.325 0.19 0.445 0.315 ;
      RECT  0.325 0.315 1.025 0.41 ;
      RECT  0.065 0.37 0.175 0.5 ;
      RECT  0.065 0.5 1.32 0.59 ;
      RECT  1.23 0.59 1.32 0.955 ;
      RECT  0.34 0.59 0.43 1.41 ;
  END
END SEN_OA31_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA31_2
#      Description : "One 3-input OR into 2-input AND"
#      Equation    : X=(A1|A2|A3)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA31_2
  CLASS CORE ;
  FOREIGN SEN_OA31_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.65 0.9 ;
      RECT  1.35 0.9 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 1.05 0.9 ;
      RECT  0.75 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.45 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1032 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.98 1.18 2.135 1.35 ;
      RECT  2.035 1.35 2.135 1.75 ;
      RECT  0.31 1.41 0.44 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  2.5 1.41 2.63 1.75 ;
      RECT  3.02 1.41 3.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.31 0.05 0.44 0.39 ;
      RECT  0.92 0.05 1.05 0.39 ;
      RECT  1.475 0.05 1.605 0.39 ;
      RECT  2.51 0.05 2.63 0.39 ;
      RECT  3.02 0.05 3.145 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.31 2.88 0.49 ;
      RECT  2.75 0.49 3.05 0.59 ;
      RECT  2.95 0.59 3.05 1.11 ;
      RECT  2.75 1.11 3.05 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.755 0.225 2.42 0.33 ;
      RECT  1.755 0.33 1.855 0.49 ;
      RECT  0.055 0.18 0.175 0.49 ;
      RECT  0.055 0.49 1.855 0.59 ;
      RECT  1.97 0.5 2.65 0.59 ;
      RECT  1.97 0.59 2.06 0.7 ;
      RECT  2.56 0.59 2.65 0.785 ;
      RECT  1.785 0.7 2.06 0.79 ;
      RECT  2.56 0.785 2.835 0.895 ;
      RECT  1.785 0.79 1.875 1.21 ;
      RECT  2.56 0.895 2.65 1.21 ;
      RECT  1.49 1.21 1.875 1.32 ;
      RECT  2.245 1.21 2.65 1.32 ;
      RECT  2.245 1.32 2.365 1.43 ;
      RECT  0.06 1.21 1.19 1.315 ;
      RECT  0.06 1.315 0.175 1.62 ;
      RECT  0.71 1.475 1.945 1.585 ;
  END
END SEN_OA31_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA31_4
#      Description : "One 3-input OR into 2-input AND"
#      Equation    : X=(A1|A2|A3)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA31_4
  CLASS CORE ;
  FOREIGN SEN_OA31_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 4.05 0.89 ;
      RECT  3.55 0.89 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2064 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.08 1.19 1.225 1.36 ;
      RECT  1.08 1.36 1.19 1.75 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  3.83 1.405 3.96 1.75 ;
      RECT  4.465 1.21 4.585 1.75 ;
      RECT  5.075 1.41 5.205 1.75 ;
      RECT  5.61 1.21 5.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      RECT  1.885 0.05 2.015 0.39 ;
      RECT  2.525 0.05 2.655 0.39 ;
      RECT  3.045 0.05 3.175 0.39 ;
      RECT  5.075 0.05 5.205 0.39 ;
      RECT  4.61 0.05 4.72 0.5 ;
      RECT  5.615 0.05 5.735 0.59 ;
      RECT  4.56 0.5 4.72 0.69 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.82 0.51 5.46 0.69 ;
      RECT  5.35 0.69 5.46 1.11 ;
      RECT  4.75 1.11 5.46 1.29 ;
    END
    ANTENNADIFFAREA 0.442 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.315 0.225 4.505 0.325 ;
      RECT  3.315 0.325 3.425 0.49 ;
      RECT  0.065 0.37 0.18 0.49 ;
      RECT  0.065 0.49 3.425 0.59 ;
      RECT  3.535 0.425 4.34 0.525 ;
      RECT  4.24 0.525 4.34 0.785 ;
      RECT  4.24 0.785 5.24 0.895 ;
      RECT  4.24 0.895 4.34 1.185 ;
      RECT  2.56 1.185 4.34 1.3 ;
      RECT  0.845 1.01 1.69 1.1 ;
      RECT  0.845 1.1 0.96 1.21 ;
      RECT  1.57 1.1 1.69 1.21 ;
      RECT  0.325 1.21 0.96 1.3 ;
      RECT  1.57 1.21 2.26 1.31 ;
      RECT  0.325 1.3 0.445 1.43 ;
      RECT  1.285 1.465 3.56 1.58 ;
  END
END SEN_OA31_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA31_8
#      Description : "One 3-input OR into 2-input AND"
#      Equation    : X=(A1|A2|A3)&B
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA31_8
  CLASS CORE ;
  FOREIGN SEN_OA31_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.91 0.71 6.65 0.91 ;
      RECT  6.55 0.91 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3402 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.315 0.695 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3402 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.51 3.45 0.71 ;
      RECT  2.55 0.71 3.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3402 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 8.25 0.915 ;
      RECT  8.15 0.915 8.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2634 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  0.59 1.4 0.71 1.75 ;
      RECT  1.11 1.4 1.23 1.75 ;
      RECT  1.63 1.4 1.75 1.75 ;
      RECT  2.15 1.23 2.27 1.75 ;
      RECT  2.68 1.495 2.855 1.75 ;
      RECT  3.205 1.495 3.38 1.75 ;
      RECT  3.725 1.495 3.9 1.75 ;
      RECT  7.12 1.45 7.24 1.75 ;
      RECT  7.64 1.455 7.76 1.75 ;
      RECT  8.18 1.21 8.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  2.655 0.05 2.825 0.195 ;
      RECT  3.195 0.05 3.365 0.195 ;
      RECT  4.465 0.05 4.585 0.27 ;
      RECT  3.925 0.05 4.045 0.275 ;
      RECT  5.01 0.05 5.13 0.31 ;
      RECT  0.565 0.05 0.735 0.32 ;
      RECT  1.085 0.05 1.255 0.32 ;
      RECT  1.605 0.05 1.775 0.32 ;
      RECT  5.55 0.05 5.67 0.36 ;
      RECT  6.08 0.05 6.2 0.36 ;
      RECT  6.6 0.05 6.72 0.36 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  2.15 0.05 2.27 0.6 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.28 0.415 2.06 0.535 ;
      RECT  0.55 0.535 2.06 0.545 ;
      RECT  0.55 0.545 0.85 1.11 ;
      RECT  0.31 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.855 0.21 8.07 0.34 ;
      RECT  6.855 0.34 6.985 0.45 ;
      RECT  2.36 0.285 3.775 0.415 ;
      RECT  3.66 0.415 3.775 0.45 ;
      RECT  3.66 0.45 6.985 0.58 ;
      RECT  4.195 0.265 4.315 0.45 ;
      RECT  8.16 0.32 8.28 0.475 ;
      RECT  7.125 0.475 8.28 0.595 ;
      RECT  7.125 0.595 7.255 1.23 ;
      RECT  0.98 0.785 2.285 0.895 ;
      RECT  2.155 0.895 2.285 1.0 ;
      RECT  2.155 1.0 5.445 1.13 ;
      RECT  5.315 1.13 5.445 1.23 ;
      RECT  5.315 1.23 8.07 1.36 ;
      RECT  2.4 1.25 5.22 1.4 ;
      RECT  4.195 1.49 7.03 1.66 ;
  END
END SEN_OA31_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OA32_1
#      Description : "One 3-input OR + one 2-input OR into 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA32_1
  CLASS CORE ;
  FOREIGN SEN_OA32_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.11 ;
      RECT  0.55 1.11 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0618 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.2 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.455 1.58 1.625 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.88 0.05 1.05 0.19 ;
      RECT  1.5 0.05 1.63 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.3 1.93 0.5 ;
      RECT  1.835 0.5 1.93 1.11 ;
      RECT  1.75 1.11 1.93 1.49 ;
    END
    ANTENNADIFFAREA 0.184 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.225 0.18 1.345 0.295 ;
      RECT  0.07 0.295 1.345 0.4 ;
      RECT  0.07 0.4 0.18 0.52 ;
      RECT  0.29 0.49 1.64 0.59 ;
      RECT  1.55 0.59 1.64 0.755 ;
      RECT  1.55 0.755 1.745 0.925 ;
      RECT  1.55 0.925 1.64 1.4 ;
      RECT  0.6 1.4 1.64 1.49 ;
      RECT  0.6 1.49 0.72 1.62 ;
  END
END SEN_OA32_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA32_2
#      Description : "One 3-input OR + one 2-input OR into 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA32_2
  CLASS CORE ;
  FOREIGN SEN_OA32_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.825 0.89 ;
      RECT  0.55 0.89 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1236 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.41 0.44 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  2.555 1.41 2.675 1.75 ;
      RECT  3.065 1.41 3.195 1.75 ;
      RECT  3.59 1.21 3.71 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  1.35 0.05 1.48 0.39 ;
      RECT  1.795 0.05 1.925 0.39 ;
      RECT  2.33 0.05 2.46 0.39 ;
      RECT  3.065 0.05 3.195 0.39 ;
      RECT  3.59 0.05 3.71 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.345 0.3 3.46 1.3 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.55 0.25 2.97 0.35 ;
      RECT  2.55 0.35 2.64 0.495 ;
      RECT  0.055 0.195 1.21 0.31 ;
      RECT  0.055 0.31 0.175 0.39 ;
      RECT  1.105 0.31 1.21 0.495 ;
      RECT  1.105 0.495 2.64 0.595 ;
      RECT  0.27 0.45 1.015 0.55 ;
      RECT  0.915 0.55 1.015 1.205 ;
      RECT  0.81 1.205 1.015 1.305 ;
      RECT  3.15 0.72 3.25 1.15 ;
      RECT  3.045 1.15 3.25 1.25 ;
      RECT  1.535 1.145 1.715 1.245 ;
      RECT  1.535 1.245 1.9 1.335 ;
      RECT  2.035 1.18 2.955 1.28 ;
      RECT  0.055 1.21 0.69 1.3 ;
      RECT  0.58 1.3 0.69 1.42 ;
      RECT  0.055 1.3 0.175 1.62 ;
      RECT  0.58 1.42 1.215 1.51 ;
      RECT  1.095 1.51 1.215 1.63 ;
      RECT  1.23 1.225 1.425 1.325 ;
      RECT  1.335 1.325 1.425 1.455 ;
      RECT  1.335 1.455 2.465 1.555 ;
      LAYER M2 ;
      RECT  0.83 1.15 3.225 1.25 ;
      LAYER V1 ;
      RECT  0.915 1.15 1.015 1.25 ;
      RECT  1.575 1.15 1.675 1.25 ;
      RECT  3.085 1.15 3.185 1.25 ;
  END
END SEN_OA32_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA32_4
#      Description : "One 3-input OR + one 2-input OR into 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA32_4
  CLASS CORE ;
  FOREIGN SEN_OA32_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 4.25 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.31 5.65 0.71 ;
      RECT  4.95 0.71 5.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2472 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  4.735 1.41 4.86 1.75 ;
      RECT  5.25 1.41 5.38 1.75 ;
      RECT  5.775 1.21 5.895 1.75 ;
      RECT  6.29 1.41 6.42 1.75 ;
      RECT  6.815 1.21 6.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  6.295 0.05 6.415 0.365 ;
      RECT  2.4 0.05 2.53 0.39 ;
      RECT  2.92 0.05 3.05 0.39 ;
      RECT  3.435 0.05 3.565 0.39 ;
      RECT  3.96 0.05 4.09 0.39 ;
      RECT  4.485 0.05 4.615 0.39 ;
      RECT  5.005 0.05 5.135 0.39 ;
      RECT  5.745 0.05 5.875 0.39 ;
      RECT  6.815 0.05 6.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.51 6.665 0.69 ;
      RECT  6.55 0.69 6.665 1.11 ;
      RECT  6.035 1.11 6.665 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.23 2.26 0.345 ;
      RECT  0.065 0.345 0.185 0.45 ;
      RECT  2.15 0.345 2.26 0.48 ;
      RECT  2.15 0.48 5.415 0.58 ;
      RECT  5.81 0.79 6.44 0.895 ;
      RECT  5.81 0.895 5.9 1.01 ;
      RECT  3.54 1.01 5.9 1.1 ;
      RECT  3.54 1.1 3.63 1.21 ;
      RECT  0.28 0.485 2.03 0.59 ;
      RECT  1.94 0.59 2.03 1.21 ;
      RECT  1.335 1.21 3.63 1.31 ;
      RECT  3.72 1.19 5.665 1.29 ;
      RECT  3.72 1.29 3.82 1.385 ;
      RECT  0.07 1.21 1.225 1.32 ;
      RECT  0.07 1.32 0.185 1.43 ;
      RECT  1.1 1.32 1.225 1.49 ;
      RECT  1.1 1.49 2.265 1.63 ;
      RECT  2.145 1.42 2.265 1.49 ;
      RECT  2.37 1.475 4.645 1.575 ;
  END
END SEN_OA32_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OA33_0P5
#      Description : "Two 3-input ORs into a 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA33_0P5
  CLASS CORE ;
  FOREIGN SEN_OA33_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0213 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.34 0.71 1.45 1.66 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0213 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0213 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0213 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0213 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0213 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.085 1.41 0.225 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.74 1.215 1.845 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  1.165 0.05 1.335 0.215 ;
      RECT  1.725 0.05 1.845 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.145 2.09 0.43 ;
      RECT  1.95 0.43 2.05 1.31 ;
      RECT  1.95 1.31 2.105 1.51 ;
    END
    ANTENNADIFFAREA 0.086 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.38 0.14 1.04 0.23 ;
      RECT  0.92 0.23 1.04 0.305 ;
      RECT  0.38 0.23 0.5 0.38 ;
      RECT  0.92 0.305 1.58 0.395 ;
      RECT  1.46 0.18 1.58 0.305 ;
      RECT  0.12 0.15 0.24 0.47 ;
      RECT  0.12 0.47 0.77 0.485 ;
      RECT  0.65 0.32 0.77 0.47 ;
      RECT  0.12 0.485 1.845 0.56 ;
      RECT  0.37 0.56 1.845 0.575 ;
      RECT  1.755 0.575 1.845 0.96 ;
      RECT  0.37 0.575 0.46 1.415 ;
      RECT  0.37 1.415 1.08 1.53 ;
  END
END SEN_OA33_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OA33_1
#      Description : "Two 3-input ORs into a 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA33_1
  CLASS CORE ;
  FOREIGN SEN_OA33_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.17 0.885 ;
      RECT  0.95 0.885 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.32 0.71 1.45 1.11 ;
      RECT  1.15 1.11 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0369 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.09 1.41 0.23 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.74 1.205 1.845 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  1.165 0.05 1.335 0.215 ;
      RECT  1.725 0.05 1.845 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.285 2.105 0.485 ;
      RECT  1.95 0.485 2.05 1.315 ;
      RECT  1.95 1.315 2.105 1.51 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.38 0.14 1.04 0.23 ;
      RECT  0.92 0.23 1.04 0.305 ;
      RECT  0.38 0.23 0.5 0.38 ;
      RECT  0.92 0.305 1.58 0.395 ;
      RECT  1.46 0.185 1.58 0.305 ;
      RECT  0.12 0.24 0.24 0.47 ;
      RECT  0.12 0.47 0.77 0.485 ;
      RECT  0.65 0.32 0.77 0.47 ;
      RECT  0.12 0.485 1.86 0.56 ;
      RECT  0.37 0.56 1.86 0.575 ;
      RECT  1.77 0.575 1.86 0.94 ;
      RECT  0.37 0.575 0.46 1.425 ;
      RECT  0.37 1.425 1.09 1.545 ;
  END
END SEN_OA33_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OA33_1P5
#      Description : "Two 3-input ORs into a 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA33_1P5
  CLASS CORE ;
  FOREIGN SEN_OA33_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.11 0.885 ;
      RECT  0.95 0.885 1.25 0.985 ;
      RECT  1.15 0.985 1.25 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.26 0.675 1.45 0.79 ;
      RECT  1.35 0.79 1.45 1.49 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.665 1.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.665 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.64 1.41 1.78 1.75 ;
      RECT  2.18 1.41 2.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  1.095 0.05 1.265 0.215 ;
      RECT  2.18 0.05 2.32 0.39 ;
      RECT  1.65 0.05 1.77 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.92 0.245 2.05 0.5 ;
      RECT  1.92 0.5 2.25 0.59 ;
      RECT  2.15 0.59 2.25 1.215 ;
      RECT  1.91 1.215 2.25 1.31 ;
      RECT  1.91 1.31 2.05 1.49 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.39 0.185 1.51 0.305 ;
      RECT  0.28 0.305 1.51 0.395 ;
      RECT  0.07 0.33 0.19 0.485 ;
      RECT  0.07 0.485 1.83 0.575 ;
      RECT  0.07 0.575 0.43 0.58 ;
      RECT  1.74 0.575 1.83 0.81 ;
      RECT  0.34 0.58 0.43 1.435 ;
      RECT  1.74 0.81 2.04 0.92 ;
      RECT  0.34 1.435 1.015 1.555 ;
  END
END SEN_OA33_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OA33_2
#      Description : "Two 3-input ORs into a 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA33_2
  CLASS CORE ;
  FOREIGN SEN_OA33_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.615 1.855 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.145 0.615 2.25 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 0.63 ;
      RECT  2.54 0.63 2.85 0.74 ;
      RECT  2.54 0.74 2.65 1.125 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.45 1.25 0.935 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.66 0.65 0.9 ;
      RECT  0.55 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0696 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.44 0.53 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  2.345 1.585 2.515 1.75 ;
      RECT  2.87 1.43 2.99 1.75 ;
      RECT  3.41 1.21 3.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  1.605 0.05 1.775 0.345 ;
      RECT  2.145 0.05 2.315 0.345 ;
      RECT  2.75 0.05 2.89 0.39 ;
      RECT  3.41 0.05 3.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.14 0.27 3.25 1.505 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.125 0.14 1.47 0.23 ;
      RECT  0.125 0.23 0.24 0.39 ;
      RECT  0.645 0.23 0.765 0.39 ;
      RECT  1.35 0.23 1.47 0.435 ;
      RECT  1.35 0.435 2.55 0.525 ;
      RECT  1.9 0.21 2.03 0.435 ;
      RECT  2.43 0.21 2.55 0.435 ;
      RECT  0.4 0.335 0.49 0.48 ;
      RECT  0.4 0.48 1.05 0.57 ;
      RECT  0.88 0.325 1.05 0.48 ;
      RECT  0.955 0.57 1.05 1.035 ;
      RECT  0.955 1.035 1.63 1.125 ;
      RECT  1.54 1.125 1.63 1.225 ;
      RECT  1.54 1.225 3.04 1.315 ;
      RECT  2.95 0.755 3.04 1.225 ;
      RECT  0.125 1.255 1.355 1.345 ;
      RECT  0.125 1.345 0.245 1.49 ;
      RECT  2.1 1.405 2.76 1.495 ;
      RECT  2.64 1.495 2.76 1.625 ;
      RECT  2.1 1.495 2.22 1.63 ;
      RECT  0.855 1.435 1.49 1.54 ;
      RECT  1.37 1.54 1.49 1.635 ;
  END
END SEN_OA33_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OA33_3
#      Description : "Two 3-input ORs into a 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA33_3
  CLASS CORE ;
  FOREIGN SEN_OA33_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.895 ;
      RECT  1.55 0.895 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.895 ;
      RECT  0.75 0.895 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.895 ;
      RECT  0.15 0.895 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.65 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.05 0.895 ;
      RECT  2.95 0.895 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1026 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.415 0.435 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  3.375 1.415 3.495 1.75 ;
      RECT  4.08 1.2 4.2 1.75 ;
      RECT  4.6 1.21 4.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.315 0.05 0.435 0.38 ;
      RECT  0.835 0.05 0.955 0.38 ;
      RECT  1.585 0.05 1.705 0.38 ;
      RECT  4.34 0.05 4.46 0.39 ;
      RECT  3.88 0.05 3.985 0.545 ;
      RECT  3.795 0.545 3.985 0.665 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.095 0.28 4.25 0.51 ;
      RECT  4.095 0.51 4.72 0.69 ;
      RECT  4.35 0.69 4.45 0.99 ;
      RECT  3.82 0.99 4.45 1.08 ;
      RECT  3.82 1.08 3.925 1.16 ;
      RECT  4.35 1.08 4.45 1.51 ;
    END
    ANTENNADIFFAREA 0.369 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.85 0.19 3.755 0.305 ;
      RECT  3.635 0.305 3.755 0.36 ;
      RECT  1.85 0.305 1.96 0.475 ;
      RECT  0.055 0.16 0.175 0.475 ;
      RECT  0.055 0.475 1.96 0.575 ;
      RECT  0.575 0.355 0.695 0.475 ;
      RECT  1.21 0.355 1.33 0.475 ;
      RECT  2.08 0.455 3.68 0.56 ;
      RECT  3.59 0.56 3.68 0.785 ;
      RECT  2.08 0.56 2.17 1.22 ;
      RECT  3.59 0.785 4.26 0.895 ;
      RECT  1.325 1.22 2.17 1.23 ;
      RECT  1.325 1.23 2.485 1.325 ;
      RECT  1.325 1.325 1.445 1.42 ;
      RECT  2.365 1.325 2.485 1.425 ;
      RECT  0.055 1.215 1.215 1.325 ;
      RECT  1.095 1.325 1.215 1.42 ;
      RECT  0.055 1.325 0.175 1.635 ;
      RECT  2.595 1.22 3.75 1.325 ;
      RECT  2.595 1.325 2.715 1.425 ;
      RECT  3.635 1.325 3.75 1.635 ;
      RECT  0.835 1.415 0.955 1.55 ;
      RECT  0.835 1.55 1.705 1.64 ;
      RECT  1.585 1.415 1.705 1.55 ;
      RECT  2.105 1.415 2.225 1.55 ;
      RECT  2.105 1.55 2.975 1.64 ;
      RECT  2.855 1.415 2.975 1.55 ;
  END
END SEN_OA33_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OA33_4
#      Description : "Two 3-input ORs into a 2-input AND"
#      Equation    : X=(A1|A2|A3)&(B1|B2|B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OA33_4
  CLASS CORE ;
  FOREIGN SEN_OA33_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.895 ;
      RECT  1.55 0.895 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.895 ;
      RECT  0.75 0.895 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.895 ;
      RECT  0.15 0.895 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END A3
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.65 0.89 ;
      RECT  2.35 0.89 2.45 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.05 0.895 ;
      RECT  2.95 0.895 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.129 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.44 0.435 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  3.33 1.41 3.455 1.75 ;
      RECT  4.035 1.4 4.155 1.75 ;
      RECT  4.555 1.4 4.675 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  4.295 0.05 4.415 0.36 ;
      RECT  0.315 0.05 0.435 0.38 ;
      RECT  0.835 0.05 0.955 0.38 ;
      RECT  1.585 0.05 1.705 0.38 ;
      RECT  3.835 0.05 3.935 0.545 ;
      RECT  4.815 0.05 4.935 0.59 ;
      RECT  3.725 0.545 3.935 0.665 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.035 0.375 4.155 0.465 ;
      RECT  4.035 0.465 4.7 0.585 ;
      RECT  4.55 0.585 4.65 1.11 ;
      RECT  3.79 0.99 3.895 1.11 ;
      RECT  3.79 1.11 4.935 1.29 ;
    END
    ANTENNADIFFAREA 0.484 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.85 0.19 3.71 0.32 ;
      RECT  3.59 0.32 3.71 0.36 ;
      RECT  1.85 0.32 1.96 0.475 ;
      RECT  0.055 0.16 0.175 0.475 ;
      RECT  0.055 0.475 1.96 0.575 ;
      RECT  2.08 0.455 3.635 0.56 ;
      RECT  3.545 0.56 3.635 0.785 ;
      RECT  2.08 0.56 2.17 1.22 ;
      RECT  3.545 0.785 4.45 0.895 ;
      RECT  1.325 1.22 2.17 1.23 ;
      RECT  1.325 1.23 2.475 1.325 ;
      RECT  1.325 1.325 1.44 1.425 ;
      RECT  2.365 1.325 2.475 1.45 ;
      RECT  2.565 0.99 2.67 1.18 ;
      RECT  2.565 1.18 3.7 1.28 ;
      RECT  3.59 1.28 3.7 1.635 ;
      RECT  0.055 1.215 1.215 1.325 ;
      RECT  1.095 1.325 1.215 1.425 ;
      RECT  0.055 1.325 0.175 1.63 ;
      RECT  0.835 1.415 0.955 1.55 ;
      RECT  0.835 1.55 1.705 1.64 ;
      RECT  1.585 1.415 1.705 1.55 ;
      RECT  2.105 1.415 2.225 1.55 ;
      RECT  2.105 1.55 2.93 1.64 ;
      RECT  2.81 1.415 2.93 1.55 ;
  END
END SEN_OA33_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI2111_0P5
#      Description : "One 2-input OR into 4-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI2111_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI2111_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0282 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0282 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0258 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0258 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.745 0.465 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0258 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.85 1.41 0.97 1.75 ;
      RECT  1.38 1.41 1.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.33 0.05 0.45 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.14 0.24 1.54 0.36 ;
      RECT  1.14 0.36 1.25 1.23 ;
      RECT  0.55 1.23 1.25 1.32 ;
      RECT  0.55 1.32 0.71 1.61 ;
      RECT  1.125 1.32 1.25 1.61 ;
    END
    ANTENNADIFFAREA 0.118 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.54 0.23 0.76 0.35 ;
      RECT  0.54 0.35 0.63 0.475 ;
      RECT  0.07 0.2 0.19 0.475 ;
      RECT  0.07 0.475 0.63 0.565 ;
  END
END SEN_OAI2111_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI2111_1
#      Description : "One 2-input OR into 4-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI2111_1
  CLASS CORE ;
  FOREIGN SEN_OAI2111_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.58 0.9 ;
      RECT  0.35 0.9 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.31 1.05 0.955 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 0.75 ;
      RECT  0.705 0.75 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.855 1.41 0.985 1.75 ;
      RECT  1.385 1.41 1.515 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.325 0.05 0.455 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.145 0.31 1.51 0.49 ;
      RECT  1.145 0.49 1.25 1.21 ;
      RECT  0.54 1.21 1.25 1.32 ;
    END
    ANTENNADIFFAREA 0.317 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.55 0.24 0.77 0.36 ;
      RECT  0.55 0.36 0.65 0.48 ;
      RECT  0.07 0.37 0.19 0.48 ;
      RECT  0.07 0.48 0.65 0.59 ;
  END
END SEN_OAI2111_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI2111_2
#      Description : "One 2-input OR into 4-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI2111_2
  CLASS CORE ;
  FOREIGN SEN_OAI2111_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.5 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.355 1.42 1.48 1.75 ;
      RECT  1.87 1.42 2.0 1.75 ;
      RECT  2.435 1.42 2.565 1.75 ;
      RECT  3.0 1.21 3.12 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  0.84 0.05 0.97 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.495 2.85 1.21 ;
      RECT  0.82 1.21 2.85 1.33 ;
    END
    ANTENNADIFFAREA 0.576 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.875 0.18 1.995 0.26 ;
      RECT  1.875 0.26 3.12 0.38 ;
      RECT  3.0 0.18 3.12 0.26 ;
      RECT  1.105 0.225 1.77 0.35 ;
      RECT  1.105 0.35 1.225 0.47 ;
      RECT  0.065 0.37 0.185 0.47 ;
      RECT  0.065 0.47 1.225 0.59 ;
      RECT  1.32 0.47 2.31 0.59 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.585 1.3 0.705 1.44 ;
      RECT  0.585 1.44 1.265 1.56 ;
  END
END SEN_OAI2111_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI2111_4
#      Description : "One 2-input OR into 4-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2&B3)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI2111_4
  CLASS CORE ;
  FOREIGN SEN_OAI2111_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.25 0.89 ;
      RECT  4.75 0.89 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.425 0.45 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.84 1.425 0.97 1.75 ;
      RECT  2.395 1.42 2.52 1.75 ;
      RECT  2.91 1.42 3.04 1.75 ;
      RECT  3.44 1.42 3.57 1.75 ;
      RECT  3.97 1.42 4.1 1.75 ;
      RECT  4.49 1.42 4.62 1.75 ;
      RECT  5.04 1.42 5.17 1.75 ;
      RECT  5.6 1.21 5.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  0.84 0.05 0.97 0.38 ;
      RECT  1.36 0.05 1.49 0.38 ;
      RECT  1.88 0.05 2.01 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.7 0.47 5.45 0.59 ;
      RECT  5.35 0.59 5.45 1.21 ;
      RECT  1.315 1.21 5.45 1.33 ;
    END
    ANTENNADIFFAREA 1.152 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.145 0.225 3.33 0.35 ;
      RECT  2.145 0.35 2.265 0.47 ;
      RECT  0.065 0.37 0.185 0.47 ;
      RECT  0.065 0.47 2.265 0.59 ;
      RECT  3.43 0.26 5.72 0.38 ;
      RECT  5.6 0.38 5.72 0.48 ;
      RECT  2.365 0.47 4.41 0.59 ;
      RECT  0.065 1.21 1.225 1.33 ;
      RECT  0.065 1.33 0.185 1.43 ;
      RECT  1.105 1.33 1.225 1.44 ;
      RECT  1.105 1.44 2.305 1.56 ;
  END
END SEN_OAI2111_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI211_0P5
#      Description : "One 2-input OR into 3-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI211_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI211_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.5 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.885 1.58 1.015 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.31 0.05 0.48 0.21 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.24 1.315 0.36 ;
      RECT  0.95 0.36 1.05 1.31 ;
      RECT  0.55 1.31 1.275 1.49 ;
    END
    ANTENNADIFFAREA 0.145 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.2 0.185 0.3 ;
      RECT  0.065 0.3 0.78 0.42 ;
  END
END SEN_OAI211_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI211_1
#      Description : "One 2-input OR into 3-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI211_1
  CLASS CORE ;
  FOREIGN SEN_OAI211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.5 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.615 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  0.885 1.45 1.015 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.31 0.05 0.48 0.32 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.24 1.315 0.36 ;
      RECT  0.95 0.36 1.05 1.24 ;
      RECT  0.56 1.24 1.325 1.36 ;
    END
    ANTENNADIFFAREA 0.29 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.3 0.185 0.41 ;
      RECT  0.065 0.41 0.78 0.52 ;
  END
END SEN_OAI211_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI211_2
#      Description : "One 2-input OR into 3-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI211_2
  CLASS CORE ;
  FOREIGN SEN_OAI211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.625 1.42 1.755 1.75 ;
      RECT  2.145 1.42 2.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.58 0.05 0.71 0.38 ;
      RECT  1.1 0.05 1.23 0.38 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.44 2.32 0.565 ;
      RECT  1.95 0.565 2.05 1.21 ;
      RECT  0.815 1.21 2.53 1.33 ;
      RECT  2.41 1.33 2.53 1.43 ;
    END
    ANTENNADIFFAREA 0.522 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.32 0.215 2.53 0.335 ;
      RECT  2.41 0.335 2.53 0.44 ;
      RECT  0.285 0.47 1.8 0.59 ;
      RECT  0.065 1.21 0.705 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  0.585 1.32 0.705 1.44 ;
      RECT  0.585 1.44 1.28 1.56 ;
  END
END SEN_OAI211_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI211_3
#      Description : "One 2-input OR into 3-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI211_3
  CLASS CORE ;
  FOREIGN SEN_OAI211_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.74 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.58 1.42 0.71 1.75 ;
      RECT  1.88 1.44 2.01 1.75 ;
      RECT  2.4 1.44 2.53 1.75 ;
      RECT  2.93 1.44 3.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  0.84 0.05 0.97 0.38 ;
      RECT  1.36 0.05 1.49 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.2 0.37 3.32 0.47 ;
      RECT  2.55 0.47 3.32 0.59 ;
      RECT  2.55 0.59 2.65 1.23 ;
      RECT  1.08 1.23 3.305 1.35 ;
      RECT  3.15 1.35 3.305 1.49 ;
    END
    ANTENNADIFFAREA 0.748 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.83 0.24 3.1 0.36 ;
      RECT  0.065 0.37 0.185 0.47 ;
      RECT  0.065 0.47 2.32 0.59 ;
      RECT  0.28 1.21 0.965 1.33 ;
      RECT  0.845 1.33 0.965 1.44 ;
      RECT  0.845 1.44 1.54 1.56 ;
  END
END SEN_OAI211_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI211_4
#      Description : "One 2-input OR into 3-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI211_4
  CLASS CORE ;
  FOREIGN SEN_OAI211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  2.585 1.42 2.715 1.75 ;
      RECT  3.105 1.42 3.235 1.75 ;
      RECT  3.625 1.42 3.755 1.75 ;
      RECT  4.145 1.42 4.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.58 0.05 0.71 0.38 ;
      RECT  1.1 0.05 1.23 0.38 ;
      RECT  1.62 0.05 1.75 0.38 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  2.145 0.05 2.25 0.68 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.44 4.32 0.565 ;
      RECT  3.55 0.565 3.65 1.21 ;
      RECT  1.315 1.21 4.53 1.33 ;
      RECT  4.41 1.33 4.53 1.43 ;
    END
    ANTENNADIFFAREA 0.955 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.34 0.215 4.53 0.335 ;
      RECT  2.34 0.335 2.45 0.385 ;
      RECT  4.41 0.335 4.53 0.44 ;
      RECT  2.375 0.475 3.28 0.595 ;
      RECT  2.375 0.595 2.465 0.77 ;
      RECT  0.285 0.47 2.03 0.59 ;
      RECT  1.94 0.59 2.03 0.77 ;
      RECT  1.94 0.77 2.465 0.86 ;
      RECT  0.065 1.205 1.225 1.325 ;
      RECT  0.065 1.325 0.185 1.43 ;
      RECT  1.105 1.325 1.225 1.45 ;
      RECT  1.105 1.45 2.32 1.57 ;
  END
END SEN_OAI211_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI211_8
#      Description : "One 2-input OR into 3-input NAND"
#      Equation    : X=!((A1|A2)&B1&B2)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI211_8
  CLASS CORE ;
  FOREIGN SEN_OAI211_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 6.25 0.89 ;
      RECT  4.95 0.89 5.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 8.45 0.89 ;
      RECT  8.35 0.89 8.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.665 0.91 ;
      RECT  0.15 0.91 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 4.25 0.91 ;
      RECT  4.15 0.91 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4992 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.59 1.41 0.71 1.75 ;
      RECT  1.11 1.41 1.23 1.75 ;
      RECT  1.63 1.41 1.75 1.75 ;
      RECT  2.15 1.41 2.27 1.75 ;
      RECT  2.67 1.41 2.79 1.75 ;
      RECT  3.19 1.41 3.31 1.75 ;
      RECT  3.685 1.48 3.855 1.75 ;
      RECT  4.205 1.48 4.375 1.75 ;
      RECT  6.78 1.41 6.9 1.75 ;
      RECT  7.3 1.41 7.425 1.75 ;
      RECT  7.815 1.41 7.94 1.75 ;
      RECT  8.34 1.41 8.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  4.7 0.05 4.82 0.35 ;
      RECT  5.22 0.05 5.34 0.35 ;
      RECT  5.74 0.05 5.86 0.35 ;
      RECT  6.26 0.05 6.38 0.35 ;
      RECT  6.78 0.05 6.9 0.35 ;
      RECT  7.3 0.05 7.42 0.35 ;
      RECT  7.82 0.05 7.94 0.35 ;
      RECT  8.34 0.05 8.46 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.28 0.44 2.05 0.565 ;
      RECT  1.345 0.565 2.05 0.61 ;
      RECT  1.88 0.61 2.05 1.11 ;
      RECT  0.34 1.11 4.05 1.22 ;
      RECT  0.34 1.22 4.635 1.29 ;
      RECT  3.855 1.29 4.635 1.39 ;
      RECT  4.465 1.39 4.635 1.41 ;
      RECT  4.465 1.41 4.825 1.47 ;
      RECT  4.465 1.47 6.435 1.59 ;
    END
    ANTENNADIFFAREA 1.76 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.605 0.18 2.79 0.23 ;
      RECT  0.07 0.23 4.405 0.35 ;
      RECT  0.07 0.35 0.19 0.45 ;
      RECT  8.6 0.34 8.72 0.44 ;
      RECT  3.945 0.44 8.72 0.49 ;
      RECT  2.36 0.49 8.72 0.56 ;
      RECT  2.36 0.56 7.185 0.61 ;
      RECT  4.395 1.015 4.815 1.13 ;
      RECT  4.725 1.13 4.815 1.18 ;
      RECT  4.725 1.18 8.72 1.29 ;
      RECT  5.98 1.11 7.16 1.18 ;
      RECT  8.6 1.29 8.72 1.41 ;
  END
END SEN_OAI211_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_0P5
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI21_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.69 0.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0321 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.675 1.43 0.795 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.39 0.05 0.51 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.22 1.06 1.22 ;
      RECT  0.35 1.22 1.06 1.31 ;
      RECT  0.35 1.31 0.45 1.44 ;
      RECT  0.94 1.31 1.06 1.52 ;
      RECT  0.08 1.44 0.45 1.56 ;
    END
    ANTENNADIFFAREA 0.134 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.11 0.21 0.23 0.44 ;
      RECT  0.11 0.44 0.79 0.56 ;
      RECT  0.67 0.21 0.79 0.44 ;
  END
END SEN_OAI21_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_1
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_1
  CLASS CORE ;
  FOREIGN SEN_OAI21_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.69 0.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.675 1.43 0.795 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.39 0.05 0.51 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.31 1.06 1.22 ;
      RECT  0.35 1.22 1.06 1.31 ;
      RECT  0.35 1.31 0.45 1.44 ;
      RECT  0.94 1.31 1.06 1.49 ;
      RECT  0.08 1.44 0.45 1.56 ;
    END
    ANTENNADIFFAREA 0.267 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.08 0.44 0.83 0.56 ;
  END
END SEN_OAI21_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_2
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_2
  CLASS CORE ;
  FOREIGN SEN_OAI21_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 0.695 ;
      RECT  1.55 0.695 1.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.41 0.445 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.565 1.25 1.685 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.325 0.05 0.445 0.35 ;
      RECT  0.845 0.05 0.965 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.45 1.59 0.56 ;
      RECT  1.35 0.56 1.45 1.03 ;
      RECT  1.15 1.03 1.945 1.15 ;
      RECT  1.825 1.15 1.945 1.23 ;
      RECT  1.15 1.15 1.25 1.24 ;
      RECT  0.82 1.24 1.25 1.35 ;
    END
    ANTENNADIFFAREA 0.369 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.13 0.24 1.85 0.36 ;
      RECT  1.13 0.36 1.25 0.44 ;
      RECT  0.065 0.34 0.185 0.44 ;
      RECT  0.065 0.44 1.25 0.56 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.19 1.43 ;
      RECT  0.585 1.3 0.705 1.44 ;
      RECT  0.585 1.44 1.28 1.56 ;
  END
END SEN_OAI21_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_3
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_3
  CLASS CORE ;
  FOREIGN SEN_OAI21_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.14 0.71 2.45 0.915 ;
      RECT  2.35 0.915 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  0.59 1.45 0.71 1.75 ;
      RECT  1.89 1.41 2.01 1.75 ;
      RECT  2.41 1.41 2.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.33 0.05 0.45 0.35 ;
      RECT  0.85 0.05 0.97 0.35 ;
      RECT  1.37 0.05 1.49 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.41 0.34 2.53 0.445 ;
      RECT  1.85 0.445 2.53 0.56 ;
      RECT  1.95 0.56 2.05 1.11 ;
      RECT  1.63 1.11 2.26 1.29 ;
      RECT  1.63 1.29 1.76 1.45 ;
      RECT  1.06 1.45 1.76 1.56 ;
    END
    ANTENNADIFFAREA 0.529 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.63 0.22 2.32 0.335 ;
      RECT  1.63 0.335 1.75 0.44 ;
      RECT  0.07 0.34 0.19 0.44 ;
      RECT  0.07 0.44 1.75 0.56 ;
      RECT  0.305 1.24 1.515 1.36 ;
  END
END SEN_OAI21_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_4
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_4
  CLASS CORE ;
  FOREIGN SEN_OAI21_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.85 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.45 0.435 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.835 1.45 0.955 1.75 ;
      RECT  2.385 1.41 2.505 1.75 ;
      RECT  2.905 1.41 3.025 1.75 ;
      RECT  3.425 1.41 3.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.575 0.05 0.695 0.35 ;
      RECT  1.095 0.05 1.215 0.35 ;
      RECT  1.615 0.05 1.735 0.35 ;
      RECT  2.135 0.05 2.255 0.36 ;
      RECT  0.055 0.05 0.175 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.62 0.5 3.34 0.62 ;
      RECT  2.75 0.62 2.85 1.11 ;
      RECT  1.35 1.11 3.25 1.2 ;
      RECT  1.35 1.2 3.31 1.29 ;
    END
    ANTENNADIFFAREA 0.668 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.425 0.17 3.545 0.27 ;
      RECT  2.39 0.27 3.545 0.39 ;
      RECT  2.39 0.39 2.505 0.45 ;
      RECT  0.27 0.45 2.505 0.56 ;
      RECT  0.055 1.24 1.215 1.36 ;
      RECT  1.095 1.36 1.215 1.44 ;
      RECT  0.055 1.36 0.175 1.63 ;
      RECT  1.095 1.44 2.28 1.56 ;
  END
END SEN_OAI21_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_16
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_16
  CLASS CORE ;
  FOREIGN SEN_OAI21_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.55 0.71 7.865 0.93 ;
      RECT  6.77 0.71 7.07 0.9 ;
      RECT  5.825 0.71 6.125 0.9 ;
      RECT  4.785 0.71 5.085 0.9 ;
      RECT  3.755 0.71 4.055 0.9 ;
      RECT  2.695 0.71 3.035 0.9 ;
      RECT  1.675 0.71 1.975 0.89 ;
      RECT  0.615 0.71 1.02 0.9 ;
      LAYER M2 ;
      RECT  0.615 0.75 7.89 0.85 ;
      LAYER V1 ;
      RECT  7.55 0.75 7.65 0.85 ;
      RECT  7.75 0.75 7.85 0.85 ;
      RECT  6.77 0.75 6.87 0.85 ;
      RECT  6.97 0.75 7.07 0.85 ;
      RECT  5.825 0.75 5.925 0.85 ;
      RECT  6.025 0.75 6.125 0.85 ;
      RECT  4.785 0.75 4.885 0.85 ;
      RECT  4.985 0.75 5.085 0.85 ;
      RECT  3.755 0.75 3.855 0.85 ;
      RECT  3.955 0.75 4.055 0.85 ;
      RECT  2.715 0.75 2.815 0.85 ;
      RECT  2.915 0.75 3.015 0.85 ;
      RECT  1.675 0.75 1.775 0.85 ;
      RECT  1.875 0.75 1.975 0.85 ;
      RECT  0.655 0.75 0.755 0.85 ;
      RECT  0.855 0.75 0.955 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.285 0.755 8.395 0.91 ;
      RECT  7.955 0.91 8.395 1.09 ;
      RECT  7.35 0.74 7.46 0.91 ;
      RECT  7.16 0.91 7.46 1.09 ;
      RECT  6.38 0.755 6.515 0.91 ;
      RECT  6.215 0.91 6.515 1.09 ;
      RECT  5.33 0.75 5.475 0.91 ;
      RECT  5.175 0.91 5.475 1.09 ;
      RECT  4.225 0.785 4.445 0.895 ;
      RECT  4.345 0.895 4.445 0.91 ;
      RECT  4.345 0.91 4.645 1.09 ;
      RECT  3.21 0.785 3.405 0.895 ;
      RECT  3.305 0.895 3.405 0.91 ;
      RECT  3.305 0.91 3.605 1.09 ;
      RECT  2.165 0.785 2.365 0.895 ;
      RECT  2.265 0.895 2.365 0.91 ;
      RECT  2.265 0.91 2.565 1.09 ;
      RECT  1.145 0.785 1.325 0.895 ;
      RECT  1.225 0.895 1.325 0.91 ;
      RECT  1.225 0.91 1.525 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.51 1.09 ;
      LAYER M2 ;
      RECT  0.17 0.95 8.295 1.05 ;
      LAYER V1 ;
      RECT  7.955 0.95 8.055 1.05 ;
      RECT  8.155 0.95 8.255 1.05 ;
      RECT  7.16 0.95 7.26 1.05 ;
      RECT  7.36 0.95 7.46 1.05 ;
      RECT  6.215 0.95 6.315 1.05 ;
      RECT  6.415 0.95 6.515 1.05 ;
      RECT  5.175 0.95 5.275 1.05 ;
      RECT  5.375 0.95 5.475 1.05 ;
      RECT  4.345 0.95 4.445 1.05 ;
      RECT  4.545 0.95 4.645 1.05 ;
      RECT  3.305 0.95 3.405 1.05 ;
      RECT  3.505 0.95 3.605 1.05 ;
      RECT  2.265 0.95 2.365 1.05 ;
      RECT  2.465 0.95 2.565 1.05 ;
      RECT  1.225 0.95 1.325 1.05 ;
      RECT  1.425 0.95 1.525 1.05 ;
      RECT  0.21 0.95 0.31 1.05 ;
      RECT  0.41 0.95 0.51 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.545 0.71 11.65 0.745 ;
      RECT  10.545 0.745 12.65 0.805 ;
      RECT  12.55 0.51 12.65 0.745 ;
      RECT  9.75 0.805 12.65 0.89 ;
      RECT  9.75 0.89 10.72 0.95 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  2.145 1.44 2.265 1.75 ;
      RECT  3.185 1.44 3.305 1.75 ;
      RECT  4.225 1.44 4.345 1.75 ;
      RECT  5.265 1.44 5.385 1.75 ;
      RECT  6.305 1.44 6.425 1.75 ;
      RECT  7.345 1.44 7.455 1.75 ;
      RECT  8.385 1.44 8.505 1.75 ;
      RECT  8.905 1.44 9.025 1.75 ;
      RECT  9.425 1.44 9.545 1.75 ;
      RECT  9.945 1.44 10.065 1.75 ;
      RECT  10.465 1.44 10.585 1.75 ;
      RECT  10.985 1.44 11.105 1.75 ;
      RECT  11.505 1.405 11.625 1.75 ;
      RECT  12.025 1.405 12.145 1.75 ;
      RECT  12.57 1.21 12.69 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  1.885 0.05 2.005 0.36 ;
      RECT  2.405 0.05 2.525 0.36 ;
      RECT  2.925 0.05 3.045 0.36 ;
      RECT  3.445 0.05 3.565 0.36 ;
      RECT  3.965 0.05 4.085 0.36 ;
      RECT  4.485 0.05 4.605 0.36 ;
      RECT  5.005 0.05 5.125 0.36 ;
      RECT  5.525 0.05 5.645 0.36 ;
      RECT  6.045 0.05 6.165 0.36 ;
      RECT  6.565 0.05 6.685 0.36 ;
      RECT  7.085 0.05 7.205 0.36 ;
      RECT  7.605 0.05 7.725 0.36 ;
      RECT  8.125 0.05 8.245 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.04 0.45 11.9 0.54 ;
      RECT  8.62 0.54 11.9 0.56 ;
      RECT  8.62 0.56 12.43 0.62 ;
      RECT  11.75 0.62 12.43 0.655 ;
      RECT  8.62 0.62 10.45 0.695 ;
      RECT  8.62 0.695 9.65 0.725 ;
      RECT  9.35 0.725 9.65 1.06 ;
      RECT  8.55 1.06 12.45 1.18 ;
      RECT  0.75 1.11 1.05 1.18 ;
      RECT  0.53 1.18 12.45 1.29 ;
      RECT  1.75 1.11 2.05 1.18 ;
      RECT  2.75 1.11 3.05 1.18 ;
      RECT  3.75 1.11 4.25 1.18 ;
      RECT  4.75 1.11 5.05 1.18 ;
      RECT  5.75 1.11 6.05 1.18 ;
      RECT  6.75 1.11 7.05 1.18 ;
      RECT  7.55 1.11 7.85 1.18 ;
      RECT  0.53 1.29 11.285 1.35 ;
      LAYER M2 ;
      RECT  0.71 1.15 8.89 1.25 ;
      LAYER V1 ;
      RECT  0.75 1.15 0.85 1.25 ;
      RECT  0.95 1.15 1.05 1.25 ;
      RECT  1.75 1.15 1.85 1.25 ;
      RECT  1.95 1.15 2.05 1.25 ;
      RECT  2.75 1.15 2.85 1.25 ;
      RECT  2.95 1.15 3.05 1.25 ;
      RECT  3.75 1.15 3.85 1.25 ;
      RECT  3.95 1.15 4.05 1.25 ;
      RECT  4.15 1.15 4.25 1.25 ;
      RECT  4.75 1.15 4.85 1.25 ;
      RECT  4.95 1.15 5.05 1.25 ;
      RECT  5.75 1.15 5.85 1.25 ;
      RECT  5.95 1.15 6.05 1.25 ;
      RECT  6.75 1.15 6.85 1.25 ;
      RECT  6.95 1.15 7.05 1.25 ;
      RECT  7.55 1.15 7.65 1.25 ;
      RECT  7.75 1.15 7.85 1.25 ;
      RECT  8.55 1.15 8.65 1.25 ;
      RECT  8.75 1.15 8.85 1.25 ;
    END
    ANTENNADIFFAREA 2.688 ;
  END X
  OBS
      LAYER M1 ;
      RECT  8.345 0.19 12.665 0.34 ;
      RECT  10.51 0.34 12.665 0.36 ;
      RECT  8.345 0.34 8.95 0.45 ;
      RECT  12.0 0.36 12.4 0.45 ;
      RECT  4.205 0.31 4.305 0.45 ;
      RECT  0.065 0.45 8.515 0.62 ;
      RECT  4.73 0.31 4.83 0.45 ;
      RECT  5.255 0.31 5.355 0.45 ;
      RECT  5.78 0.31 5.88 0.45 ;
      RECT  6.305 0.31 6.405 0.45 ;
      RECT  6.83 0.31 6.93 0.45 ;
      RECT  7.35 0.31 7.45 0.45 ;
      RECT  7.855 0.31 7.955 0.45 ;
      LAYER M2 ;
      RECT  4.165 0.35 12.4 0.45 ;
      LAYER V1 ;
      RECT  4.205 0.35 4.305 0.45 ;
      RECT  4.73 0.35 4.83 0.45 ;
      RECT  5.255 0.35 5.355 0.45 ;
      RECT  5.78 0.35 5.88 0.45 ;
      RECT  6.305 0.35 6.405 0.45 ;
      RECT  6.83 0.35 6.93 0.45 ;
      RECT  7.35 0.35 7.45 0.45 ;
      RECT  7.855 0.35 7.955 0.45 ;
      RECT  8.61 0.35 8.71 0.45 ;
      RECT  8.81 0.35 8.91 0.45 ;
      RECT  12.04 0.35 12.14 0.45 ;
      RECT  12.26 0.35 12.36 0.45 ;
  END
END SEN_OAI21_16
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_6
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_6
  CLASS CORE ;
  FOREIGN SEN_OAI21_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.495 0.71 2.795 0.925 ;
      RECT  1.665 0.71 1.965 0.925 ;
      RECT  0.675 0.71 1.015 0.925 ;
      LAYER M2 ;
      RECT  0.675 0.75 3.09 0.85 ;
      LAYER V1 ;
      RECT  2.495 0.75 2.595 0.85 ;
      RECT  2.695 0.75 2.795 0.85 ;
      RECT  1.665 0.75 1.765 0.85 ;
      RECT  1.865 0.75 1.965 0.85 ;
      RECT  0.715 0.75 0.815 0.85 ;
      RECT  0.915 0.75 1.015 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.095 0.73 3.185 0.91 ;
      RECT  2.885 0.91 3.185 1.09 ;
      RECT  2.235 0.73 2.355 0.91 ;
      RECT  2.055 0.91 2.355 1.09 ;
      RECT  1.195 0.72 1.315 0.91 ;
      RECT  1.195 0.91 1.525 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.58 1.09 ;
      LAYER M2 ;
      RECT  0.235 0.95 3.29 1.05 ;
      LAYER V1 ;
      RECT  2.885 0.95 2.985 1.05 ;
      RECT  3.085 0.95 3.185 1.05 ;
      RECT  2.055 0.95 2.155 1.05 ;
      RECT  2.255 0.95 2.355 1.05 ;
      RECT  1.225 0.95 1.325 1.05 ;
      RECT  1.425 0.95 1.525 1.05 ;
      RECT  0.275 0.95 0.375 1.05 ;
      RECT  0.475 0.95 0.575 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 4.85 0.71 ;
      RECT  3.75 0.71 4.85 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.105 1.43 1.225 1.75 ;
      RECT  2.145 1.43 2.265 1.75 ;
      RECT  3.185 1.43 3.305 1.75 ;
      RECT  3.705 1.44 3.825 1.75 ;
      RECT  4.225 1.38 4.345 1.75 ;
      RECT  4.77 1.21 4.89 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.325 0.05 0.445 0.385 ;
      RECT  0.845 0.05 0.965 0.385 ;
      RECT  1.365 0.05 1.485 0.385 ;
      RECT  1.885 0.05 2.005 0.385 ;
      RECT  2.405 0.05 2.525 0.385 ;
      RECT  2.925 0.05 3.045 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.43 4.655 0.515 ;
      RECT  3.445 0.515 4.655 0.56 ;
      RECT  3.445 0.56 3.66 0.69 ;
      RECT  3.53 0.69 3.66 1.11 ;
      RECT  3.35 1.11 4.65 1.2 ;
      RECT  0.75 1.11 1.05 1.2 ;
      RECT  0.535 1.2 4.65 1.29 ;
      RECT  1.75 1.11 1.85 1.2 ;
      RECT  2.55 1.11 2.65 1.2 ;
      RECT  0.535 1.29 3.49 1.34 ;
    END
    ANTENNADIFFAREA 1.008 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.175 0.21 4.915 0.34 ;
      RECT  3.175 0.34 3.305 0.475 ;
      RECT  0.065 0.38 0.185 0.475 ;
      RECT  0.065 0.475 3.305 0.605 ;
  END
END SEN_OAI21_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_8
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_8
  CLASS CORE ;
  FOREIGN SEN_OAI21_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.685 0.71 3.985 0.925 ;
      RECT  2.71 0.71 3.05 0.925 ;
      RECT  1.675 0.71 2.045 0.925 ;
      RECT  0.635 0.71 1.05 0.91 ;
      LAYER M2 ;
      RECT  0.635 0.75 4.29 0.85 ;
      LAYER V1 ;
      RECT  3.685 0.75 3.785 0.85 ;
      RECT  3.885 0.75 3.985 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  1.745 0.75 1.845 0.85 ;
      RECT  1.945 0.75 2.045 0.85 ;
      RECT  0.675 0.75 0.775 0.85 ;
      RECT  0.875 0.75 0.975 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.135 0.755 4.225 0.91 ;
      RECT  4.075 0.91 4.375 1.09 ;
      RECT  3.27 0.735 3.36 0.91 ;
      RECT  3.27 0.91 3.595 1.09 ;
      RECT  2.175 0.745 2.265 0.91 ;
      RECT  2.175 0.91 2.475 1.09 ;
      RECT  1.175 0.72 1.265 0.91 ;
      RECT  1.175 0.91 1.525 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.525 1.09 ;
      LAYER M2 ;
      RECT  0.185 0.95 4.49 1.05 ;
      LAYER V1 ;
      RECT  4.075 0.95 4.175 1.05 ;
      RECT  4.275 0.95 4.375 1.05 ;
      RECT  3.295 0.95 3.395 1.05 ;
      RECT  3.495 0.95 3.595 1.05 ;
      RECT  2.175 0.95 2.275 1.05 ;
      RECT  2.375 0.95 2.475 1.05 ;
      RECT  1.225 0.95 1.325 1.05 ;
      RECT  1.425 0.95 1.525 1.05 ;
      RECT  0.225 0.95 0.325 1.05 ;
      RECT  0.425 0.95 0.525 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.51 6.45 0.71 ;
      RECT  4.95 0.71 6.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  2.145 1.44 2.265 1.75 ;
      RECT  3.185 1.44 3.305 1.75 ;
      RECT  4.225 1.44 4.345 1.75 ;
      RECT  4.745 1.44 4.865 1.75 ;
      RECT  5.265 1.44 5.385 1.75 ;
      RECT  5.785 1.44 5.905 1.75 ;
      RECT  6.33 1.21 6.45 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  1.885 0.05 2.005 0.36 ;
      RECT  2.405 0.05 2.525 0.36 ;
      RECT  2.925 0.05 3.045 0.36 ;
      RECT  3.445 0.05 3.565 0.36 ;
      RECT  3.965 0.05 4.085 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.48 0.46 6.215 0.595 ;
      RECT  4.48 0.595 4.65 1.11 ;
      RECT  4.48 1.11 6.18 1.18 ;
      RECT  0.75 1.11 1.05 1.18 ;
      RECT  0.55 1.18 6.18 1.29 ;
      RECT  1.75 1.11 2.05 1.18 ;
      RECT  2.75 1.11 3.05 1.18 ;
      RECT  3.75 1.11 3.85 1.18 ;
      RECT  0.55 1.29 4.65 1.35 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.195 0.21 6.475 0.34 ;
      RECT  4.195 0.34 4.365 0.45 ;
      RECT  0.065 0.4 0.185 0.45 ;
      RECT  0.065 0.45 4.365 0.62 ;
  END
END SEN_OAI21_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_G_12
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_G_12
  CLASS CORE ;
  FOREIGN SEN_OAI21_G_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.55 0.71 5.855 0.9 ;
      RECT  4.75 0.71 5.05 0.895 ;
      RECT  3.55 0.71 3.85 0.895 ;
      RECT  2.55 0.71 2.85 0.895 ;
      RECT  1.55 0.71 1.85 0.895 ;
      RECT  0.55 0.71 0.85 0.895 ;
      LAYER M2 ;
      RECT  0.51 0.75 5.89 0.85 ;
      LAYER V1 ;
      RECT  5.55 0.75 5.65 0.85 ;
      RECT  5.75 0.75 5.85 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.25 0.91 ;
      RECT  5.95 0.91 6.25 1.09 ;
      RECT  5.35 0.71 5.45 0.91 ;
      RECT  5.15 0.91 5.45 1.09 ;
      RECT  4.15 0.71 4.25 0.91 ;
      RECT  4.15 0.91 4.45 1.09 ;
      RECT  3.15 0.71 3.25 0.91 ;
      RECT  3.15 0.91 3.45 1.09 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  2.15 0.91 2.45 1.09 ;
      RECT  1.15 0.71 1.25 0.91 ;
      RECT  1.15 0.91 1.45 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.45 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.95 6.29 1.05 ;
      LAYER V1 ;
      RECT  5.95 0.95 6.05 1.05 ;
      RECT  6.15 0.95 6.25 1.05 ;
      RECT  5.15 0.95 5.25 1.05 ;
      RECT  5.35 0.95 5.45 1.05 ;
      RECT  4.15 0.95 4.25 1.05 ;
      RECT  4.35 0.95 4.45 1.05 ;
      RECT  3.15 0.95 3.25 1.05 ;
      RECT  3.35 0.95 3.45 1.05 ;
      RECT  2.15 0.95 2.25 1.05 ;
      RECT  2.35 0.95 2.45 1.05 ;
      RECT  1.15 0.95 1.25 1.05 ;
      RECT  1.35 0.95 1.45 1.05 ;
      RECT  0.15 0.95 0.25 1.05 ;
      RECT  0.35 0.95 0.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.515 0.71 9.25 0.895 ;
      RECT  9.15 0.895 9.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.6 1.85 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  2.145 1.44 2.265 1.75 ;
      RECT  3.185 1.44 3.305 1.75 ;
      RECT  4.225 1.44 4.345 1.75 ;
      RECT  5.265 1.44 5.385 1.75 ;
      RECT  6.305 1.44 6.425 1.75 ;
      RECT  6.825 1.385 6.945 1.75 ;
      RECT  7.345 1.385 7.465 1.75 ;
      RECT  7.865 1.385 7.985 1.75 ;
      RECT  8.385 1.385 8.505 1.75 ;
      RECT  8.905 1.385 9.025 1.75 ;
      RECT  9.41 1.41 9.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      RECT  3.445 0.05 3.565 0.36 ;
      RECT  3.965 0.05 4.085 0.36 ;
      RECT  4.485 0.05 4.605 0.36 ;
      RECT  5.005 0.05 5.125 0.36 ;
      RECT  5.525 0.05 5.645 0.36 ;
      RECT  6.045 0.05 6.165 0.36 ;
      RECT  0.325 0.05 0.445 0.41 ;
      RECT  0.845 0.05 0.965 0.41 ;
      RECT  1.365 0.05 1.485 0.41 ;
      RECT  1.885 0.05 2.005 0.41 ;
      RECT  2.405 0.05 2.525 0.41 ;
      RECT  2.925 0.05 3.045 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.45 9.335 0.54 ;
      RECT  6.52 0.54 9.335 0.62 ;
      RECT  6.52 0.62 7.4 0.66 ;
      RECT  7.15 0.66 7.4 1.045 ;
      RECT  6.35 1.045 7.4 1.11 ;
      RECT  6.35 1.11 8.85 1.18 ;
      RECT  3.75 1.11 4.05 1.18 ;
      RECT  3.75 1.18 8.85 1.205 ;
      RECT  4.55 1.11 5.05 1.18 ;
      RECT  5.55 1.11 5.85 1.18 ;
      RECT  3.75 1.205 9.28 1.21 ;
      RECT  2.75 1.11 3.05 1.205 ;
      RECT  0.54 1.205 3.05 1.21 ;
      RECT  0.54 1.21 9.28 1.295 ;
      RECT  0.54 1.295 6.65 1.35 ;
      RECT  9.15 1.295 9.28 1.49 ;
      LAYER M2 ;
      RECT  2.71 1.15 6.89 1.25 ;
      LAYER V1 ;
      RECT  2.75 1.15 2.85 1.25 ;
      RECT  2.95 1.15 3.05 1.25 ;
      RECT  3.75 1.15 3.85 1.25 ;
      RECT  3.95 1.15 4.05 1.25 ;
      RECT  4.55 1.15 4.65 1.25 ;
      RECT  4.75 1.15 4.85 1.25 ;
      RECT  4.95 1.15 5.05 1.25 ;
      RECT  5.55 1.15 5.65 1.25 ;
      RECT  5.75 1.15 5.85 1.25 ;
      RECT  6.35 1.15 6.45 1.25 ;
      RECT  6.55 1.15 6.65 1.25 ;
      RECT  6.75 1.15 6.85 1.25 ;
    END
    ANTENNADIFFAREA 2.016 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.26 0.165 7.48 0.19 ;
      RECT  6.26 0.19 9.545 0.36 ;
      RECT  6.26 0.36 6.89 0.45 ;
      RECT  3.195 0.31 3.295 0.45 ;
      RECT  3.195 0.45 6.43 0.5 ;
      RECT  3.72 0.31 3.82 0.45 ;
      RECT  4.24 0.31 4.34 0.45 ;
      RECT  4.75 0.31 4.85 0.45 ;
      RECT  5.275 0.31 5.375 0.45 ;
      RECT  5.76 0.31 5.86 0.45 ;
      RECT  0.065 0.4 0.185 0.5 ;
      RECT  0.065 0.5 6.43 0.62 ;
      LAYER M2 ;
      RECT  3.155 0.35 6.89 0.45 ;
      LAYER V1 ;
      RECT  3.195 0.35 3.295 0.45 ;
      RECT  3.72 0.35 3.82 0.45 ;
      RECT  4.24 0.35 4.34 0.45 ;
      RECT  4.75 0.35 4.85 0.45 ;
      RECT  5.275 0.35 5.375 0.45 ;
      RECT  5.76 0.35 5.86 0.45 ;
      RECT  6.35 0.35 6.45 0.45 ;
      RECT  6.55 0.35 6.65 0.45 ;
      RECT  6.75 0.35 6.85 0.45 ;
  END
END SEN_OAI21_G_12
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_G_16
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_G_16
  CLASS CORE ;
  FOREIGN SEN_OAI21_G_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.71 8.05 0.895 ;
      RECT  6.755 0.71 7.055 0.9 ;
      RECT  5.75 0.71 6.05 0.9 ;
      RECT  4.75 0.71 5.05 0.9 ;
      RECT  3.55 0.71 3.85 0.895 ;
      RECT  2.55 0.71 2.85 0.895 ;
      RECT  1.55 0.71 1.85 0.895 ;
      RECT  0.55 0.71 0.85 0.895 ;
      LAYER M2 ;
      RECT  0.51 0.75 8.09 0.85 ;
      LAYER V1 ;
      RECT  7.75 0.75 7.85 0.85 ;
      RECT  7.95 0.75 8.05 0.85 ;
      RECT  6.755 0.75 6.855 0.85 ;
      RECT  6.955 0.75 7.055 0.85 ;
      RECT  5.75 0.75 5.85 0.85 ;
      RECT  5.95 0.75 6.05 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.315 0.71 8.45 0.91 ;
      RECT  8.15 0.91 8.45 1.09 ;
      RECT  7.35 0.71 7.45 0.91 ;
      RECT  7.15 0.91 7.45 1.09 ;
      RECT  6.35 0.71 6.45 0.91 ;
      RECT  6.15 0.91 6.45 1.09 ;
      RECT  5.35 0.71 5.45 0.91 ;
      RECT  5.15 0.91 5.45 1.09 ;
      RECT  4.15 0.71 4.25 0.91 ;
      RECT  4.15 0.91 4.45 1.09 ;
      RECT  3.15 0.71 3.25 0.91 ;
      RECT  3.15 0.91 3.45 1.09 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  2.15 0.91 2.45 1.09 ;
      RECT  1.15 0.71 1.25 0.91 ;
      RECT  1.15 0.91 1.45 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.45 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.95 8.49 1.05 ;
      LAYER V1 ;
      RECT  8.15 0.95 8.25 1.05 ;
      RECT  8.35 0.95 8.45 1.05 ;
      RECT  7.15 0.95 7.25 1.05 ;
      RECT  7.35 0.95 7.45 1.05 ;
      RECT  6.15 0.95 6.25 1.05 ;
      RECT  6.35 0.95 6.45 1.05 ;
      RECT  5.15 0.95 5.25 1.05 ;
      RECT  5.35 0.95 5.45 1.05 ;
      RECT  4.15 0.95 4.25 1.05 ;
      RECT  4.35 0.95 4.45 1.05 ;
      RECT  3.15 0.95 3.25 1.05 ;
      RECT  3.35 0.95 3.45 1.05 ;
      RECT  2.15 0.95 2.25 1.05 ;
      RECT  2.35 0.95 2.45 1.05 ;
      RECT  1.15 0.95 1.25 1.05 ;
      RECT  1.35 0.95 1.45 1.05 ;
      RECT  0.15 0.95 0.25 1.05 ;
      RECT  0.35 0.95 0.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.75 0.71 12.65 0.81 ;
      RECT  9.97 0.81 12.65 0.895 ;
      RECT  9.97 0.895 10.94 0.92 ;
      RECT  12.55 0.895 12.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0368 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  2.145 1.44 2.265 1.75 ;
      RECT  3.185 1.44 3.305 1.75 ;
      RECT  4.225 1.44 4.345 1.75 ;
      RECT  5.265 1.44 5.385 1.75 ;
      RECT  6.305 1.44 6.425 1.75 ;
      RECT  7.345 1.44 7.465 1.75 ;
      RECT  8.385 1.44 8.505 1.75 ;
      RECT  8.905 1.44 9.025 1.75 ;
      RECT  9.425 1.44 9.545 1.75 ;
      RECT  9.945 1.44 10.065 1.75 ;
      RECT  10.465 1.44 10.585 1.75 ;
      RECT  10.985 1.38 11.105 1.75 ;
      RECT  11.505 1.38 11.625 1.75 ;
      RECT  12.025 1.38 12.145 1.75 ;
      RECT  12.57 1.21 12.69 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  1.885 0.05 2.005 0.36 ;
      RECT  2.405 0.05 2.525 0.36 ;
      RECT  2.925 0.05 3.045 0.36 ;
      RECT  3.445 0.05 3.565 0.36 ;
      RECT  3.965 0.05 4.085 0.36 ;
      RECT  4.485 0.05 4.605 0.36 ;
      RECT  5.005 0.05 5.125 0.36 ;
      RECT  5.525 0.05 5.645 0.36 ;
      RECT  6.045 0.05 6.165 0.36 ;
      RECT  6.565 0.05 6.685 0.36 ;
      RECT  7.085 0.05 7.205 0.36 ;
      RECT  7.605 0.05 7.725 0.36 ;
      RECT  8.125 0.05 8.245 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.495 0.45 11.415 0.47 ;
      RECT  9.54 0.47 11.415 0.5 ;
      RECT  9.54 0.5 12.455 0.56 ;
      RECT  8.62 0.56 12.455 0.62 ;
      RECT  8.62 0.62 10.65 0.69 ;
      RECT  9.55 0.69 10.65 0.7 ;
      RECT  9.55 0.7 9.87 1.11 ;
      RECT  8.55 1.11 12.45 1.18 ;
      RECT  6.75 1.11 7.05 1.18 ;
      RECT  6.75 1.18 12.45 1.23 ;
      RECT  7.55 1.11 8.05 1.18 ;
      RECT  0.55 1.11 1.05 1.23 ;
      RECT  0.55 1.23 12.45 1.29 ;
      RECT  1.55 1.11 1.85 1.23 ;
      RECT  2.755 1.11 3.055 1.23 ;
      RECT  3.75 1.11 4.05 1.23 ;
      RECT  4.75 1.11 5.05 1.23 ;
      RECT  5.75 1.11 6.05 1.23 ;
      RECT  0.55 1.29 10.65 1.35 ;
      LAYER M2 ;
      RECT  0.71 1.15 10.09 1.25 ;
      LAYER V1 ;
      RECT  0.75 1.15 0.85 1.25 ;
      RECT  0.95 1.15 1.05 1.25 ;
      RECT  1.55 1.15 1.65 1.25 ;
      RECT  1.75 1.15 1.85 1.25 ;
      RECT  2.755 1.15 2.855 1.25 ;
      RECT  2.955 1.15 3.055 1.25 ;
      RECT  3.75 1.15 3.85 1.25 ;
      RECT  3.95 1.15 4.05 1.25 ;
      RECT  4.75 1.15 4.85 1.25 ;
      RECT  4.95 1.15 5.05 1.25 ;
      RECT  5.75 1.15 5.85 1.25 ;
      RECT  5.95 1.15 6.05 1.25 ;
      RECT  6.75 1.15 6.85 1.25 ;
      RECT  6.95 1.15 7.05 1.25 ;
      RECT  7.55 1.15 7.65 1.25 ;
      RECT  7.75 1.15 7.85 1.25 ;
      RECT  7.95 1.15 8.05 1.25 ;
      RECT  8.55 1.15 8.65 1.25 ;
      RECT  8.75 1.15 8.85 1.25 ;
      RECT  8.95 1.15 9.05 1.25 ;
      RECT  9.15 1.15 9.25 1.25 ;
      RECT  9.35 1.15 9.45 1.25 ;
      RECT  9.55 1.15 9.65 1.25 ;
      RECT  9.75 1.15 9.85 1.25 ;
      RECT  9.95 1.15 10.05 1.25 ;
    END
    ANTENNADIFFAREA 2.688 ;
  END X
  OBS
      LAYER M1 ;
      RECT  8.35 0.19 12.66 0.36 ;
      RECT  8.35 0.36 9.4 0.45 ;
      RECT  12.55 0.36 12.66 0.49 ;
      RECT  3.72 0.31 3.82 0.45 ;
      RECT  0.065 0.45 8.53 0.62 ;
      RECT  4.24 0.31 4.34 0.45 ;
      RECT  4.76 0.31 4.86 0.45 ;
      RECT  5.28 0.31 5.38 0.45 ;
      RECT  5.8 0.31 5.9 0.45 ;
      RECT  6.31 0.31 6.41 0.45 ;
      RECT  6.83 0.31 6.93 0.45 ;
      RECT  7.355 0.31 7.455 0.45 ;
      RECT  7.865 0.31 7.965 0.45 ;
      LAYER M2 ;
      RECT  3.68 0.35 12.69 0.45 ;
      LAYER V1 ;
      RECT  3.72 0.35 3.82 0.45 ;
      RECT  4.24 0.35 4.34 0.45 ;
      RECT  4.76 0.35 4.86 0.45 ;
      RECT  5.28 0.35 5.38 0.45 ;
      RECT  5.8 0.35 5.9 0.45 ;
      RECT  6.31 0.35 6.41 0.45 ;
      RECT  6.83 0.35 6.93 0.45 ;
      RECT  7.355 0.35 7.455 0.45 ;
      RECT  7.865 0.35 7.965 0.45 ;
      RECT  8.35 0.35 8.45 0.45 ;
      RECT  8.65 0.35 8.75 0.45 ;
      RECT  8.95 0.35 9.05 0.45 ;
      RECT  9.25 0.35 9.35 0.45 ;
      RECT  12.55 0.35 12.65 0.45 ;
  END
END SEN_OAI21_G_16
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_G_6
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_G_6
  CLASS CORE ;
  FOREIGN SEN_OAI21_G_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.895 ;
      RECT  1.55 0.71 1.85 0.895 ;
      RECT  0.55 0.71 0.85 0.895 ;
      LAYER M2 ;
      RECT  0.51 0.75 2.89 0.85 ;
      LAYER V1 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.14 0.71 3.25 0.91 ;
      RECT  2.95 0.91 3.25 1.09 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  1.95 0.91 2.25 1.09 ;
      RECT  1.15 0.71 1.25 0.91 ;
      RECT  1.15 0.91 1.45 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.45 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.95 3.29 1.05 ;
      LAYER V1 ;
      RECT  2.95 0.95 3.05 1.05 ;
      RECT  3.15 0.95 3.25 1.05 ;
      RECT  1.95 0.95 2.05 1.05 ;
      RECT  2.15 0.95 2.25 1.05 ;
      RECT  1.15 0.95 1.25 1.05 ;
      RECT  1.35 0.95 1.45 1.05 ;
      RECT  0.15 0.95 0.25 1.05 ;
      RECT  0.35 0.95 0.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 4.85 0.71 ;
      RECT  3.77 0.71 4.85 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.105 1.425 1.225 1.75 ;
      RECT  2.145 1.425 2.265 1.75 ;
      RECT  3.185 1.425 3.3 1.75 ;
      RECT  3.72 1.38 3.84 1.75 ;
      RECT  4.24 1.38 4.36 1.75 ;
      RECT  4.79 1.21 4.91 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.325 0.05 0.445 0.4 ;
      RECT  0.845 0.05 0.965 0.4 ;
      RECT  1.365 0.05 1.485 0.4 ;
      RECT  1.885 0.05 2.005 0.4 ;
      RECT  2.405 0.05 2.525 0.4 ;
      RECT  2.925 0.05 3.045 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.41 0.475 4.66 0.595 ;
      RECT  3.54 0.595 3.67 1.11 ;
      RECT  3.35 1.11 4.65 1.205 ;
      RECT  0.535 1.205 4.65 1.29 ;
      RECT  0.535 1.29 3.48 1.335 ;
    END
    ANTENNADIFFAREA 1.008 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.185 0.24 4.93 0.36 ;
      RECT  3.185 0.36 3.315 0.49 ;
      RECT  0.065 0.4 0.185 0.49 ;
      RECT  0.065 0.49 3.315 0.62 ;
  END
END SEN_OAI21_G_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_G_8
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_G_8
  CLASS CORE ;
  FOREIGN SEN_OAI21_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 3.85 0.895 ;
      RECT  2.55 0.71 2.85 0.895 ;
      RECT  1.55 0.71 1.85 0.895 ;
      RECT  0.55 0.71 0.85 0.895 ;
      LAYER M2 ;
      RECT  0.51 0.75 3.89 0.85 ;
      LAYER V1 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.145 0.71 4.265 0.91 ;
      RECT  3.95 0.91 4.265 1.09 ;
      RECT  3.15 0.71 3.25 0.91 ;
      RECT  3.15 0.91 3.45 1.09 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  2.15 0.91 2.45 1.09 ;
      RECT  1.15 0.71 1.25 0.91 ;
      RECT  1.15 0.91 1.45 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.45 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.95 4.29 1.05 ;
      LAYER V1 ;
      RECT  3.95 0.95 4.05 1.05 ;
      RECT  4.15 0.95 4.25 1.05 ;
      RECT  3.15 0.95 3.25 1.05 ;
      RECT  3.35 0.95 3.45 1.05 ;
      RECT  2.15 0.95 2.25 1.05 ;
      RECT  2.35 0.95 2.45 1.05 ;
      RECT  1.15 0.95 1.25 1.05 ;
      RECT  1.35 0.95 1.45 1.05 ;
      RECT  0.15 0.95 0.25 1.05 ;
      RECT  0.35 0.95 0.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.51 6.45 0.71 ;
      RECT  4.825 0.71 6.45 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.105 1.415 1.225 1.75 ;
      RECT  2.145 1.415 2.265 1.75 ;
      RECT  3.185 1.44 3.305 1.75 ;
      RECT  4.225 1.44 4.345 1.75 ;
      RECT  4.745 1.415 4.865 1.75 ;
      RECT  5.265 1.415 5.38 1.75 ;
      RECT  5.785 1.415 5.905 1.75 ;
      RECT  6.34 1.21 6.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  3.445 0.05 3.565 0.36 ;
      RECT  3.965 0.05 4.085 0.36 ;
      RECT  0.325 0.05 0.445 0.4 ;
      RECT  0.845 0.05 0.965 0.4 ;
      RECT  1.365 0.05 1.485 0.4 ;
      RECT  1.885 0.05 2.005 0.4 ;
      RECT  2.405 0.05 2.525 0.4 ;
      RECT  2.925 0.05 3.045 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.485 0.45 6.215 0.58 ;
      RECT  4.485 0.58 4.655 1.11 ;
      RECT  4.485 1.11 6.25 1.18 ;
      RECT  3.75 1.11 3.85 1.18 ;
      RECT  3.75 1.18 6.25 1.205 ;
      RECT  0.535 1.205 6.25 1.29 ;
      RECT  0.535 1.29 4.65 1.325 ;
      RECT  2.54 1.325 4.65 1.35 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.195 0.21 6.495 0.34 ;
      RECT  4.195 0.34 4.365 0.45 ;
      RECT  3.135 0.45 4.365 0.49 ;
      RECT  0.065 0.4 0.185 0.49 ;
      RECT  0.065 0.49 4.365 0.62 ;
  END
END SEN_OAI21_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_S_0P5
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_S_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI21_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.94 1.41 1.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.36 0.05 0.48 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.18 1.06 0.475 ;
      RECT  0.75 0.475 1.06 0.565 ;
      RECT  0.75 0.565 0.85 1.445 ;
      RECT  0.595 1.445 0.85 1.565 ;
    END
    ANTENNADIFFAREA 0.091 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.57 0.23 0.815 0.35 ;
      RECT  0.57 0.35 0.66 0.51 ;
      RECT  0.07 0.185 0.19 0.51 ;
      RECT  0.07 0.51 0.66 0.6 ;
  END
END SEN_OAI21_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_S_1
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_S_1
  CLASS CORE ;
  FOREIGN SEN_OAI21_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.67 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.67 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0543 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0336 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.94 1.41 1.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.35 0.05 0.47 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.94 0.275 1.06 0.51 ;
      RECT  0.75 0.51 1.06 0.6 ;
      RECT  0.75 0.6 0.85 1.44 ;
      RECT  0.595 1.44 0.85 1.56 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.57 0.24 0.815 0.36 ;
      RECT  0.57 0.36 0.66 0.49 ;
      RECT  0.065 0.275 0.185 0.49 ;
      RECT  0.065 0.49 0.66 0.58 ;
  END
END SEN_OAI21_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_S_1P5
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_S_1P5
  CLASS CORE ;
  FOREIGN SEN_OAI21_S_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 0.91 ;
      RECT  0.75 0.91 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.081 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0507 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.37 0.445 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.6 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.87 0.05 0.99 0.41 ;
      RECT  0.3 0.05 0.42 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.43 1.46 1.23 ;
      RECT  0.795 1.23 1.46 1.35 ;
      RECT  1.35 1.35 1.46 1.49 ;
    END
    ANTENNADIFFAREA 0.237 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.12 0.21 1.735 0.3 ;
      RECT  1.615 0.3 1.735 0.43 ;
      RECT  1.12 0.3 1.21 0.5 ;
      RECT  0.535 0.5 1.21 0.62 ;
      RECT  0.065 1.18 0.705 1.27 ;
      RECT  0.065 1.27 0.185 1.4 ;
      RECT  0.585 1.27 0.705 1.44 ;
      RECT  0.585 1.44 1.26 1.56 ;
  END
END SEN_OAI21_S_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_S_2
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_S_2
  CLASS CORE ;
  FOREIGN SEN_OAI21_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1086 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.45 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1086 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0672 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.37 0.435 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.61 1.21 1.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.315 0.05 0.435 0.43 ;
      RECT  0.835 0.05 0.955 0.43 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.335 1.46 1.21 ;
      RECT  0.785 1.21 1.46 1.33 ;
    END
    ANTENNADIFFAREA 0.264 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.095 0.155 1.735 0.245 ;
      RECT  1.615 0.245 1.735 0.42 ;
      RECT  1.095 0.245 1.215 0.52 ;
      RECT  0.055 0.3 0.175 0.52 ;
      RECT  0.055 0.52 1.215 0.61 ;
      RECT  0.575 0.275 0.695 0.52 ;
      RECT  0.055 1.18 0.695 1.27 ;
      RECT  0.575 1.27 0.695 1.43 ;
      RECT  0.055 1.27 0.175 1.615 ;
      RECT  0.575 1.43 1.265 1.55 ;
  END
END SEN_OAI21_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_S_3
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_S_3
  CLASS CORE ;
  FOREIGN SEN_OAI21_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.45 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1632 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1014 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  0.59 1.39 0.71 1.75 ;
      RECT  1.9 1.45 2.02 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.85 0.05 0.97 0.41 ;
      RECT  1.38 0.05 1.5 0.41 ;
      RECT  0.34 0.05 0.45 0.62 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.85 0.465 2.05 0.585 ;
      RECT  1.95 0.585 2.05 1.11 ;
      RECT  1.11 1.11 2.05 1.24 ;
      RECT  1.11 1.24 2.33 1.29 ;
      RECT  1.95 1.29 2.33 1.36 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.64 0.24 2.33 0.36 ;
      RECT  1.64 0.36 1.76 0.5 ;
      RECT  0.54 0.5 1.76 0.62 ;
      RECT  0.28 1.18 0.97 1.3 ;
      RECT  0.85 1.3 0.97 1.44 ;
      RECT  0.85 1.44 1.54 1.56 ;
  END
END SEN_OAI21_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_S_4
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_S_4
  CLASS CORE ;
  FOREIGN SEN_OAI21_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.85 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2169 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2169 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.54 0.71 3.05 0.895 ;
      RECT  2.95 0.895 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1341 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.33 1.39 0.45 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  0.85 1.39 0.97 1.75 ;
      RECT  2.4 1.38 2.52 1.75 ;
      RECT  2.94 1.21 3.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.67 0.05 0.79 0.38 ;
      RECT  1.24 0.05 1.36 0.38 ;
      RECT  1.805 0.05 1.925 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.28 0.45 3.045 0.57 ;
      RECT  2.35 0.57 2.45 1.11 ;
      RECT  1.345 1.11 2.85 1.29 ;
    END
    ANTENNADIFFAREA 0.505 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.07 0.24 2.76 0.36 ;
      RECT  2.07 0.36 2.19 0.47 ;
      RECT  0.36 0.47 2.19 0.59 ;
      RECT  0.07 1.18 1.235 1.3 ;
      RECT  0.07 1.3 0.19 1.4 ;
      RECT  1.105 1.3 1.235 1.44 ;
      RECT  1.105 1.44 2.31 1.56 ;
  END
END SEN_OAI21_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_S_8
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_S_8
  CLASS CORE ;
  FOREIGN SEN_OAI21_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.665 3.46 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4338 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.65 0.905 ;
      RECT  0.55 0.905 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4338 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.51 5.05 0.71 ;
      RECT  4.15 0.71 5.05 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2682 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.39 0.445 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.845 1.39 0.965 1.75 ;
      RECT  1.365 1.39 1.485 1.75 ;
      RECT  1.885 1.41 2.005 1.75 ;
      RECT  4.235 1.38 4.355 1.75 ;
      RECT  4.755 1.38 4.875 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  2.12 0.05 2.29 0.31 ;
      RECT  2.64 0.05 2.815 0.31 ;
      RECT  3.16 0.05 3.33 0.31 ;
      RECT  0.585 0.05 0.705 0.395 ;
      RECT  1.105 0.05 1.225 0.395 ;
      RECT  1.625 0.05 1.745 0.395 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.68 0.45 4.86 0.575 ;
      RECT  4.755 0.575 4.86 0.62 ;
      RECT  3.68 0.575 3.85 1.105 ;
      RECT  3.68 1.105 5.135 1.11 ;
      RECT  2.35 1.11 5.135 1.29 ;
    END
    ANTENNADIFFAREA 0.966 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.015 0.165 5.135 0.24 ;
      RECT  3.455 0.24 5.135 0.36 ;
      RECT  3.455 0.36 3.575 0.4 ;
      RECT  1.86 0.4 3.575 0.485 ;
      RECT  0.275 0.485 3.575 0.52 ;
      RECT  0.275 0.52 1.99 0.605 ;
      RECT  0.065 1.18 2.26 1.3 ;
      RECT  1.565 1.3 2.26 1.32 ;
      RECT  0.065 1.3 0.185 1.4 ;
      RECT  2.12 1.32 2.26 1.42 ;
      RECT  2.12 1.42 2.81 1.44 ;
      RECT  2.12 1.44 3.875 1.56 ;
  END
END SEN_OAI21_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_0P75
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_0P75
  CLASS CORE ;
  FOREIGN SEN_OAI21_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0471 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.2 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.94 1.41 1.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.325 0.05 0.445 0.43 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.425 1.04 0.54 ;
      RECT  0.75 0.54 0.85 1.31 ;
      RECT  0.55 1.31 0.85 1.49 ;
    END
    ANTENNADIFFAREA 0.163 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.535 0.215 0.755 0.335 ;
      RECT  0.535 0.335 0.625 0.53 ;
      RECT  0.065 0.325 0.185 0.53 ;
      RECT  0.065 0.53 0.625 0.62 ;
  END
END SEN_OAI21_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_5
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_5
  CLASS CORE ;
  FOREIGN SEN_OAI21_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 2.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3165 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.585 1.39 0.705 1.75 ;
      RECT  1.105 1.39 1.225 1.75 ;
      RECT  2.925 1.38 3.045 1.75 ;
      RECT  3.445 1.38 3.565 1.75 ;
      RECT  3.98 1.21 4.1 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.325 0.05 0.445 0.4 ;
      RECT  0.845 0.05 0.965 0.4 ;
      RECT  1.365 0.05 1.485 0.4 ;
      RECT  1.885 0.05 2.005 0.4 ;
      RECT  2.405 0.05 2.525 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.31 4.085 0.475 ;
      RECT  2.9 0.475 4.085 0.595 ;
      RECT  3.15 0.595 3.26 1.11 ;
      RECT  1.575 1.11 3.86 1.29 ;
    END
    ANTENNADIFFAREA 0.859 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.665 0.26 3.86 0.38 ;
      RECT  2.665 0.38 2.785 0.49 ;
      RECT  0.065 0.39 0.185 0.49 ;
      RECT  0.065 0.49 2.785 0.61 ;
      RECT  0.275 1.18 1.485 1.3 ;
      RECT  1.365 1.3 1.485 1.425 ;
      RECT  1.365 1.425 2.575 1.545 ;
  END
END SEN_OAI21_5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_T_0P5
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_T_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI21_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 0.9 ;
      RECT  0.35 0.9 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0315 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.875 1.41 1.005 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.845 0.21 0.965 0.51 ;
      RECT  0.75 0.51 0.965 0.6 ;
      RECT  0.75 0.6 0.85 1.21 ;
      RECT  0.55 1.21 0.85 1.3 ;
      RECT  0.55 1.3 0.705 1.49 ;
    END
    ANTENNADIFFAREA 0.097 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.54 0.215 0.755 0.335 ;
      RECT  0.54 0.335 0.63 0.475 ;
      RECT  0.065 0.32 0.185 0.475 ;
      RECT  0.065 0.475 0.63 0.565 ;
  END
END SEN_OAI21_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_T_1
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_T_1
  CLASS CORE ;
  FOREIGN SEN_OAI21_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.315 0.925 ;
      RECT  1.15 0.925 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0633 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.305 1.21 0.425 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.38 1.41 1.51 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.495 0.49 ;
      RECT  1.405 0.49 1.495 1.11 ;
      RECT  1.35 1.11 1.495 1.2 ;
      RECT  1.105 1.2 1.495 1.29 ;
      RECT  1.105 1.29 1.25 1.49 ;
    END
    ANTENNADIFFAREA 0.195 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 1.225 0.59 ;
      RECT  1.105 0.37 1.225 0.48 ;
  END
END SEN_OAI21_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_T_2
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_T_2
  CLASS CORE ;
  FOREIGN SEN_OAI21_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.91 ;
      RECT  0.95 0.91 1.85 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1872 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.85 0.9 ;
      RECT  0.15 0.9 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1872 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.45 0.91 ;
      RECT  2.15 0.91 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1266 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.39 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.6 1.495 1.77 1.75 ;
      RECT  2.12 1.495 2.29 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.1 0.05 1.23 0.385 ;
      RECT  1.62 0.05 1.75 0.385 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.39 2.25 0.71 ;
      RECT  1.95 0.71 2.25 0.8 ;
      RECT  1.95 0.8 2.05 1.315 ;
      RECT  0.82 1.235 1.485 1.315 ;
      RECT  0.82 1.315 2.525 1.36 ;
      RECT  1.365 1.36 2.525 1.405 ;
      RECT  2.405 1.405 2.525 1.535 ;
      RECT  1.365 1.405 1.485 1.55 ;
      RECT  1.885 1.405 2.005 1.55 ;
    END
    ANTENNADIFFAREA 0.353 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.885 0.21 2.525 0.3 ;
      RECT  2.405 0.3 2.525 0.43 ;
      RECT  1.885 0.3 2.005 0.475 ;
      RECT  0.275 0.475 2.005 0.6 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.185 1.435 ;
      RECT  0.585 1.3 0.705 1.48 ;
      RECT  0.585 1.48 1.275 1.6 ;
  END
END SEN_OAI21_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_T_3
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_T_3
  CLASS CORE ;
  FOREIGN SEN_OAI21_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.45 0.91 ;
      RECT  1.55 0.91 2.45 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 0.91 ;
      RECT  0.55 0.91 1.45 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1899 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.56 1.465 0.73 1.75 ;
      RECT  1.08 1.465 1.25 1.75 ;
      RECT  2.94 1.42 3.05 1.75 ;
      RECT  3.48 1.21 3.6 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  1.88 0.05 2.01 0.385 ;
      RECT  2.4 0.05 2.53 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.445 0.32 3.565 0.45 ;
      RECT  2.94 0.45 3.565 0.54 ;
      RECT  2.94 0.54 3.05 1.21 ;
      RECT  2.68 1.21 3.355 1.33 ;
      RECT  2.68 1.33 2.85 1.465 ;
      RECT  1.575 1.465 2.85 1.58 ;
    END
    ANTENNADIFFAREA 0.527 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.665 0.215 3.355 0.335 ;
      RECT  2.665 0.335 2.785 0.475 ;
      RECT  0.065 0.375 0.185 0.475 ;
      RECT  0.065 0.475 2.785 0.595 ;
      RECT  0.275 1.255 2.575 1.375 ;
  END
END SEN_OAI21_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_T_4
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_T_4
  CLASS CORE ;
  FOREIGN SEN_OAI21_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 3.45 0.91 ;
      RECT  2.35 0.91 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 0.91 ;
      RECT  0.55 0.91 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.85 0.905 ;
      RECT  4.75 0.905 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2532 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.54 1.415 0.67 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.1 1.415 1.23 1.75 ;
      RECT  1.62 1.415 1.75 1.75 ;
      RECT  3.71 1.44 3.83 1.75 ;
      RECT  4.22 1.41 4.35 1.75 ;
      RECT  4.765 1.21 4.885 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  1.88 0.05 2.01 0.385 ;
      RECT  2.4 0.05 2.53 0.385 ;
      RECT  2.92 0.05 3.05 0.385 ;
      RECT  3.44 0.05 3.57 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.94 0.45 4.655 0.57 ;
      RECT  3.94 0.57 4.06 1.11 ;
      RECT  3.94 1.11 4.65 1.23 ;
      RECT  2.11 1.23 4.65 1.29 ;
      RECT  2.11 1.29 4.05 1.35 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.705 0.24 4.915 0.36 ;
      RECT  3.705 0.36 3.825 0.475 ;
      RECT  0.065 0.375 0.185 0.475 ;
      RECT  0.065 0.475 3.825 0.595 ;
      RECT  0.35 1.205 2.0 1.325 ;
      RECT  0.35 1.325 0.45 1.4 ;
      RECT  1.885 1.325 2.0 1.44 ;
      RECT  0.065 1.4 0.45 1.57 ;
      RECT  1.885 1.44 3.62 1.56 ;
  END
END SEN_OAI21_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_T_6
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_T_6
  CLASS CORE ;
  FOREIGN SEN_OAI21_T_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.71 5.05 0.91 ;
      RECT  3.15 0.91 5.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5616 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.91 2.05 1.095 ;
      RECT  0.15 1.095 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5616 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.51 7.05 0.71 ;
      RECT  5.935 0.71 7.05 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3798 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 7.2 1.85 ;
      RECT  0.615 1.415 0.745 1.75 ;
      RECT  1.205 1.415 1.335 1.75 ;
      RECT  1.81 1.415 1.94 1.75 ;
      RECT  2.385 1.415 2.515 1.75 ;
      RECT  5.595 1.41 5.725 1.75 ;
      RECT  6.115 1.41 6.245 1.75 ;
      RECT  6.635 1.41 6.765 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      RECT  0.32 0.05 0.45 0.375 ;
      RECT  5.075 0.05 5.205 0.395 ;
      RECT  0.845 0.05 0.965 0.585 ;
      RECT  1.365 0.05 1.485 0.585 ;
      RECT  1.885 0.05 2.005 0.585 ;
      RECT  2.405 0.05 2.525 0.585 ;
      RECT  3.0 0.05 3.12 0.585 ;
      RECT  3.52 0.05 3.64 0.585 ;
      RECT  4.04 0.05 4.16 0.585 ;
      RECT  4.56 0.05 4.665 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.535 0.45 6.81 0.58 ;
      RECT  5.535 0.58 5.665 1.11 ;
      RECT  5.34 1.11 7.05 1.235 ;
      RECT  2.975 1.235 7.05 1.29 ;
      RECT  2.975 1.29 5.46 1.365 ;
    END
    ANTENNADIFFAREA 1.092 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.315 0.23 7.07 0.36 ;
      RECT  5.315 0.36 5.445 0.485 ;
      RECT  4.755 0.485 5.445 0.615 ;
      RECT  4.755 0.615 4.86 0.675 ;
      RECT  0.065 0.375 0.185 0.465 ;
      RECT  0.065 0.465 0.735 0.595 ;
      RECT  0.605 0.595 0.735 0.675 ;
      RECT  0.605 0.675 4.86 0.805 ;
      RECT  0.34 1.2 2.83 1.325 ;
      RECT  0.34 1.325 0.46 1.43 ;
      RECT  2.695 1.325 2.83 1.455 ;
      RECT  2.695 1.455 5.24 1.585 ;
  END
END SEN_OAI21_T_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_T_8
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_T_8
  CLASS CORE ;
  FOREIGN SEN_OAI21_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.71 6.05 0.91 ;
      RECT  3.55 0.91 6.05 1.095 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7488 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.75 0.91 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7488 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.06 0.71 8.65 0.905 ;
      RECT  8.55 0.905 8.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5064 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.3 1.445 0.47 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  0.82 1.445 0.99 1.75 ;
      RECT  1.34 1.445 1.51 1.75 ;
      RECT  1.86 1.445 2.03 1.75 ;
      RECT  2.38 1.445 2.55 1.75 ;
      RECT  2.9 1.445 3.07 1.75 ;
      RECT  6.515 1.12 6.635 1.75 ;
      RECT  7.025 1.41 7.155 1.75 ;
      RECT  7.545 1.41 7.675 1.75 ;
      RECT  8.065 1.41 8.195 1.75 ;
      RECT  8.6 1.21 8.72 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  0.84 0.05 0.97 0.36 ;
      RECT  1.36 0.05 1.49 0.36 ;
      RECT  1.88 0.05 2.01 0.36 ;
      RECT  2.4 0.05 2.53 0.36 ;
      RECT  2.92 0.05 3.05 0.36 ;
      RECT  3.44 0.05 3.57 0.36 ;
      RECT  3.96 0.05 4.09 0.36 ;
      RECT  4.48 0.05 4.61 0.36 ;
      RECT  5.0 0.05 5.13 0.36 ;
      RECT  5.52 0.05 5.65 0.36 ;
      RECT  6.04 0.05 6.17 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.745 0.45 8.5 0.62 ;
      RECT  6.745 0.62 6.925 0.71 ;
      RECT  6.14 0.71 6.925 0.89 ;
      RECT  6.75 0.89 6.925 1.11 ;
      RECT  6.14 0.89 6.31 1.185 ;
      RECT  6.75 1.11 8.45 1.29 ;
      RECT  3.42 1.185 6.31 1.345 ;
    END
    ANTENNADIFFAREA 1.328 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.47 0.19 8.71 0.36 ;
      RECT  8.59 0.36 8.71 0.43 ;
      RECT  6.47 0.36 6.64 0.45 ;
      RECT  0.065 0.4 0.185 0.45 ;
      RECT  0.065 0.45 6.64 0.62 ;
      RECT  0.065 1.185 3.33 1.355 ;
      RECT  0.065 1.355 0.185 1.43 ;
      RECT  3.16 1.355 3.33 1.435 ;
      RECT  3.16 1.435 6.425 1.615 ;
  END
END SEN_OAI21_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_G_0P5
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_G_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI21_G_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.91 ;
      RECT  0.35 0.91 0.45 1.135 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.94 1.41 1.07 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.845 0.26 1.05 0.45 ;
      RECT  0.75 0.45 1.05 0.54 ;
      RECT  0.75 0.54 0.85 1.31 ;
      RECT  0.55 1.31 0.85 1.49 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.54 0.215 0.755 0.335 ;
      RECT  0.54 0.335 0.63 0.45 ;
      RECT  0.065 0.21 0.19 0.45 ;
      RECT  0.065 0.45 0.63 0.54 ;
  END
END SEN_OAI21_G_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_G_1
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_G_1
  CLASS CORE ;
  FOREIGN SEN_OAI21_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.915 1.41 1.045 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.32 0.05 0.45 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.845 0.31 1.05 0.45 ;
      RECT  0.75 0.45 1.05 0.55 ;
      RECT  0.75 0.55 0.85 1.11 ;
      RECT  0.55 1.11 0.85 1.29 ;
    END
    ANTENNADIFFAREA 0.197 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.555 0.24 0.755 0.36 ;
      RECT  0.555 0.36 0.645 0.495 ;
      RECT  0.065 0.365 0.185 0.495 ;
      RECT  0.065 0.495 0.645 0.585 ;
  END
END SEN_OAI21_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_G_2
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_G_2
  CLASS CORE ;
  FOREIGN SEN_OAI21_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.9 ;
      RECT  0.75 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.245 1.22 1.445 1.34 ;
      RECT  1.34 1.34 1.445 1.75 ;
      RECT  0.325 1.19 0.445 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.81 1.41 1.94 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.58 0.05 0.71 0.385 ;
      RECT  1.1 0.05 1.22 0.385 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.32 1.675 0.555 ;
      RECT  1.55 0.555 1.65 1.04 ;
      RECT  0.95 1.04 1.65 1.13 ;
      RECT  0.95 1.13 1.05 1.24 ;
      RECT  1.55 1.13 1.65 1.34 ;
      RECT  0.795 1.24 1.05 1.36 ;
      RECT  1.55 1.34 1.675 1.54 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.31 0.14 1.93 0.23 ;
      RECT  1.815 0.23 1.93 0.43 ;
      RECT  1.31 0.23 1.415 0.475 ;
      RECT  0.34 0.38 0.445 0.475 ;
      RECT  0.34 0.475 1.415 0.6 ;
      RECT  1.295 0.6 1.415 0.715 ;
      RECT  0.065 0.99 0.65 1.08 ;
      RECT  0.065 1.08 0.185 1.22 ;
      RECT  0.56 1.08 0.65 1.46 ;
      RECT  0.56 1.46 1.25 1.58 ;
  END
END SEN_OAI21_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21_G_4
#      Description : "One 2-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21_G_4
  CLASS CORE ;
  FOREIGN SEN_OAI21_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.45 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.285 1.225 2.48 1.345 ;
      RECT  2.39 1.345 2.48 1.75 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  2.855 1.23 2.975 1.75 ;
      RECT  3.39 1.21 3.51 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.41 0.05 1.54 0.385 ;
      RECT  2.03 0.05 2.16 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.44 3.285 0.56 ;
      RECT  2.55 0.56 2.65 1.015 ;
      RECT  1.95 1.015 3.25 1.135 ;
      RECT  1.95 1.135 2.05 1.24 ;
      RECT  3.115 1.135 3.25 1.49 ;
      RECT  1.315 1.24 2.05 1.36 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.335 0.215 3.495 0.335 ;
      RECT  3.375 0.335 3.495 0.435 ;
      RECT  2.335 0.335 2.455 0.475 ;
      RECT  0.065 0.375 0.185 0.475 ;
      RECT  0.065 0.475 2.455 0.595 ;
      RECT  0.065 1.205 1.225 1.325 ;
      RECT  0.065 1.325 0.185 1.425 ;
      RECT  1.105 1.325 1.225 1.46 ;
      RECT  1.105 1.46 2.3 1.58 ;
  END
END SEN_OAI21_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21B_0P5
#      Description : "One 2-input OR into 2-input NAND (other input inverted)"
#      Equation    : X=!((A1|A2)&!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21B_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI21B_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.705 0.65 0.91 ;
      RECT  0.35 0.91 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0198 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  0.845 1.41 0.975 1.75 ;
      RECT  1.375 1.415 1.505 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.325 0.05 0.455 0.365 ;
      RECT  1.375 0.05 1.505 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.85 0.2 0.97 0.635 ;
      RECT  0.75 0.635 0.97 0.725 ;
      RECT  0.75 0.725 0.85 1.11 ;
      RECT  0.55 1.11 0.85 1.29 ;
      RECT  0.55 1.29 0.71 1.49 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.21 0.19 0.455 ;
      RECT  0.07 0.455 0.71 0.545 ;
      RECT  0.59 0.21 0.71 0.455 ;
      RECT  1.115 0.18 1.235 0.815 ;
      RECT  0.98 0.815 1.235 0.925 ;
      RECT  1.115 0.925 1.235 1.63 ;
  END
END SEN_OAI21B_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21B_1
#      Description : "One 2-input OR into 2-input NAND (other input inverted)"
#      Equation    : X=!((A1|A2)&!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21B_1
  CLASS CORE ;
  FOREIGN SEN_OAI21B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.7 0.65 1.54 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.5 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0294 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.15 1.41 0.28 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.08 1.41 1.21 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.365 0.05 0.495 0.39 ;
      RECT  1.41 0.05 1.54 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.855 0.5 1.05 0.69 ;
      RECT  0.855 0.69 0.945 0.71 ;
      RECT  0.75 0.71 0.945 0.81 ;
      RECT  0.75 0.81 0.85 1.3 ;
    END
    ANTENNADIFFAREA 0.213 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.095 0.37 0.215 0.5 ;
      RECT  0.095 0.5 0.765 0.59 ;
      RECT  0.645 0.37 0.765 0.5 ;
      RECT  1.155 0.21 1.26 0.78 ;
      RECT  1.035 0.78 1.26 0.9 ;
      RECT  1.155 0.9 1.26 1.21 ;
      RECT  1.155 1.21 1.535 1.3 ;
      RECT  1.415 1.3 1.535 1.58 ;
  END
END SEN_OAI21B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21B_2
#      Description : "One 2-input OR into 2-input NAND (other input inverted)"
#      Equation    : X=!((A1|A2)&!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21B_2
  CLASS CORE ;
  FOREIGN SEN_OAI21B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.7 1.06 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.5 2.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0588 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.42 1.41 1.55 1.75 ;
      RECT  1.95 1.41 2.08 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.32 0.05 0.49 0.39 ;
      RECT  0.87 0.05 0.995 0.39 ;
      RECT  2.19 0.05 2.32 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.565 0.695 ;
      RECT  1.35 0.695 1.45 1.11 ;
      RECT  0.84 1.11 1.85 1.29 ;
    END
    ANTENNADIFFAREA 0.334 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.14 0.19 1.78 0.28 ;
      RECT  1.66 0.28 1.78 0.44 ;
      RECT  1.14 0.28 1.26 0.49 ;
      RECT  0.065 0.37 0.185 0.49 ;
      RECT  0.065 0.49 1.26 0.59 ;
      RECT  1.93 0.44 2.04 0.79 ;
      RECT  1.6 0.79 2.04 0.89 ;
      RECT  1.95 0.89 2.04 1.21 ;
      RECT  1.95 1.21 2.335 1.3 ;
      RECT  2.215 1.3 2.335 1.43 ;
      RECT  0.065 1.21 0.72 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.6 1.3 0.72 1.52 ;
      RECT  0.6 1.52 1.265 1.61 ;
      RECT  1.145 1.38 1.265 1.52 ;
  END
END SEN_OAI21B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21B_3
#      Description : "One 2-input OR into 2-input NAND (other input inverted)"
#      Equation    : X=!((A1|A2)&!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21B_3
  CLASS CORE ;
  FOREIGN SEN_OAI21B_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.7 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.7 3.25 0.89 ;
      RECT  2.95 0.89 3.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0882 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.61 1.21 0.73 1.75 ;
      RECT  1.965 1.41 2.095 1.75 ;
      RECT  2.555 1.21 2.665 1.75 ;
      RECT  3.14 1.21 3.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.335 0.05 0.465 0.39 ;
      RECT  0.87 0.05 1.0 0.39 ;
      RECT  1.395 0.05 1.525 0.39 ;
      RECT  2.69 0.05 2.82 0.39 ;
      RECT  3.215 0.05 3.335 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.895 0.51 2.65 0.7 ;
      RECT  1.95 0.7 2.05 1.11 ;
      RECT  1.35 1.11 2.45 1.21 ;
      RECT  1.115 1.21 2.45 1.29 ;
      RECT  1.115 1.29 1.45 1.31 ;
    END
    ANTENNADIFFAREA 0.536 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.66 0.25 2.35 0.35 ;
      RECT  1.66 0.35 1.78 0.49 ;
      RECT  0.065 0.37 0.185 0.49 ;
      RECT  0.065 0.49 1.78 0.59 ;
      RECT  2.955 0.33 3.075 0.5 ;
      RECT  2.755 0.5 3.075 0.59 ;
      RECT  2.755 0.59 2.845 0.79 ;
      RECT  2.185 0.79 2.845 0.89 ;
      RECT  2.755 0.89 2.845 1.21 ;
      RECT  2.755 1.21 2.975 1.3 ;
      RECT  2.855 1.3 2.975 1.45 ;
      RECT  0.35 1.01 0.995 1.1 ;
      RECT  0.35 1.1 0.45 1.25 ;
      RECT  0.875 1.1 0.995 1.46 ;
      RECT  0.875 1.46 1.57 1.56 ;
  END
END SEN_OAI21B_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21B_4
#      Description : "One 2-input OR into 2-input NAND (other input inverted)"
#      Equation    : X=!((A1|A2)&!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21B_4
  CLASS CORE ;
  FOREIGN SEN_OAI21B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.7 4.05 0.89 ;
      RECT  3.95 0.89 4.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1176 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.335 1.41 0.465 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  0.87 1.21 1.0 1.75 ;
      RECT  2.43 1.21 2.55 1.75 ;
      RECT  2.945 1.38 3.075 1.75 ;
      RECT  3.47 1.21 3.6 1.75 ;
      RECT  4.01 1.21 4.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  0.335 0.05 0.465 0.39 ;
      RECT  0.87 0.05 1.0 0.39 ;
      RECT  1.395 0.05 1.525 0.39 ;
      RECT  1.92 0.05 2.04 0.39 ;
      RECT  3.475 0.05 3.605 0.39 ;
      RECT  4.015 0.05 4.135 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.415 0.51 3.105 0.69 ;
      RECT  2.75 0.69 2.85 0.91 ;
      RECT  1.95 0.91 2.85 1.1 ;
      RECT  1.95 1.1 2.065 1.11 ;
      RECT  2.655 1.1 2.85 1.11 ;
      RECT  1.55 1.11 2.065 1.21 ;
      RECT  2.655 1.11 3.36 1.29 ;
      RECT  1.375 1.21 2.065 1.31 ;
    END
    ANTENNADIFFAREA 0.668 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.18 0.28 3.34 0.38 ;
      RECT  2.18 0.38 2.3 0.48 ;
      RECT  3.22 0.38 3.34 0.5 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 2.3 0.59 ;
      RECT  3.74 0.37 3.86 0.5 ;
      RECT  3.555 0.5 3.86 0.59 ;
      RECT  3.555 0.59 3.645 0.79 ;
      RECT  2.99 0.79 3.645 0.89 ;
      RECT  3.555 0.89 3.645 1.01 ;
      RECT  3.555 1.01 3.86 1.1 ;
      RECT  3.74 1.1 3.86 1.33 ;
      RECT  0.61 1.01 1.25 1.12 ;
      RECT  0.61 1.12 0.74 1.21 ;
      RECT  1.15 1.12 1.25 1.46 ;
      RECT  0.065 1.21 0.74 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  1.15 1.46 2.3 1.56 ;
      RECT  2.18 1.34 2.3 1.46 ;
  END
END SEN_OAI21B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21B_6
#      Description : "One 2-input OR into 2-input NAND (other input inverted)"
#      Equation    : X=!((A1|A2)&!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21B_6
  CLASS CORE ;
  FOREIGN SEN_OAI21B_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 0.71 ;
      RECT  0.95 0.71 2.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.91 ;
      RECT  0.55 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1602 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.455 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.86 1.44 0.99 1.75 ;
      RECT  1.395 1.45 1.525 1.75 ;
      RECT  1.915 1.45 2.045 1.75 ;
      RECT  2.415 1.45 2.585 1.75 ;
      RECT  2.945 1.45 3.075 1.75 ;
      RECT  3.465 1.45 3.595 1.75 ;
      RECT  3.985 1.45 4.115 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  0.325 0.05 0.455 0.36 ;
      RECT  0.865 0.05 0.995 0.36 ;
      RECT  1.395 0.05 1.525 0.36 ;
      RECT  1.915 0.05 2.045 0.36 ;
      RECT  2.435 0.05 2.565 0.36 ;
      RECT  4.505 0.05 4.635 0.36 ;
      RECT  5.025 0.05 5.155 0.36 ;
      RECT  5.545 0.05 5.675 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.905 0.51 4.14 0.63 ;
      RECT  2.905 0.63 4.05 0.69 ;
      RECT  3.92 0.69 4.05 0.91 ;
      RECT  3.92 0.91 4.65 1.01 ;
      RECT  2.64 1.01 4.65 1.12 ;
      RECT  4.53 1.12 4.65 1.24 ;
      RECT  4.53 1.24 5.93 1.36 ;
      RECT  5.81 1.36 5.93 1.46 ;
    END
    ANTENNADIFFAREA 1.08 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.685 0.215 4.375 0.345 ;
      RECT  2.685 0.345 2.815 0.45 ;
      RECT  4.245 0.345 4.375 0.46 ;
      RECT  1.14 0.36 1.26 0.45 ;
      RECT  1.14 0.45 2.815 0.58 ;
      RECT  4.245 0.46 5.93 0.58 ;
      RECT  5.81 0.36 5.93 0.46 ;
      RECT  2.45 0.79 3.825 0.89 ;
      RECT  2.45 0.89 2.55 1.04 ;
      RECT  0.07 0.35 0.19 0.45 ;
      RECT  0.07 0.45 0.86 0.57 ;
      RECT  0.77 0.57 0.86 1.04 ;
      RECT  0.77 1.04 2.55 1.13 ;
      RECT  0.77 1.13 0.86 1.23 ;
      RECT  0.07 1.23 0.86 1.35 ;
      RECT  0.07 1.35 0.19 1.45 ;
      RECT  1.09 1.23 4.385 1.36 ;
      RECT  4.24 1.36 4.385 1.455 ;
      RECT  4.24 1.455 5.72 1.585 ;
  END
END SEN_OAI21B_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI21B_8
#      Description : "One 2-input OR into 2-input NAND (other input inverted)"
#      Equation    : X=!((A1|A2)&!B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI21B_8
  CLASS CORE ;
  FOREIGN SEN_OAI21B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 5.45 0.89 ;
      RECT  5.35 0.89 5.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.71 7.45 0.89 ;
      RECT  7.35 0.89 7.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2052 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.455 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.945 1.44 1.075 1.75 ;
      RECT  1.625 1.41 1.755 1.75 ;
      RECT  2.145 1.41 2.275 1.75 ;
      RECT  2.665 1.41 2.795 1.75 ;
      RECT  3.185 1.41 3.315 1.75 ;
      RECT  5.775 1.44 5.905 1.75 ;
      RECT  6.295 1.44 6.425 1.75 ;
      RECT  6.815 1.44 6.945 1.75 ;
      RECT  7.335 1.44 7.465 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  0.585 0.05 0.715 0.36 ;
      RECT  1.105 0.05 1.235 0.36 ;
      RECT  3.695 0.05 3.825 0.36 ;
      RECT  4.215 0.05 4.345 0.36 ;
      RECT  4.735 0.05 4.865 0.36 ;
      RECT  5.255 0.05 5.385 0.36 ;
      RECT  5.775 0.05 5.905 0.36 ;
      RECT  6.295 0.05 6.425 0.36 ;
      RECT  6.815 0.05 6.945 0.36 ;
      RECT  7.335 0.05 7.465 0.36 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 3.32 0.69 ;
      RECT  3.15 0.69 3.32 1.11 ;
      RECT  1.345 1.11 4.25 1.22 ;
      RECT  1.345 1.22 5.425 1.29 ;
      RECT  4.135 1.29 5.425 1.35 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.89 0.205 3.585 0.23 ;
      RECT  1.36 0.23 3.585 0.36 ;
      RECT  1.36 0.36 1.48 0.45 ;
      RECT  3.415 0.36 3.585 0.45 ;
      RECT  3.415 0.45 7.72 0.58 ;
      RECT  7.6 0.36 7.72 0.45 ;
      RECT  3.415 0.58 6.185 0.62 ;
      RECT  0.28 0.45 1.24 0.57 ;
      RECT  1.15 0.57 1.24 0.78 ;
      RECT  1.15 0.78 2.965 0.905 ;
      RECT  1.15 0.905 1.24 1.23 ;
      RECT  0.07 1.23 1.24 1.35 ;
      RECT  0.07 1.35 0.19 1.45 ;
      RECT  5.515 1.2 6.195 1.23 ;
      RECT  5.515 1.23 7.72 1.35 ;
      RECT  7.6 1.35 7.72 1.45 ;
      RECT  5.515 1.35 5.665 1.465 ;
      RECT  3.44 1.38 3.56 1.465 ;
      RECT  3.44 1.465 5.665 1.595 ;
      RECT  4.975 1.595 5.665 1.615 ;
  END
END SEN_OAI21B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI221_0P5
#      Description : "Two 2-input ORs into 3-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI221_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI221_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.585 0.91 ;
      RECT  0.35 0.91 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.705 0.71 0.85 1.15 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.91 ;
      RECT  1.15 0.91 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.105 1.44 1.235 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.325 0.05 0.455 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.61 0.2 1.73 0.45 ;
      RECT  1.35 0.45 1.73 0.54 ;
      RECT  1.35 0.54 1.45 1.26 ;
      RECT  0.755 1.26 1.45 1.31 ;
      RECT  0.55 1.31 1.45 1.35 ;
      RECT  1.35 1.35 1.45 1.36 ;
      RECT  0.55 1.35 0.855 1.49 ;
      RECT  1.35 1.36 1.49 1.54 ;
    END
    ANTENNADIFFAREA 0.146 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.85 0.14 1.47 0.23 ;
      RECT  1.35 0.23 1.47 0.36 ;
      RECT  0.85 0.23 0.97 0.385 ;
      RECT  0.07 0.21 0.19 0.475 ;
      RECT  0.07 0.475 1.24 0.565 ;
      RECT  0.59 0.21 0.71 0.475 ;
      RECT  1.12 0.32 1.24 0.475 ;
  END
END SEN_OAI221_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI221_1
#      Description : "Two 2-input ORs into 3-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI221_1
  CLASS CORE ;
  FOREIGN SEN_OAI221_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.575 0.89 ;
      RECT  0.35 0.89 0.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.665 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.5 1.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.195 1.585 1.365 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.5 1.46 1.405 ;
      RECT  0.54 1.405 1.65 1.495 ;
      RECT  1.55 1.495 1.65 1.63 ;
    END
    ANTENNADIFFAREA 0.299 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.615 0.18 1.735 0.27 ;
      RECT  0.79 0.27 1.735 0.39 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 1.25 0.59 ;
  END
END SEN_OAI221_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI221_2
#      Description : "Two 2-input ORs into 3-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI221_2
  CLASS CORE ;
  FOREIGN SEN_OAI221_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 2.65 0.71 ;
      RECT  2.15 0.71 2.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.405 0.45 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  2.16 1.415 2.29 1.75 ;
      RECT  2.67 1.4 2.8 1.75 ;
      RECT  3.2 1.21 3.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  0.895 0.05 1.025 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.47 3.11 0.59 ;
      RECT  2.75 0.59 2.85 1.01 ;
      RECT  1.75 1.01 2.85 1.115 ;
      RECT  1.75 1.115 1.85 1.21 ;
      RECT  2.75 1.115 2.85 1.21 ;
      RECT  0.795 1.21 1.85 1.33 ;
      RECT  2.75 1.21 3.05 1.3 ;
      RECT  2.95 1.3 3.05 1.49 ;
    END
    ANTENNADIFFAREA 0.456 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.1 0.17 2.705 0.2 ;
      RECT  1.45 0.2 2.705 0.225 ;
      RECT  1.45 0.225 3.32 0.285 ;
      RECT  1.45 0.285 2.245 0.315 ;
      RECT  2.595 0.285 3.32 0.34 ;
      RECT  3.2 0.34 3.32 0.45 ;
      RECT  0.065 0.37 0.185 0.47 ;
      RECT  0.065 0.47 2.46 0.59 ;
      RECT  2.345 0.375 2.46 0.47 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.585 1.3 0.705 1.465 ;
      RECT  0.585 1.465 1.25 1.585 ;
      RECT  1.95 1.205 2.6 1.325 ;
      RECT  1.95 1.325 2.05 1.465 ;
      RECT  1.36 1.465 2.05 1.585 ;
  END
END SEN_OAI221_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI221_4
#      Description : "Two 2-input ORs into 3-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI221_4
  CLASS CORE ;
  FOREIGN SEN_OAI221_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  2.75 0.89 2.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.5 4.85 0.71 ;
      RECT  3.95 0.71 4.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.85 0.89 ;
      RECT  5.75 0.89 5.85 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.0 1.85 ;
      RECT  0.58 1.415 0.71 1.75 ;
      RECT  1.1 1.415 1.23 1.75 ;
      RECT  3.695 1.48 3.865 1.75 ;
      RECT  4.215 1.48 4.385 1.75 ;
      RECT  4.755 1.41 4.885 1.75 ;
      RECT  5.275 1.41 5.405 1.75 ;
      RECT  5.795 1.41 5.925 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      RECT  0.35 0.05 0.48 0.37 ;
      RECT  0.925 0.05 1.055 0.37 ;
      RECT  1.485 0.05 1.615 0.37 ;
      RECT  2.045 0.05 2.175 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.465 5.68 0.585 ;
      RECT  4.95 0.585 5.05 1.075 ;
      RECT  3.15 1.075 5.05 1.11 ;
      RECT  3.15 1.11 5.65 1.195 ;
      RECT  3.15 1.195 3.25 1.205 ;
      RECT  4.95 1.195 5.65 1.29 ;
      RECT  2.41 1.205 3.25 1.325 ;
      RECT  2.41 1.325 2.53 1.44 ;
      RECT  1.33 1.44 2.53 1.56 ;
    END
    ANTENNADIFFAREA 0.993 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.54 0.22 5.93 0.34 ;
      RECT  0.065 0.36 0.185 0.46 ;
      RECT  0.065 0.46 4.61 0.58 ;
      RECT  0.285 1.205 2.32 1.325 ;
      RECT  3.46 1.285 4.665 1.39 ;
      RECT  3.46 1.39 3.56 1.48 ;
      RECT  2.62 1.48 3.56 1.6 ;
  END
END SEN_OAI221_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI222_1
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&(C1|C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI222_1
  CLASS CORE ;
  FOREIGN SEN_OAI222_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.5 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.55 0.89 1.65 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.14 1.405 1.27 1.75 ;
      RECT  1.975 1.41 2.105 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.325 0.05 0.455 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.44 1.86 0.56 ;
      RECT  1.35 0.56 1.45 1.21 ;
      RECT  0.95 1.21 1.61 1.315 ;
      RECT  0.95 1.315 1.05 1.41 ;
      RECT  0.6 1.41 1.05 1.53 ;
    END
    ANTENNADIFFAREA 0.315 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.8 0.23 2.13 0.35 ;
      RECT  0.07 0.37 0.19 0.47 ;
      RECT  0.07 0.47 1.255 0.59 ;
  END
END SEN_OAI222_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI222_2
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&(C1|C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI222_2
  CLASS CORE ;
  FOREIGN SEN_OAI222_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.5 1.45 0.71 ;
      RECT  1.35 0.71 1.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.68 2.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.51 3.85 0.71 ;
      RECT  3.33 0.71 3.85 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  1.62 1.445 1.75 1.75 ;
      RECT  3.48 1.41 3.61 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.91 0.05 1.08 0.21 ;
      RECT  0.32 0.05 0.45 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.475 3.65 0.595 ;
      RECT  2.95 0.595 3.09 1.21 ;
      RECT  1.14 1.045 2.26 1.145 ;
      RECT  1.14 1.145 1.24 1.21 ;
      RECT  2.145 1.145 2.26 1.21 ;
      RECT  0.795 1.21 1.24 1.33 ;
      RECT  2.145 1.21 3.09 1.31 ;
    END
    ANTENNADIFFAREA 0.552 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.32 0.23 2.58 0.3 ;
      RECT  0.585 0.3 2.58 0.35 ;
      RECT  0.585 0.35 1.44 0.41 ;
      RECT  0.585 0.41 0.705 0.49 ;
      RECT  0.065 0.37 0.185 0.49 ;
      RECT  0.065 0.49 0.705 0.59 ;
      RECT  2.725 0.22 3.93 0.34 ;
      RECT  2.725 0.34 2.845 0.47 ;
      RECT  1.57 0.47 2.845 0.59 ;
      RECT  3.2 1.21 3.885 1.3 ;
      RECT  3.765 1.3 3.885 1.43 ;
      RECT  3.2 1.3 3.33 1.45 ;
      RECT  2.66 1.45 3.33 1.57 ;
      RECT  0.065 1.21 0.705 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  0.585 1.32 0.705 1.45 ;
      RECT  0.585 1.45 1.28 1.57 ;
      RECT  1.33 1.235 2.005 1.355 ;
      RECT  1.885 1.355 2.005 1.45 ;
      RECT  1.885 1.45 2.55 1.57 ;
  END
END SEN_OAI222_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI222_4
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&(C1|C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI222_4
  CLASS CORE ;
  FOREIGN SEN_OAI222_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.7 1.85 0.9 ;
      RECT  1.35 0.9 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.7 0.85 0.9 ;
      RECT  0.35 0.9 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.7 3.45 0.9 ;
      RECT  2.95 0.9 3.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.5 4.65 0.71 ;
      RECT  3.75 0.71 4.65 0.9 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.7 5.25 0.9 ;
      RECT  5.15 0.9 5.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.7 6.65 0.9 ;
      RECT  6.15 0.9 6.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.42 0.445 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.845 1.42 0.965 1.75 ;
      RECT  3.68 1.47 3.85 1.75 ;
      RECT  4.2 1.47 4.37 1.75 ;
      RECT  6.01 1.42 6.18 1.75 ;
      RECT  6.53 1.42 6.7 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  0.585 0.05 0.705 0.375 ;
      RECT  1.105 0.05 1.225 0.375 ;
      RECT  1.62 0.05 1.745 0.38 ;
      RECT  2.145 0.05 2.265 0.38 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.825 0.47 6.71 0.59 ;
      RECT  5.55 0.59 5.66 1.21 ;
      RECT  3.15 1.06 4.85 1.17 ;
      RECT  4.75 1.17 4.85 1.21 ;
      RECT  3.15 1.17 3.305 1.22 ;
      RECT  4.75 1.21 5.66 1.33 ;
      RECT  1.95 1.09 2.85 1.215 ;
      RECT  1.325 1.215 2.85 1.22 ;
      RECT  1.325 1.22 3.305 1.29 ;
      RECT  2.755 1.29 3.305 1.33 ;
      RECT  1.325 1.29 2.05 1.335 ;
    END
    ANTENNADIFFAREA 1.112 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.64 0.215 5.81 0.23 ;
      RECT  2.355 0.23 6.935 0.35 ;
      RECT  6.815 0.35 6.935 0.455 ;
      RECT  0.325 0.38 0.445 0.47 ;
      RECT  0.325 0.47 4.46 0.59 ;
      RECT  4.355 0.445 4.46 0.47 ;
      RECT  4.355 0.59 4.46 0.615 ;
      RECT  0.06 1.21 1.23 1.33 ;
      RECT  0.06 1.33 0.19 1.435 ;
      RECT  1.1 1.33 1.23 1.465 ;
      RECT  1.1 1.465 2.26 1.585 ;
      RECT  2.14 1.385 2.26 1.465 ;
      RECT  5.77 1.21 6.94 1.33 ;
      RECT  6.81 1.33 6.94 1.415 ;
      RECT  5.77 1.33 5.9 1.45 ;
      RECT  4.695 1.45 5.9 1.57 ;
      RECT  3.445 1.26 4.605 1.38 ;
      RECT  3.445 1.38 3.57 1.48 ;
      RECT  4.485 1.38 4.605 1.515 ;
      RECT  2.405 1.395 2.525 1.48 ;
      RECT  2.405 1.48 3.57 1.6 ;
  END
END SEN_OAI222_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI222_0P5
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&(C1|C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI222_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI222_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.91 ;
      RECT  0.35 0.91 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.91 ;
      RECT  1.14 0.91 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.12 1.44 1.25 1.75 ;
      RECT  1.94 1.41 2.07 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.325 0.05 0.445 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.645 0.32 1.765 0.51 ;
      RECT  1.645 0.51 1.85 0.6 ;
      RECT  1.75 0.6 1.85 1.455 ;
      RECT  0.55 1.26 1.45 1.35 ;
      RECT  1.35 1.35 1.45 1.455 ;
      RECT  0.55 1.35 0.85 1.49 ;
      RECT  1.35 1.455 1.85 1.575 ;
    END
    ANTENNADIFFAREA 0.166 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.14 1.245 0.23 ;
      RECT  1.125 0.23 1.245 0.39 ;
      RECT  0.585 0.23 0.705 0.455 ;
      RECT  0.065 0.21 0.185 0.455 ;
      RECT  0.065 0.455 0.705 0.545 ;
      RECT  1.375 0.14 2.035 0.23 ;
      RECT  1.915 0.23 2.035 0.4 ;
      RECT  1.375 0.23 1.495 0.51 ;
      RECT  0.805 0.32 1.025 0.44 ;
      RECT  0.935 0.44 1.025 0.51 ;
      RECT  0.935 0.51 1.495 0.6 ;
  END
END SEN_OAI222_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI222_0P75
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&(C1|C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI222_0P75
  CLASS CORE ;
  FOREIGN SEN_OAI222_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.905 ;
      RECT  0.35 0.905 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.695 0.85 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.25 0.905 ;
      RECT  1.15 0.905 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.51 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.12 1.415 1.25 1.75 ;
      RECT  1.94 1.21 2.06 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.645 0.32 1.765 0.51 ;
      RECT  1.645 0.51 1.85 0.6 ;
      RECT  1.75 0.6 1.85 1.455 ;
      RECT  0.535 1.205 1.45 1.325 ;
      RECT  1.35 1.325 1.45 1.455 ;
      RECT  1.35 1.455 1.85 1.575 ;
    END
    ANTENNADIFFAREA 0.239 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.375 0.14 2.035 0.23 ;
      RECT  1.915 0.23 2.035 0.405 ;
      RECT  1.375 0.23 1.495 0.42 ;
      RECT  0.805 0.42 1.495 0.535 ;
      RECT  0.585 0.215 1.285 0.33 ;
      RECT  0.585 0.33 0.705 0.475 ;
      RECT  0.065 0.345 0.185 0.475 ;
      RECT  0.065 0.475 0.705 0.565 ;
  END
END SEN_OAI222_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI222_3
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2)&(C1|C2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI222_3
  CLASS CORE ;
  FOREIGN SEN_OAI222_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.25 0.9 ;
      RECT  1.55 0.9 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.45 0.9 ;
      RECT  3.35 0.9 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B2
  PIN C1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END C1
  PIN C2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 5.05 0.89 ;
      RECT  4.95 0.89 5.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 5.2 1.85 ;
      RECT  0.58 1.415 0.71 1.75 ;
      RECT  2.66 1.42 2.79 1.75 ;
      RECT  3.18 1.42 3.31 1.75 ;
      RECT  4.485 1.415 4.615 1.75 ;
      RECT  5.01 1.21 5.13 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.45 4.92 0.57 ;
      RECT  3.55 0.57 3.65 1.21 ;
      RECT  1.055 1.21 4.14 1.33 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.835 0.24 5.13 0.36 ;
      RECT  5.01 0.36 5.13 0.46 ;
      RECT  0.065 0.375 0.185 0.475 ;
      RECT  0.065 0.475 3.37 0.595 ;
      RECT  1.835 1.0 3.095 1.12 ;
      RECT  0.275 1.205 0.965 1.325 ;
      RECT  0.845 1.325 0.965 1.44 ;
      RECT  0.845 1.44 1.535 1.56 ;
      RECT  4.285 1.205 4.92 1.325 ;
      RECT  4.285 1.325 4.375 1.44 ;
      RECT  3.66 1.44 4.375 1.56 ;
  END
END SEN_OAI222_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_0P5
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI22_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.5 1.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.15 1.41 1.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.32 0.05 0.45 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.815 0.32 1.05 0.45 ;
      RECT  0.95 0.45 1.05 1.42 ;
      RECT  0.54 1.42 1.05 1.54 ;
    END
    ANTENNADIFFAREA 0.118 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.14 1.265 0.23 ;
      RECT  1.145 0.23 1.265 0.39 ;
      RECT  0.585 0.23 0.705 0.47 ;
      RECT  0.065 0.22 0.185 0.47 ;
      RECT  0.065 0.47 0.705 0.56 ;
  END
END SEN_OAI22_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_1
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_1
  CLASS CORE ;
  FOREIGN SEN_OAI22_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.5 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.085 1.41 0.215 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.195 1.41 1.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.36 0.05 0.52 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.45 1.05 1.44 ;
      RECT  0.62 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.226 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.67 0.17 1.32 0.26 ;
      RECT  1.2 0.26 1.32 0.39 ;
      RECT  0.67 0.26 0.79 0.48 ;
      RECT  0.075 0.48 0.79 0.59 ;
  END
END SEN_OAI22_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_2
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_2
  CLASS CORE ;
  FOREIGN SEN_OAI22_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 0.71 ;
      RECT  1.35 0.71 1.66 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.71 ;
      RECT  1.95 0.71 2.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.9 ;
      RECT  0.75 0.9 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  2.135 1.41 2.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.32 0.05 0.45 0.37 ;
      RECT  0.84 0.05 0.97 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.56 0.41 2.255 0.54 ;
      RECT  2.135 0.54 2.255 0.59 ;
      RECT  1.75 0.54 1.85 1.22 ;
      RECT  0.82 1.22 1.85 1.34 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.13 0.2 2.525 0.32 ;
      RECT  2.39 0.32 2.525 0.39 ;
      RECT  1.13 0.32 1.25 0.47 ;
      RECT  0.065 0.37 0.185 0.47 ;
      RECT  0.065 0.47 1.25 0.59 ;
      RECT  1.955 1.21 2.515 1.3 ;
      RECT  2.395 1.3 2.515 1.43 ;
      RECT  1.955 1.3 2.045 1.48 ;
      RECT  1.355 1.43 1.475 1.48 ;
      RECT  1.355 1.48 2.045 1.6 ;
      RECT  0.065 1.21 0.705 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  0.585 1.32 0.705 1.48 ;
      RECT  0.585 1.48 1.225 1.6 ;
      RECT  1.105 1.43 1.225 1.48 ;
  END
END SEN_OAI22_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_3
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_3
  CLASS CORE ;
  FOREIGN SEN_OAI22_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.715 0.71 2.06 0.89 ;
      RECT  1.715 0.89 1.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 3.25 0.71 ;
      RECT  2.55 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  2.66 1.41 2.79 1.75 ;
      RECT  3.195 1.21 3.315 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.835 0.45 3.045 0.57 ;
      RECT  2.925 0.57 3.045 0.62 ;
      RECT  2.15 0.57 2.25 1.21 ;
      RECT  1.075 1.21 2.29 1.33 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.625 0.24 3.305 0.36 ;
      RECT  3.185 0.36 3.305 0.41 ;
      RECT  1.625 0.36 1.745 0.48 ;
      RECT  0.065 0.37 0.185 0.48 ;
      RECT  0.065 0.48 1.745 0.59 ;
      RECT  0.275 1.21 0.965 1.32 ;
      RECT  0.845 1.32 0.965 1.455 ;
      RECT  0.845 1.455 1.54 1.575 ;
      RECT  2.4 1.21 3.07 1.32 ;
      RECT  2.4 1.32 2.53 1.445 ;
      RECT  1.83 1.445 2.53 1.565 ;
  END
END SEN_OAI22_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_4
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_4
  CLASS CORE ;
  FOREIGN SEN_OAI22_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.71 ;
      RECT  2.35 0.71 3.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.745 0.7 4.25 0.9 ;
      RECT  4.15 0.9 4.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.42 0.45 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.84 1.42 0.97 1.75 ;
      RECT  3.625 1.42 3.755 1.75 ;
      RECT  4.145 1.42 4.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.32 0.05 0.45 0.38 ;
      RECT  0.84 0.05 0.97 0.38 ;
      RECT  1.36 0.05 1.49 0.38 ;
      RECT  1.88 0.05 2.01 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.54 0.42 4.32 0.54 ;
      RECT  3.35 0.54 3.455 1.01 ;
      RECT  1.95 1.01 3.455 1.12 ;
      RECT  1.95 1.12 2.05 1.22 ;
      RECT  1.315 1.22 2.05 1.34 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.145 0.2 4.53 0.32 ;
      RECT  4.41 0.32 4.53 0.39 ;
      RECT  2.145 0.32 2.26 0.47 ;
      RECT  0.065 0.37 0.19 0.47 ;
      RECT  0.065 0.47 2.26 0.59 ;
      RECT  0.065 1.21 1.225 1.33 ;
      RECT  0.065 1.33 0.185 1.43 ;
      RECT  1.105 1.33 1.225 1.48 ;
      RECT  1.105 1.48 2.265 1.6 ;
      RECT  2.145 1.42 2.265 1.48 ;
      RECT  2.28 1.21 4.53 1.33 ;
      RECT  4.41 1.33 4.53 1.43 ;
  END
END SEN_OAI22_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_12
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_12
  CLASS CORE ;
  FOREIGN SEN_OAI22_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.775 0.71 12.175 0.9 ;
      RECT  10.875 0.71 11.175 0.9 ;
      RECT  9.78 0.71 10.05 0.9 ;
      RECT  8.915 0.71 9.225 0.9 ;
      RECT  7.855 0.71 8.155 0.9 ;
      RECT  6.95 0.71 7.34 0.9 ;
      LAYER M2 ;
      RECT  7.0 0.75 12.115 0.85 ;
      LAYER V1 ;
      RECT  11.775 0.75 11.875 0.85 ;
      RECT  11.975 0.75 12.075 0.85 ;
      RECT  11.015 0.75 11.115 0.85 ;
      RECT  9.845 0.75 9.945 0.85 ;
      RECT  8.99 0.75 9.09 0.85 ;
      RECT  7.855 0.75 7.955 0.85 ;
      RECT  8.055 0.75 8.155 0.85 ;
      RECT  7.04 0.75 7.14 0.85 ;
      RECT  7.24 0.75 7.34 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  12.45 0.75 12.545 0.89 ;
      RECT  12.36 0.89 12.545 1.09 ;
      RECT  11.415 0.71 11.505 0.91 ;
      RECT  11.34 0.91 11.505 1.09 ;
      RECT  10.375 0.775 10.615 0.895 ;
      RECT  10.375 0.895 10.475 1.09 ;
      RECT  9.455 0.715 9.635 0.845 ;
      RECT  9.455 0.845 9.555 1.09 ;
      RECT  8.425 0.715 8.525 0.93 ;
      RECT  8.425 0.93 8.68 1.09 ;
      RECT  7.43 0.755 7.52 0.91 ;
      RECT  7.43 0.91 7.73 1.09 ;
      RECT  6.475 0.71 6.66 1.09 ;
      LAYER M2 ;
      RECT  6.52 0.95 12.56 1.05 ;
      LAYER V1 ;
      RECT  12.42 0.95 12.52 1.05 ;
      RECT  11.405 0.95 11.505 1.05 ;
      RECT  10.375 0.95 10.475 1.05 ;
      RECT  9.455 0.95 9.555 1.05 ;
      RECT  8.425 0.95 8.525 1.05 ;
      RECT  7.43 0.95 7.53 1.05 ;
      RECT  7.63 0.95 7.73 1.05 ;
      RECT  6.56 0.95 6.66 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.525 0.71 5.905 0.885 ;
      RECT  4.74 0.71 5.04 0.9 ;
      RECT  3.71 0.71 4.01 0.9 ;
      RECT  2.695 0.71 2.995 0.9 ;
      RECT  1.605 0.71 1.895 0.9 ;
      RECT  0.625 0.71 0.965 0.9 ;
      LAYER M2 ;
      RECT  0.62 0.75 6.09 0.85 ;
      LAYER V1 ;
      RECT  5.765 0.75 5.865 0.85 ;
      RECT  4.83 0.75 4.93 0.85 ;
      RECT  3.745 0.75 3.845 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.64 0.75 1.74 0.85 ;
      RECT  0.66 0.75 0.76 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.215 0.755 6.305 0.91 ;
      RECT  5.995 0.91 6.305 1.09 ;
      RECT  5.285 0.715 5.385 0.93 ;
      RECT  5.19 0.93 5.385 1.09 ;
      RECT  4.255 0.715 4.345 0.91 ;
      RECT  4.255 0.91 4.445 1.09 ;
      RECT  3.155 0.715 3.245 0.91 ;
      RECT  3.155 0.91 3.36 1.09 ;
      RECT  2.155 0.715 2.245 0.91 ;
      RECT  2.155 0.91 2.33 1.09 ;
      RECT  1.15 0.715 1.25 0.91 ;
      RECT  1.15 0.91 1.375 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.43 1.09 ;
      LAYER M2 ;
      RECT  0.17 0.95 6.135 1.05 ;
      LAYER V1 ;
      RECT  5.995 0.95 6.095 1.05 ;
      RECT  5.285 0.95 5.385 1.05 ;
      RECT  4.305 0.95 4.405 1.05 ;
      RECT  3.185 0.95 3.285 1.05 ;
      RECT  2.155 0.95 2.255 1.05 ;
      RECT  1.15 0.95 1.25 1.05 ;
      RECT  0.21 0.95 0.31 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  3.18 1.44 3.31 1.75 ;
      RECT  4.22 1.44 4.35 1.75 ;
      RECT  5.26 1.44 5.39 1.75 ;
      RECT  6.3 1.44 6.43 1.75 ;
      RECT  7.34 1.44 7.47 1.75 ;
      RECT  8.38 1.44 8.51 1.75 ;
      RECT  9.42 1.44 9.55 1.75 ;
      RECT  10.46 1.44 10.59 1.75 ;
      RECT  11.5 1.44 11.63 1.75 ;
      RECT  12.565 1.21 12.685 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      RECT  0.845 0.05 0.97 0.36 ;
      RECT  1.36 0.05 1.49 0.36 ;
      RECT  1.88 0.05 2.01 0.36 ;
      RECT  2.4 0.05 2.53 0.36 ;
      RECT  2.92 0.05 3.05 0.36 ;
      RECT  3.44 0.05 3.57 0.36 ;
      RECT  3.96 0.05 4.09 0.36 ;
      RECT  4.48 0.05 4.61 0.36 ;
      RECT  5.0 0.05 5.13 0.36 ;
      RECT  5.52 0.05 5.65 0.36 ;
      RECT  6.04 0.05 6.165 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.12 0.5 12.455 0.62 ;
      RECT  10.15 0.62 10.25 1.11 ;
      RECT  11.595 0.62 11.685 1.11 ;
      RECT  9.75 1.11 10.25 1.18 ;
      RECT  11.595 1.11 12.25 1.18 ;
      RECT  7.555 0.5 8.815 0.62 ;
      RECT  8.245 0.62 8.335 1.11 ;
      RECT  7.865 1.11 8.335 1.18 ;
      RECT  6.53 0.5 7.255 0.62 ;
      RECT  6.75 0.62 6.86 1.11 ;
      RECT  6.75 1.11 7.25 1.18 ;
      RECT  0.55 1.11 1.05 1.18 ;
      RECT  0.55 1.18 12.25 1.35 ;
      RECT  1.55 1.11 2.05 1.18 ;
      RECT  2.55 1.11 3.05 1.18 ;
      RECT  3.55 1.11 4.05 1.18 ;
      RECT  4.55 1.11 5.05 1.18 ;
      RECT  5.55 1.11 5.89 1.18 ;
      RECT  8.905 1.11 9.255 1.18 ;
      RECT  10.75 1.11 11.25 1.18 ;
    END
    ANTENNADIFFAREA 2.592 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.27 0.19 12.665 0.36 ;
      RECT  6.27 0.36 6.44 0.45 ;
      RECT  7.35 0.36 7.45 0.49 ;
      RECT  8.93 0.36 9.03 0.49 ;
      RECT  1.625 0.31 1.725 0.45 ;
      RECT  0.065 0.45 6.44 0.62 ;
      RECT  2.15 0.31 2.25 0.45 ;
      RECT  2.685 0.31 2.785 0.45 ;
      RECT  3.2 0.31 3.3 0.45 ;
      RECT  3.725 0.31 3.825 0.45 ;
      RECT  4.22 0.31 4.32 0.45 ;
      RECT  4.75 0.31 4.85 0.45 ;
      RECT  5.25 0.31 5.35 0.45 ;
      RECT  5.78 0.31 5.88 0.45 ;
      LAYER M2 ;
      RECT  1.58 0.35 9.07 0.45 ;
      LAYER V1 ;
      RECT  1.625 0.35 1.725 0.45 ;
      RECT  2.15 0.35 2.25 0.45 ;
      RECT  2.685 0.35 2.785 0.45 ;
      RECT  3.2 0.35 3.3 0.45 ;
      RECT  3.725 0.35 3.825 0.45 ;
      RECT  4.22 0.35 4.32 0.45 ;
      RECT  4.75 0.35 4.85 0.45 ;
      RECT  5.25 0.35 5.35 0.45 ;
      RECT  5.78 0.35 5.88 0.45 ;
      RECT  7.35 0.35 7.45 0.45 ;
      RECT  8.93 0.35 9.03 0.45 ;
  END
END SEN_OAI22_12
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_6
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_6
  CLASS CORE ;
  FOREIGN SEN_OAI22_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.71 6.05 0.89 ;
      RECT  4.75 0.71 5.05 0.89 ;
      RECT  3.75 0.71 4.05 0.89 ;
      LAYER M2 ;
      RECT  3.71 0.75 6.09 0.85 ;
      LAYER V1 ;
      RECT  5.75 0.75 5.85 0.85 ;
      RECT  5.95 0.75 6.05 0.85 ;
      RECT  4.75 0.75 4.85 0.85 ;
      RECT  4.95 0.75 5.05 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  3.95 0.75 4.05 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.45 0.89 ;
      RECT  6.15 0.89 6.25 1.09 ;
      RECT  5.35 0.71 5.45 0.91 ;
      RECT  5.15 0.91 5.45 1.09 ;
      RECT  4.35 0.71 4.45 0.91 ;
      RECT  4.35 0.91 4.65 1.09 ;
      RECT  3.35 0.695 3.45 1.115 ;
      LAYER M2 ;
      RECT  3.31 0.95 6.29 1.05 ;
      LAYER V1 ;
      RECT  6.15 0.95 6.25 1.05 ;
      RECT  5.15 0.95 5.25 1.05 ;
      RECT  5.35 0.95 5.45 1.05 ;
      RECT  4.35 0.95 4.45 1.05 ;
      RECT  4.55 0.95 4.65 1.05 ;
      RECT  3.35 0.95 3.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 2.85 0.89 ;
      RECT  1.55 0.71 1.85 0.9 ;
      RECT  0.55 0.71 0.85 0.89 ;
      LAYER M2 ;
      RECT  0.51 0.75 2.89 0.85 ;
      LAYER V1 ;
      RECT  2.55 0.75 2.65 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  1.55 0.75 1.65 0.85 ;
      RECT  1.75 0.75 1.85 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
      RECT  0.75 0.75 0.85 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.25 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
      RECT  2.15 0.71 2.25 0.91 ;
      RECT  2.15 0.91 2.45 1.09 ;
      RECT  1.155 0.71 1.245 0.91 ;
      RECT  1.155 0.91 1.455 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.45 1.09 ;
      LAYER M2 ;
      RECT  0.11 0.95 3.09 1.05 ;
      LAYER V1 ;
      RECT  2.95 0.95 3.05 1.05 ;
      RECT  2.15 0.95 2.25 1.05 ;
      RECT  2.35 0.95 2.45 1.05 ;
      RECT  1.155 0.95 1.255 1.05 ;
      RECT  1.355 0.95 1.455 1.05 ;
      RECT  0.15 0.95 0.25 1.05 ;
      RECT  0.35 0.95 0.45 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3888 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  1.1 1.425 1.23 1.75 ;
      RECT  2.14 1.425 2.27 1.75 ;
      RECT  3.18 1.425 3.31 1.75 ;
      RECT  4.24 1.425 4.37 1.75 ;
      RECT  5.28 1.425 5.41 1.75 ;
      RECT  6.36 1.21 6.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.84 0.05 0.97 0.39 ;
      RECT  1.36 0.05 1.49 0.39 ;
      RECT  1.88 0.05 2.01 0.39 ;
      RECT  2.4 0.05 2.53 0.39 ;
      RECT  2.92 0.05 3.05 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.44 0.45 6.24 0.58 ;
      RECT  3.54 0.58 3.66 1.205 ;
      RECT  5.54 0.58 5.66 1.205 ;
      RECT  0.535 1.205 5.975 1.335 ;
    END
    ANTENNADIFFAREA 1.314 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.18 0.215 6.51 0.345 ;
      RECT  3.18 0.345 3.31 0.48 ;
      RECT  0.065 0.39 0.185 0.48 ;
      RECT  0.065 0.48 3.31 0.61 ;
  END
END SEN_OAI22_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_8
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_8
  CLASS CORE ;
  FOREIGN SEN_OAI22_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.77 0.71 8.07 0.9 ;
      RECT  6.74 0.71 7.105 0.895 ;
      RECT  5.815 0.71 6.115 0.9 ;
      RECT  4.795 0.71 5.115 0.9 ;
      LAYER M2 ;
      RECT  4.775 0.75 8.11 0.85 ;
      LAYER V1 ;
      RECT  7.77 0.75 7.87 0.85 ;
      RECT  7.97 0.75 8.07 0.85 ;
      RECT  6.815 0.75 6.915 0.85 ;
      RECT  5.905 0.75 6.005 0.85 ;
      RECT  4.815 0.75 4.915 0.85 ;
      RECT  5.015 0.75 5.115 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.16 0.755 8.335 0.91 ;
      RECT  8.16 0.91 8.395 1.09 ;
      RECT  7.38 0.72 7.48 0.91 ;
      RECT  7.38 0.91 7.68 1.09 ;
      RECT  6.35 0.72 6.45 0.91 ;
      RECT  6.35 0.91 6.65 1.09 ;
      RECT  5.385 0.715 5.485 0.91 ;
      RECT  5.385 0.91 5.575 1.09 ;
      RECT  4.395 0.755 4.485 0.91 ;
      RECT  4.395 0.91 4.635 1.09 ;
      LAYER M2 ;
      RECT  4.385 0.95 8.34 1.05 ;
      LAYER V1 ;
      RECT  8.16 0.95 8.26 1.05 ;
      RECT  7.38 0.95 7.48 1.05 ;
      RECT  7.58 0.95 7.68 1.05 ;
      RECT  6.35 0.95 6.45 1.05 ;
      RECT  6.55 0.95 6.65 1.05 ;
      RECT  5.385 0.95 5.485 1.05 ;
      RECT  4.425 0.95 4.525 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.56 0.71 3.86 0.9 ;
      RECT  2.665 0.71 2.965 0.9 ;
      RECT  1.64 0.71 1.94 0.9 ;
      RECT  0.575 0.71 0.915 0.9 ;
      LAYER M2 ;
      RECT  0.735 0.75 4.09 0.85 ;
      LAYER V1 ;
      RECT  3.56 0.75 3.66 0.85 ;
      RECT  3.76 0.75 3.86 0.85 ;
      RECT  2.71 0.75 2.81 0.85 ;
      RECT  1.745 0.75 1.845 0.85 ;
      RECT  0.775 0.75 0.875 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.135 0.755 4.265 0.91 ;
      RECT  3.95 0.91 4.265 1.09 ;
      RECT  3.165 0.715 3.255 0.91 ;
      RECT  3.165 0.91 3.315 1.09 ;
      RECT  2.155 0.715 2.245 0.91 ;
      RECT  2.155 0.91 2.33 1.09 ;
      RECT  1.155 0.715 1.245 0.91 ;
      RECT  1.155 0.91 1.365 1.09 ;
      RECT  0.15 0.71 0.25 0.91 ;
      RECT  0.15 0.91 0.35 1.09 ;
      LAYER M2 ;
      RECT  0.17 0.95 4.09 1.05 ;
      LAYER V1 ;
      RECT  3.95 0.95 4.05 1.05 ;
      RECT  3.165 0.95 3.265 1.05 ;
      RECT  2.16 0.95 2.26 1.05 ;
      RECT  1.155 0.95 1.255 1.05 ;
      RECT  0.21 0.95 0.31 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  1.105 1.44 1.225 1.75 ;
      RECT  2.145 1.44 2.265 1.75 ;
      RECT  3.185 1.44 3.305 1.75 ;
      RECT  4.225 1.44 4.345 1.75 ;
      RECT  5.265 1.44 5.385 1.75 ;
      RECT  6.305 1.44 6.425 1.75 ;
      RECT  7.345 1.44 7.465 1.75 ;
      RECT  8.4 1.21 8.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  0.325 0.05 0.445 0.36 ;
      RECT  0.845 0.05 0.965 0.36 ;
      RECT  1.365 0.05 1.485 0.36 ;
      RECT  1.885 0.05 2.005 0.36 ;
      RECT  2.405 0.05 2.525 0.36 ;
      RECT  2.925 0.05 3.045 0.36 ;
      RECT  3.445 0.05 3.565 0.36 ;
      RECT  3.965 0.05 4.085 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.445 0.465 8.295 0.585 ;
      RECT  5.205 0.585 5.295 1.11 ;
      RECT  7.2 0.585 7.29 1.11 ;
      RECT  4.75 1.11 5.295 1.18 ;
      RECT  6.75 1.11 7.29 1.18 ;
      RECT  0.55 1.11 1.05 1.18 ;
      RECT  0.55 1.18 8.05 1.35 ;
      RECT  1.55 1.11 2.05 1.18 ;
      RECT  2.55 1.11 3.05 1.18 ;
      RECT  3.55 1.11 3.85 1.18 ;
      RECT  5.75 1.11 6.25 1.18 ;
      RECT  7.88 1.11 8.05 1.18 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.185 0.19 8.505 0.36 ;
      RECT  4.185 0.36 4.355 0.45 ;
      RECT  0.065 0.45 4.355 0.62 ;
  END
END SEN_OAI22_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_S_0P5
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_S_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI22_S_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0285 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.15 1.41 1.28 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.325 0.05 0.455 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.81 0.345 1.05 0.465 ;
      RECT  0.95 0.465 1.05 1.44 ;
      RECT  0.54 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.112 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.59 0.14 1.285 0.23 ;
      RECT  1.165 0.23 1.285 0.395 ;
      RECT  0.59 0.23 0.71 0.47 ;
      RECT  0.07 0.185 0.19 0.47 ;
      RECT  0.07 0.47 0.71 0.56 ;
  END
END SEN_OAI22_S_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_S_1
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_S_1
  CLASS CORE ;
  FOREIGN SEN_OAI22_S_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.68 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0561 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0561 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0561 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.68 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0561 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.15 1.21 1.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.325 0.05 0.455 0.38 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.81 0.345 1.05 0.465 ;
      RECT  0.95 0.465 1.05 1.44 ;
      RECT  0.54 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.59 0.14 1.285 0.23 ;
      RECT  1.165 0.23 1.285 0.4 ;
      RECT  0.59 0.23 0.71 0.47 ;
      RECT  0.07 0.315 0.19 0.47 ;
      RECT  0.07 0.47 0.71 0.56 ;
  END
END SEN_OAI22_S_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_S_2
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_S_2
  CLASS CORE ;
  FOREIGN SEN_OAI22_S_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1122 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.62 2.25 1.115 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1122 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.05 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1122 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1122 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  2.13 1.415 2.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.3 0.05 0.47 0.32 ;
      RECT  0.82 0.05 0.99 0.32 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.395 0.31 2.515 0.41 ;
      RECT  1.33 0.41 2.515 0.53 ;
      RECT  1.33 0.53 1.45 1.11 ;
      RECT  0.845 1.11 1.735 1.29 ;
    END
    ANTENNADIFFAREA 0.418 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.105 0.2 2.305 0.32 ;
      RECT  1.105 0.32 1.225 0.41 ;
      RECT  0.065 0.31 0.185 0.41 ;
      RECT  0.065 0.41 1.225 0.53 ;
      RECT  0.065 1.225 0.705 1.315 ;
      RECT  0.065 1.315 0.185 1.445 ;
      RECT  0.585 1.315 0.705 1.52 ;
      RECT  0.585 1.52 1.225 1.61 ;
      RECT  1.105 1.38 1.225 1.52 ;
      RECT  1.875 1.205 2.515 1.325 ;
      RECT  2.395 1.325 2.515 1.425 ;
      RECT  1.875 1.325 1.995 1.45 ;
      RECT  1.315 1.45 1.995 1.57 ;
  END
END SEN_OAI22_S_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_S_3
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_S_3
  CLASS CORE ;
  FOREIGN SEN_OAI22_S_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.05 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1683 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.71 3.05 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1683 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1683 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1683 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.07 1.21 0.19 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.59 1.215 0.71 1.75 ;
      RECT  2.665 1.45 2.795 1.75 ;
      RECT  3.21 1.21 3.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.305 0.05 0.475 0.32 ;
      RECT  0.825 0.05 0.995 0.32 ;
      RECT  1.345 0.05 1.515 0.32 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.84 0.41 3.1 0.53 ;
      RECT  2.15 0.53 2.255 1.24 ;
      RECT  1.06 1.24 2.255 1.365 ;
    END
    ANTENNADIFFAREA 0.564 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.63 0.2 3.31 0.32 ;
      RECT  1.63 0.32 1.75 0.415 ;
      RECT  3.19 0.32 3.31 0.42 ;
      RECT  0.07 0.315 0.19 0.415 ;
      RECT  0.07 0.415 1.75 0.535 ;
      RECT  0.34 1.035 0.97 1.125 ;
      RECT  0.34 1.125 0.45 1.255 ;
      RECT  0.85 1.125 0.97 1.455 ;
      RECT  0.85 1.455 1.54 1.575 ;
      RECT  2.41 1.24 3.1 1.36 ;
      RECT  2.41 1.36 2.53 1.455 ;
      RECT  1.84 1.455 2.53 1.575 ;
  END
END SEN_OAI22_S_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_S_4
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_S_4
  CLASS CORE ;
  FOREIGN SEN_OAI22_S_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.635 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2241 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2241 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.795 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2241 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2241 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.45 0.45 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.84 1.45 0.97 1.75 ;
      RECT  3.49 1.45 3.62 1.75 ;
      RECT  4.05 1.45 4.18 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.38 0.05 0.51 0.35 ;
      RECT  1.035 0.05 1.165 0.35 ;
      RECT  1.62 0.05 1.75 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.145 0.32 2.265 0.435 ;
      RECT  2.145 0.435 4.45 0.525 ;
      RECT  2.665 0.32 2.785 0.435 ;
      RECT  3.185 0.32 3.305 0.435 ;
      RECT  3.795 0.32 3.915 0.435 ;
      RECT  4.315 0.29 4.45 0.435 ;
      RECT  2.35 0.525 2.45 1.11 ;
      RECT  1.35 1.11 3.05 1.29 ;
    END
    ANTENNADIFFAREA 0.841 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.885 0.14 4.175 0.23 ;
      RECT  2.405 0.23 2.525 0.345 ;
      RECT  2.925 0.23 3.045 0.345 ;
      RECT  3.49 0.23 3.61 0.345 ;
      RECT  4.055 0.23 4.175 0.345 ;
      RECT  1.885 0.23 2.005 0.44 ;
      RECT  0.065 0.34 0.185 0.44 ;
      RECT  0.065 0.44 2.005 0.56 ;
      RECT  0.065 1.24 1.225 1.36 ;
      RECT  1.105 1.36 1.225 1.44 ;
      RECT  0.065 1.36 0.185 1.46 ;
      RECT  1.105 1.44 2.315 1.56 ;
      RECT  3.185 1.24 4.485 1.36 ;
      RECT  3.185 1.36 3.305 1.44 ;
      RECT  2.615 1.44 3.305 1.56 ;
  END
END SEN_OAI22_S_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_S_8
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_S_8
  CLASS CORE ;
  FOREIGN SEN_OAI22_S_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.615 0.67 5.85 0.89 ;
      RECT  5.75 0.89 5.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.35 0.71 7.45 0.89 ;
      RECT  7.35 0.89 7.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.66 3.65 0.89 ;
      RECT  2.55 0.89 2.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.25 0.445 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  0.845 1.25 0.965 1.75 ;
      RECT  1.365 1.25 1.485 1.75 ;
      RECT  1.885 1.25 2.005 1.75 ;
      RECT  6.055 1.42 6.185 1.75 ;
      RECT  6.61 1.405 6.74 1.75 ;
      RECT  7.17 1.405 7.3 1.75 ;
      RECT  7.71 1.405 7.84 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  0.56 0.05 0.73 0.325 ;
      RECT  1.08 0.05 1.25 0.325 ;
      RECT  1.6 0.05 1.77 0.325 ;
      RECT  2.12 0.05 2.29 0.325 ;
      RECT  2.64 0.05 2.81 0.325 ;
      RECT  3.16 0.05 3.33 0.325 ;
      RECT  3.68 0.05 3.85 0.325 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.18 0.415 7.635 0.53 ;
      RECT  4.35 0.53 7.635 0.56 ;
      RECT  4.35 0.56 4.52 1.11 ;
      RECT  2.75 1.11 5.65 1.18 ;
      RECT  2.38 1.18 5.65 1.29 ;
    END
    ANTENNADIFFAREA 1.535 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.96 0.195 7.895 0.325 ;
      RECT  3.96 0.325 4.09 0.415 ;
      RECT  0.34 0.325 0.445 0.415 ;
      RECT  0.34 0.415 4.09 0.545 ;
      RECT  1.585 1.01 2.29 1.04 ;
      RECT  0.065 1.04 2.29 1.16 ;
      RECT  0.065 1.16 0.185 1.26 ;
      RECT  2.12 1.16 2.29 1.44 ;
      RECT  2.12 1.44 3.875 1.56 ;
      RECT  2.12 1.56 2.825 1.59 ;
      RECT  5.76 1.18 8.155 1.3 ;
      RECT  5.76 1.3 6.5 1.33 ;
      RECT  5.76 1.33 5.93 1.41 ;
      RECT  5.225 1.41 5.93 1.44 ;
      RECT  4.175 1.44 5.93 1.56 ;
  END
END SEN_OAI22_S_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_0P75
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_0P75
  CLASS CORE ;
  FOREIGN SEN_OAI22_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.905 ;
      RECT  0.35 0.905 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.14 1.21 1.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.32 0.05 0.45 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.795 0.41 1.05 0.53 ;
      RECT  0.95 0.53 1.05 1.45 ;
      RECT  0.535 1.45 1.05 1.57 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.2 1.295 0.32 ;
      RECT  0.585 0.32 0.705 0.45 ;
      RECT  0.065 0.32 0.185 0.45 ;
      RECT  0.065 0.45 0.705 0.54 ;
  END
END SEN_OAI22_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_T_0P5
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_T_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI22_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.645 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0504 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 0.65 0.91 ;
      RECT  0.35 0.91 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0468 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.14 1.21 1.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.795 0.32 1.05 0.44 ;
      RECT  0.95 0.44 1.05 1.44 ;
      RECT  0.535 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.108 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.585 0.14 1.26 0.23 ;
      RECT  1.14 0.23 1.26 0.41 ;
      RECT  0.585 0.23 0.705 0.475 ;
      RECT  0.065 0.345 0.185 0.475 ;
      RECT  0.065 0.475 0.705 0.565 ;
  END
END SEN_OAI22_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_T_1
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_T_1
  CLASS CORE ;
  FOREIGN SEN_OAI22_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.65 0.815 ;
      RECT  1.15 0.815 1.65 0.915 ;
      RECT  1.15 0.915 1.25 1.09 ;
      RECT  1.55 0.915 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1008 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0936 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.24 1.21 0.36 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.545 1.415 1.675 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.325 0.05 0.455 0.365 ;
      RECT  0.845 0.05 0.975 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.345 0.44 1.54 0.56 ;
      RECT  1.345 0.56 1.455 0.635 ;
      RECT  0.94 0.635 1.455 0.725 ;
      RECT  0.94 0.725 1.06 1.29 ;
    END
    ANTENNADIFFAREA 0.324 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.11 0.23 1.8 0.35 ;
      RECT  1.11 0.35 1.23 0.455 ;
      RECT  0.07 0.355 0.19 0.455 ;
      RECT  0.07 0.455 1.23 0.545 ;
      RECT  0.07 0.545 0.75 0.575 ;
      RECT  1.24 1.205 1.93 1.325 ;
      RECT  1.81 1.325 1.93 1.425 ;
  END
END SEN_OAI22_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_T_1P5
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_T_1P5
  CLASS CORE ;
  FOREIGN SEN_OAI22_T_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.85 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1506 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1398 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1398 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.36 1.415 0.49 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  2.285 1.415 2.415 1.75 ;
      RECT  2.81 1.21 2.93 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  0.325 0.05 0.455 0.385 ;
      RECT  0.845 0.05 0.975 0.385 ;
      RECT  1.41 0.05 1.54 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.955 0.435 2.695 0.555 ;
      RECT  2.15 0.555 2.25 1.0 ;
      RECT  1.74 1.0 2.25 1.1 ;
      RECT  1.74 1.1 1.86 1.22 ;
      RECT  0.86 1.22 1.86 1.34 ;
    END
    ANTENNADIFFAREA 0.352 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.72 0.215 2.93 0.335 ;
      RECT  2.81 0.335 2.93 0.435 ;
      RECT  1.72 0.335 1.84 0.475 ;
      RECT  0.07 0.375 0.19 0.475 ;
      RECT  0.07 0.475 1.84 0.595 ;
      RECT  0.07 1.205 0.77 1.325 ;
      RECT  0.07 1.325 0.19 1.425 ;
      RECT  0.65 1.325 0.77 1.455 ;
      RECT  0.65 1.455 1.34 1.575 ;
      RECT  2.03 1.205 2.72 1.325 ;
      RECT  2.03 1.325 2.15 1.455 ;
      RECT  1.43 1.455 2.15 1.575 ;
  END
END SEN_OAI22_T_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_T_2
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_T_2
  CLASS CORE ;
  FOREIGN SEN_OAI22_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.65 0.895 ;
      RECT  2.15 0.895 2.25 1.14 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.65 0.91 ;
      RECT  3.55 0.91 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2016 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1872 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1872 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.51 1.415 0.64 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  2.815 1.415 2.945 1.75 ;
      RECT  3.335 1.415 3.465 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.425 0.05 0.555 0.385 ;
      RECT  0.945 0.05 1.075 0.385 ;
      RECT  1.465 0.05 1.595 0.385 ;
      RECT  1.985 0.05 2.115 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.6 0.295 3.72 0.4 ;
      RECT  2.46 0.4 3.72 0.515 ;
      RECT  2.75 0.515 2.85 1.0 ;
      RECT  2.35 1.0 2.85 1.09 ;
      RECT  2.35 1.09 2.45 1.23 ;
      RECT  1.16 1.23 2.45 1.35 ;
    END
    ANTENNADIFFAREA 0.468 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.25 0.2 3.505 0.31 ;
      RECT  2.25 0.31 2.37 0.475 ;
      RECT  0.12 0.475 2.37 0.595 ;
      RECT  0.12 1.2 1.025 1.325 ;
      RECT  0.905 1.325 1.025 1.465 ;
      RECT  0.905 1.465 1.645 1.585 ;
      RECT  2.56 1.205 3.72 1.325 ;
      RECT  3.6 1.325 3.72 1.425 ;
      RECT  2.56 1.325 2.68 1.465 ;
      RECT  1.965 1.465 2.68 1.585 ;
  END
END SEN_OAI22_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_T_3
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_T_3
  CLASS CORE ;
  FOREIGN SEN_OAI22_T_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.69 4.05 0.89 ;
      RECT  3.55 0.89 3.65 0.98 ;
      RECT  2.94 0.98 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1944 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.71 5.25 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3024 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.45 0.89 ;
      RECT  1.75 0.89 1.85 0.91 ;
      RECT  1.35 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.25 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2808 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.08 1.21 0.2 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.595 1.415 0.725 1.75 ;
      RECT  3.54 1.39 3.67 1.75 ;
      RECT  4.09 1.4 4.22 1.75 ;
      RECT  4.61 1.4 4.74 1.75 ;
      RECT  5.13 1.4 5.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.335 0.05 0.465 0.385 ;
      RECT  0.855 0.05 0.985 0.385 ;
      RECT  1.375 0.05 1.505 0.385 ;
      RECT  1.895 0.05 2.025 0.385 ;
      RECT  2.415 0.05 2.545 0.385 ;
      RECT  2.935 0.05 3.06 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.425 5.305 0.545 ;
      RECT  3.35 0.545 3.45 0.71 ;
      RECT  2.75 0.71 3.45 0.89 ;
      RECT  2.75 0.89 2.85 1.205 ;
      RECT  1.095 1.205 3.11 1.325 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.15 0.215 5.515 0.335 ;
      RECT  5.395 0.335 5.515 0.435 ;
      RECT  3.15 0.335 3.25 0.475 ;
      RECT  0.08 0.375 0.2 0.475 ;
      RECT  0.08 0.475 3.25 0.595 ;
      RECT  3.225 1.19 5.515 1.28 ;
      RECT  3.835 1.28 5.515 1.31 ;
      RECT  3.225 1.28 3.345 1.43 ;
      RECT  5.395 1.31 5.515 1.41 ;
      RECT  3.835 1.31 3.955 1.57 ;
      RECT  2.16 1.43 3.345 1.55 ;
      RECT  2.16 1.55 2.28 1.635 ;
      RECT  0.29 1.205 0.98 1.325 ;
      RECT  0.86 1.325 0.98 1.43 ;
      RECT  0.86 1.43 2.07 1.55 ;
  END
END SEN_OAI22_T_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_T_4
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_T_4
  CLASS CORE ;
  FOREIGN SEN_OAI22_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.71 4.85 0.89 ;
      RECT  4.15 0.89 4.25 0.91 ;
      RECT  3.55 0.91 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.25 0.89 ;
      RECT  5.15 0.89 5.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4032 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 3.25 0.89 ;
      RECT  2.15 0.89 2.25 0.91 ;
      RECT  1.75 0.91 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.65 0.9 ;
      RECT  0.75 0.9 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3744 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  4.745 1.435 4.87 1.75 ;
      RECT  5.26 1.435 5.39 1.75 ;
      RECT  5.78 1.435 5.91 1.75 ;
      RECT  6.3 1.435 6.43 1.75 ;
      RECT  6.82 1.41 6.945 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  1.88 0.05 2.01 0.385 ;
      RECT  2.4 0.05 2.53 0.385 ;
      RECT  2.92 0.05 3.05 0.385 ;
      RECT  3.44 0.05 3.57 0.385 ;
      RECT  3.96 0.05 4.09 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.435 0.41 6.735 0.52 ;
      RECT  4.95 0.52 5.05 1.01 ;
      RECT  4.35 1.01 5.05 1.1 ;
      RECT  4.35 1.1 4.45 1.255 ;
      RECT  1.34 1.255 4.45 1.375 ;
    END
    ANTENNADIFFAREA 0.868 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.225 0.205 6.945 0.32 ;
      RECT  6.825 0.32 6.945 0.41 ;
      RECT  4.225 0.32 4.345 0.475 ;
      RECT  0.065 0.375 0.185 0.475 ;
      RECT  0.065 0.475 4.345 0.595 ;
      RECT  0.065 1.205 1.225 1.325 ;
      RECT  0.065 1.325 0.185 1.425 ;
      RECT  1.105 1.325 1.225 1.465 ;
      RECT  1.105 1.465 2.81 1.585 ;
      RECT  4.55 1.225 6.735 1.345 ;
      RECT  4.55 1.345 4.65 1.465 ;
      RECT  2.9 1.465 4.65 1.585 ;
  END
END SEN_OAI22_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI22_T_8
#      Description : "Two 2-input ORs into 2-input NAND"
#      Equation    : X=!((A1|A2)&(B1|B2))
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI22_T_8
  CLASS CORE ;
  FOREIGN SEN_OAI22_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 8.895 0.89 ;
      RECT  7.35 0.89 7.45 0.98 ;
      RECT  5.945 0.98 7.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.15 0.71 12.65 0.89 ;
      RECT  9.35 0.89 10.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8064 ;
  END A2
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 7.115 0.89 ;
      RECT  3.95 0.89 4.05 0.91 ;
      RECT  3.15 0.91 4.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7488 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 3.05 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7488 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.415 0.45 1.75 ;
      RECT  0.0 1.75 13.4 1.85 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  1.36 1.415 1.49 1.75 ;
      RECT  1.88 1.415 2.01 1.75 ;
      RECT  8.365 1.485 8.535 1.75 ;
      RECT  8.885 1.485 9.055 1.75 ;
      RECT  9.405 1.485 9.575 1.75 ;
      RECT  9.945 1.415 10.075 1.75 ;
      RECT  10.465 1.415 10.595 1.75 ;
      RECT  10.985 1.415 11.115 1.75 ;
      RECT  11.505 1.415 11.635 1.75 ;
      RECT  12.045 1.415 12.175 1.75 ;
      RECT  12.62 1.415 12.75 1.75 ;
      RECT  13.19 1.21 13.31 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 13.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 13.4 0.05 ;
      RECT  3.44 0.05 3.57 0.36 ;
      RECT  3.96 0.05 4.09 0.36 ;
      RECT  4.48 0.05 4.61 0.36 ;
      RECT  5.0 0.05 5.13 0.36 ;
      RECT  5.52 0.05 5.65 0.36 ;
      RECT  6.04 0.05 6.17 0.36 ;
      RECT  6.56 0.05 6.69 0.36 ;
      RECT  7.08 0.05 7.21 0.36 ;
      RECT  7.6 0.05 7.73 0.36 ;
      RECT  8.12 0.05 8.25 0.36 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  1.88 0.05 2.01 0.385 ;
      RECT  2.4 0.05 2.53 0.385 ;
      RECT  2.92 0.05 3.05 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 13.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.62 0.42 13.085 0.54 ;
      RECT  9.08 0.54 13.085 0.55 ;
      RECT  9.08 0.55 11.555 0.59 ;
      RECT  9.08 0.59 9.25 0.98 ;
      RECT  7.55 0.98 9.25 1.15 ;
      RECT  7.55 1.15 7.75 1.205 ;
      RECT  4.15 1.205 7.75 1.255 ;
      RECT  2.38 1.255 7.75 1.375 ;
    END
    ANTENNADIFFAREA 1.731 ;
  END X
  OBS
      LAYER M1 ;
      RECT  8.36 0.16 11.83 0.21 ;
      RECT  8.36 0.21 13.3 0.33 ;
      RECT  13.18 0.33 13.3 0.43 ;
      RECT  8.36 0.33 8.53 0.45 ;
      RECT  3.435 0.45 8.53 0.485 ;
      RECT  0.065 0.4 0.185 0.485 ;
      RECT  0.065 0.485 8.53 0.62 ;
      RECT  9.415 1.185 13.09 1.24 ;
      RECT  7.935 1.24 13.09 1.325 ;
      RECT  7.935 1.325 9.575 1.395 ;
      RECT  7.935 1.395 8.135 1.465 ;
      RECT  5.215 1.465 8.135 1.585 ;
      RECT  7.28 1.585 8.135 1.61 ;
      RECT  0.065 1.185 2.29 1.325 ;
      RECT  0.065 1.325 0.185 1.405 ;
      RECT  2.12 1.325 2.29 1.465 ;
      RECT  2.12 1.465 4.915 1.585 ;
  END
END SEN_OAI22_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_1
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_1
  CLASS CORE ;
  FOREIGN SEN_OAI31_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.67 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.505 0.92 ;
      RECT  0.35 0.92 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.7 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0642 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.16 1.575 1.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.595 0.05 0.725 0.38 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 1.38 ;
      RECT  0.82 1.38 1.25 1.48 ;
    END
    ANTENNADIFFAREA 0.207 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.37 0.455 0.47 ;
      RECT  0.34 0.47 1.03 0.59 ;
  END
END SEN_OAI31_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_2
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_2
  CLASS CORE ;
  FOREIGN SEN_OAI31_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 0.7 ;
      RECT  0.15 0.7 0.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1284 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.41 0.455 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  2.135 1.44 2.27 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.585 0.05 0.715 0.36 ;
      RECT  1.105 0.05 1.235 0.36 ;
      RECT  1.615 0.05 1.745 0.36 ;
      RECT  0.065 0.05 0.195 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.47 2.25 1.23 ;
      RECT  1.335 1.23 2.52 1.35 ;
      RECT  2.4 1.35 2.52 1.45 ;
    END
    ANTENNADIFFAREA 0.412 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.875 0.17 2.52 0.29 ;
      RECT  2.4 0.29 2.52 0.39 ;
      RECT  1.875 0.29 2.0 0.45 ;
      RECT  0.34 0.35 0.45 0.45 ;
      RECT  0.34 0.45 2.0 0.57 ;
      RECT  1.11 1.1 1.23 1.21 ;
      RECT  0.07 1.21 1.23 1.32 ;
      RECT  0.07 1.32 0.19 1.43 ;
      RECT  0.8 1.45 1.79 1.57 ;
  END
END SEN_OAI31_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_3
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_3
  CLASS CORE ;
  FOREIGN SEN_OAI31_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.25 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.65 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1926 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  0.585 1.44 0.715 1.75 ;
      RECT  2.665 1.44 2.795 1.75 ;
      RECT  3.2 1.21 3.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.585 0.05 0.715 0.38 ;
      RECT  1.105 0.05 1.235 0.38 ;
      RECT  1.625 0.05 1.755 0.38 ;
      RECT  2.145 0.05 2.275 0.38 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.64 0.47 3.335 0.59 ;
      RECT  2.75 0.59 2.85 1.22 ;
      RECT  1.84 1.22 3.075 1.34 ;
    END
    ANTENNADIFFAREA 0.529 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.41 0.24 3.09 0.36 ;
      RECT  2.41 0.36 2.53 0.47 ;
      RECT  0.305 0.47 2.53 0.59 ;
      RECT  0.305 1.23 1.54 1.35 ;
      RECT  1.06 1.45 2.32 1.57 ;
  END
END SEN_OAI31_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_4
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_4
  CLASS CORE ;
  FOREIGN SEN_OAI31_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2568 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.455 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.845 1.44 0.975 1.75 ;
      RECT  3.64 1.44 3.77 1.75 ;
      RECT  4.16 1.44 4.29 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.345 0.05 0.475 0.37 ;
      RECT  0.895 0.05 1.025 0.37 ;
      RECT  1.435 0.05 1.565 0.37 ;
      RECT  2.005 0.05 2.135 0.37 ;
      RECT  2.59 0.05 2.72 0.37 ;
      RECT  3.12 0.05 3.25 0.37 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.46 4.33 0.58 ;
      RECT  3.55 0.58 3.65 1.205 ;
      RECT  3.55 1.205 4.545 1.21 ;
      RECT  2.32 1.015 2.65 1.135 ;
      RECT  2.55 1.135 2.65 1.21 ;
      RECT  2.55 1.21 4.545 1.32 ;
      RECT  4.425 1.32 4.545 1.61 ;
    END
    ANTENNADIFFAREA 0.711 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.345 0.23 4.545 0.35 ;
      RECT  4.425 0.35 4.545 0.4 ;
      RECT  3.345 0.35 3.45 0.46 ;
      RECT  0.07 0.36 0.19 0.46 ;
      RECT  0.07 0.46 3.45 0.58 ;
      RECT  0.07 1.23 2.27 1.35 ;
      RECT  2.15 1.35 2.27 1.41 ;
      RECT  0.07 1.35 0.19 1.45 ;
      RECT  1.32 1.44 2.06 1.52 ;
      RECT  1.32 1.52 3.3 1.56 ;
      RECT  2.55 1.44 3.3 1.52 ;
      RECT  1.93 1.56 2.685 1.62 ;
  END
END SEN_OAI31_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_12
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_12
  CLASS CORE ;
  FOREIGN SEN_OAI31_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  9.22 0.735 9.45 0.89 ;
      RECT  9.22 0.89 9.32 1.29 ;
      RECT  7.95 0.71 8.05 1.15 ;
      RECT  7.87 1.15 8.05 1.25 ;
      RECT  6.35 0.71 6.45 1.29 ;
      RECT  4.75 0.71 4.85 1.29 ;
      RECT  3.15 0.71 3.25 1.29 ;
      RECT  1.55 0.71 1.66 1.29 ;
      RECT  0.15 0.71 0.25 1.29 ;
      LAYER M2 ;
      RECT  0.11 1.15 9.36 1.25 ;
      LAYER V1 ;
      RECT  9.22 1.15 9.32 1.25 ;
      RECT  7.91 1.15 8.01 1.25 ;
      RECT  6.35 1.15 6.45 1.25 ;
      RECT  4.75 1.15 4.85 1.25 ;
      RECT  3.15 1.15 3.25 1.25 ;
      RECT  1.55 1.15 1.65 1.25 ;
      RECT  0.15 1.15 0.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7452 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.95 0.735 9.13 0.89 ;
      RECT  8.95 0.89 9.05 1.045 ;
      RECT  8.15 0.735 8.45 0.89 ;
      RECT  8.15 0.89 8.25 1.045 ;
      RECT  7.35 0.71 7.65 0.89 ;
      RECT  7.53 0.89 7.65 1.07 ;
      RECT  6.55 0.71 6.85 0.89 ;
      RECT  6.75 0.89 6.85 1.05 ;
      RECT  5.75 0.71 6.05 0.89 ;
      RECT  5.75 0.89 5.85 1.05 ;
      RECT  5.15 0.71 5.385 0.89 ;
      RECT  5.15 0.89 5.25 1.05 ;
      RECT  4.35 0.71 4.65 0.89 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  2.745 0.71 3.05 0.89 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  0.35 0.71 0.65 0.9 ;
      LAYER M2 ;
      RECT  0.31 0.75 9.13 0.85 ;
      LAYER V1 ;
      RECT  8.99 0.75 9.09 0.85 ;
      RECT  8.305 0.75 8.405 0.85 ;
      RECT  7.35 0.75 7.45 0.85 ;
      RECT  7.55 0.75 7.65 0.85 ;
      RECT  6.55 0.75 6.65 0.85 ;
      RECT  6.75 0.75 6.85 0.85 ;
      RECT  5.75 0.75 5.85 0.85 ;
      RECT  5.95 0.75 6.05 0.85 ;
      RECT  5.15 0.75 5.25 0.85 ;
      RECT  4.35 0.75 4.45 0.85 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
      RECT  0.35 0.75 0.45 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7452 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.66 0.735 8.77 0.95 ;
      RECT  8.53 0.95 8.77 1.05 ;
      RECT  7.145 0.715 7.255 0.95 ;
      RECT  6.99 0.95 7.255 1.05 ;
      RECT  5.545 0.71 5.655 0.95 ;
      RECT  5.475 0.95 5.655 1.05 ;
      RECT  3.945 0.71 4.055 1.095 ;
      RECT  2.345 0.71 2.455 1.095 ;
      RECT  0.745 0.71 0.855 1.095 ;
      LAYER M2 ;
      RECT  0.71 0.95 8.77 1.05 ;
      LAYER V1 ;
      RECT  8.63 0.95 8.73 1.05 ;
      RECT  7.065 0.95 7.165 1.05 ;
      RECT  5.515 0.95 5.615 1.05 ;
      RECT  3.95 0.95 4.05 1.05 ;
      RECT  2.35 0.95 2.45 1.05 ;
      RECT  0.75 0.95 0.85 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7452 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.65 0.71 12.65 0.785 ;
      RECT  10.135 0.785 12.65 0.89 ;
      RECT  12.55 0.89 12.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7344 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.84 1.4 0.97 1.75 ;
      RECT  0.0 1.75 12.8 1.85 ;
      RECT  2.4 1.42 2.53 1.75 ;
      RECT  3.96 1.425 4.09 1.75 ;
      RECT  5.52 1.415 5.665 1.75 ;
      RECT  7.06 1.46 7.23 1.75 ;
      RECT  8.62 1.48 8.79 1.75 ;
      RECT  9.75 1.415 9.865 1.75 ;
      RECT  10.255 1.415 10.385 1.75 ;
      RECT  10.775 1.415 10.905 1.75 ;
      RECT  11.295 1.415 11.425 1.75 ;
      RECT  11.815 1.415 11.945 1.75 ;
      RECT  12.335 1.415 12.46 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      RECT  6.54 0.05 6.71 0.305 ;
      RECT  7.06 0.05 7.23 0.305 ;
      RECT  7.58 0.05 7.75 0.305 ;
      RECT  8.1 0.05 8.27 0.305 ;
      RECT  8.62 0.05 8.79 0.305 ;
      RECT  9.14 0.05 9.31 0.305 ;
      RECT  4.46 0.05 4.63 0.345 ;
      RECT  4.98 0.05 5.15 0.345 ;
      RECT  5.5 0.05 5.67 0.345 ;
      RECT  6.02 0.05 6.19 0.345 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  1.88 0.05 2.01 0.385 ;
      RECT  2.4 0.05 2.53 0.385 ;
      RECT  2.92 0.05 3.05 0.385 ;
      RECT  3.44 0.05 3.57 0.385 ;
      RECT  3.96 0.05 4.085 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  10.32 0.44 12.51 0.485 ;
      RECT  9.74 0.485 12.51 0.565 ;
      RECT  9.74 0.565 11.1 0.61 ;
      RECT  9.74 0.61 10.5 0.695 ;
      RECT  9.74 0.695 9.99 1.04 ;
      RECT  9.41 1.04 9.99 1.11 ;
      RECT  9.41 1.11 12.45 1.18 ;
      RECT  9.41 1.18 12.72 1.29 ;
      RECT  9.41 1.29 9.66 1.38 ;
      RECT  12.55 1.29 12.72 1.49 ;
      RECT  6.74 1.16 7.65 1.34 ;
      RECT  6.74 1.34 9.13 1.37 ;
      RECT  8.15 1.14 9.13 1.34 ;
      RECT  7.44 1.37 9.13 1.38 ;
      RECT  6.74 1.37 6.95 1.405 ;
      RECT  7.44 1.38 9.66 1.39 ;
      RECT  7.44 1.39 8.45 1.59 ;
      RECT  8.88 1.39 9.66 1.63 ;
      RECT  5.15 1.14 6.05 1.31 ;
      RECT  5.88 1.31 6.05 1.405 ;
      RECT  5.15 1.31 5.32 1.415 ;
      RECT  5.88 1.405 6.95 1.615 ;
      RECT  3.74 1.205 4.46 1.335 ;
      RECT  4.33 1.335 4.46 1.415 ;
      RECT  3.74 1.335 3.865 1.44 ;
      RECT  4.33 1.415 5.32 1.585 ;
      RECT  2.14 1.205 2.86 1.33 ;
      RECT  2.14 1.33 2.265 1.44 ;
      RECT  2.735 1.33 2.86 1.44 ;
      RECT  0.55 1.215 1.25 1.305 ;
      RECT  0.55 1.305 0.65 1.41 ;
      RECT  1.15 1.305 1.25 1.44 ;
      RECT  0.065 1.41 0.65 1.5 ;
      RECT  1.15 1.44 2.265 1.56 ;
      RECT  2.735 1.44 3.865 1.565 ;
      RECT  0.065 1.5 0.185 1.63 ;
    END
    ANTENNADIFFAREA 2.038 ;
  END X
  OBS
      LAYER M1 ;
      RECT  9.4 0.16 11.35 0.22 ;
      RECT  9.4 0.22 12.72 0.34 ;
      RECT  9.4 0.34 10.255 0.375 ;
      RECT  12.6 0.34 12.72 0.44 ;
      RECT  9.4 0.375 9.65 0.395 ;
      RECT  6.27 0.395 9.65 0.435 ;
      RECT  4.16 0.435 9.65 0.49 ;
      RECT  0.065 0.4 0.185 0.49 ;
      RECT  0.065 0.49 9.65 0.62 ;
      RECT  8.145 0.62 9.65 0.645 ;
  END
END SEN_OAI31_12
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_6
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_6
  CLASS CORE ;
  FOREIGN SEN_OAI31_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.85 0.89 ;
      RECT  4.55 0.89 4.65 1.29 ;
      RECT  3.15 0.71 3.25 1.29 ;
      RECT  1.55 0.71 1.66 1.29 ;
      RECT  0.15 0.71 0.25 1.29 ;
      LAYER M2 ;
      RECT  0.11 1.15 4.695 1.25 ;
      LAYER V1 ;
      RECT  4.55 1.15 4.65 1.25 ;
      RECT  3.15 1.15 3.25 1.25 ;
      RECT  1.55 1.15 1.65 1.25 ;
      RECT  0.15 1.15 0.25 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3726 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.34 0.71 4.46 1.095 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  2.745 0.71 3.05 0.89 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  0.35 0.71 0.65 0.9 ;
      LAYER M2 ;
      RECT  0.31 0.75 4.49 0.85 ;
      LAYER V1 ;
      RECT  4.35 0.75 4.45 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
      RECT  0.35 0.75 0.45 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3726 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.945 0.71 4.055 1.095 ;
      RECT  2.345 0.71 2.455 1.095 ;
      RECT  0.745 0.71 0.855 1.095 ;
      LAYER M2 ;
      RECT  0.71 0.95 4.09 1.05 ;
      LAYER V1 ;
      RECT  3.95 0.95 4.05 1.05 ;
      RECT  2.35 0.95 2.45 1.05 ;
      RECT  0.75 0.95 0.85 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3726 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.33 0.71 6.45 0.89 ;
      RECT  6.35 0.89 6.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3672 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  0.0 1.75 6.6 1.85 ;
      RECT  2.4 1.42 2.53 1.75 ;
      RECT  3.96 1.425 4.09 1.75 ;
      RECT  5.035 1.415 5.165 1.75 ;
      RECT  5.555 1.415 5.685 1.75 ;
      RECT  6.075 1.415 6.205 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  1.88 0.05 2.01 0.385 ;
      RECT  2.4 0.05 2.53 0.385 ;
      RECT  2.92 0.05 3.05 0.385 ;
      RECT  3.44 0.05 3.57 0.385 ;
      RECT  3.96 0.05 4.09 0.385 ;
      RECT  4.48 0.05 4.61 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.44 6.25 0.57 ;
      RECT  4.95 0.57 5.08 1.11 ;
      RECT  4.75 1.11 6.25 1.18 ;
      RECT  4.75 1.18 6.51 1.29 ;
      RECT  4.75 1.29 4.88 1.435 ;
      RECT  3.74 1.205 4.46 1.335 ;
      RECT  4.33 1.335 4.46 1.435 ;
      RECT  3.74 1.335 3.865 1.44 ;
      RECT  4.33 1.435 4.88 1.565 ;
      RECT  2.14 1.205 2.86 1.33 ;
      RECT  2.14 1.33 2.265 1.44 ;
      RECT  2.735 1.33 2.86 1.44 ;
      RECT  0.55 1.215 1.25 1.305 ;
      RECT  0.55 1.305 0.65 1.41 ;
      RECT  1.15 1.305 1.25 1.44 ;
      RECT  0.065 1.41 0.65 1.5 ;
      RECT  1.15 1.44 2.265 1.56 ;
      RECT  2.735 1.44 3.865 1.565 ;
      RECT  0.065 1.5 0.185 1.63 ;
    END
    ANTENNADIFFAREA 1.06 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.73 0.22 6.51 0.35 ;
      RECT  4.73 0.35 4.86 0.48 ;
      RECT  0.065 0.39 0.185 0.48 ;
      RECT  0.065 0.48 4.86 0.61 ;
  END
END SEN_OAI31_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_8
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_8
  CLASS CORE ;
  FOREIGN SEN_OAI31_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.25 1.29 ;
      RECT  4.75 0.71 4.85 1.29 ;
      RECT  3.15 0.71 3.25 1.29 ;
      RECT  1.55 0.71 1.66 1.29 ;
      RECT  0.15 0.71 0.25 1.15 ;
      RECT  0.15 1.15 0.42 1.25 ;
      LAYER M2 ;
      RECT  0.18 1.15 6.29 1.25 ;
      LAYER V1 ;
      RECT  6.15 1.15 6.25 1.25 ;
      RECT  4.75 1.15 4.85 1.25 ;
      RECT  3.15 1.15 3.25 1.25 ;
      RECT  1.55 1.15 1.65 1.25 ;
      RECT  0.25 1.15 0.35 1.25 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4968 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.71 6.05 0.89 ;
      RECT  5.75 0.89 5.85 1.05 ;
      RECT  5.15 0.71 5.385 0.89 ;
      RECT  5.15 0.89 5.25 1.05 ;
      RECT  4.35 0.71 4.65 0.89 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  2.745 0.71 3.05 0.89 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.15 0.71 1.45 0.89 ;
      RECT  0.35 0.71 0.65 0.9 ;
      LAYER M2 ;
      RECT  0.31 0.75 6.09 0.85 ;
      LAYER V1 ;
      RECT  5.75 0.75 5.85 0.85 ;
      RECT  5.95 0.75 6.05 0.85 ;
      RECT  5.15 0.75 5.25 0.85 ;
      RECT  4.35 0.75 4.45 0.85 ;
      RECT  4.55 0.75 4.65 0.85 ;
      RECT  3.55 0.75 3.65 0.85 ;
      RECT  3.75 0.75 3.85 0.85 ;
      RECT  2.75 0.75 2.85 0.85 ;
      RECT  2.95 0.75 3.05 0.85 ;
      RECT  1.95 0.75 2.05 0.85 ;
      RECT  2.15 0.75 2.25 0.85 ;
      RECT  1.15 0.75 1.25 0.85 ;
      RECT  1.35 0.75 1.45 0.85 ;
      RECT  0.35 0.75 0.45 0.85 ;
      RECT  0.55 0.75 0.65 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4968 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.545 0.71 5.655 0.95 ;
      RECT  5.475 0.95 5.655 1.05 ;
      RECT  3.945 0.71 4.055 1.095 ;
      RECT  2.345 0.71 2.455 1.095 ;
      RECT  0.745 0.71 0.855 1.095 ;
      LAYER M2 ;
      RECT  0.71 0.95 5.655 1.05 ;
      LAYER V1 ;
      RECT  5.515 0.95 5.615 1.05 ;
      RECT  3.95 0.95 4.05 1.05 ;
      RECT  2.35 0.95 2.45 1.05 ;
      RECT  0.75 0.95 0.85 1.05 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4968 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.93 0.71 8.45 0.89 ;
      RECT  8.35 0.89 8.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.84 1.415 0.97 1.75 ;
      RECT  0.0 1.75 8.6 1.85 ;
      RECT  2.4 1.42 2.53 1.75 ;
      RECT  3.96 1.425 4.09 1.75 ;
      RECT  5.52 1.415 5.665 1.75 ;
      RECT  6.6 1.415 6.715 1.75 ;
      RECT  7.105 1.415 7.235 1.75 ;
      RECT  7.625 1.415 7.755 1.75 ;
      RECT  8.145 1.415 8.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      RECT  4.48 0.05 4.61 0.35 ;
      RECT  5.0 0.05 5.13 0.35 ;
      RECT  5.52 0.05 5.65 0.35 ;
      RECT  6.04 0.05 6.17 0.35 ;
      RECT  0.32 0.05 0.45 0.385 ;
      RECT  0.84 0.05 0.97 0.385 ;
      RECT  1.36 0.05 1.49 0.385 ;
      RECT  1.88 0.05 2.01 0.385 ;
      RECT  2.4 0.05 2.53 0.385 ;
      RECT  2.92 0.05 3.05 0.385 ;
      RECT  3.44 0.05 3.57 0.385 ;
      RECT  3.96 0.05 4.09 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.55 0.44 8.32 0.57 ;
      RECT  6.55 0.57 6.72 1.11 ;
      RECT  6.34 1.11 8.25 1.18 ;
      RECT  6.34 1.18 8.53 1.29 ;
      RECT  8.41 1.29 8.53 1.4 ;
      RECT  6.34 1.29 6.51 1.415 ;
      RECT  5.15 1.14 6.05 1.31 ;
      RECT  5.15 1.31 5.32 1.415 ;
      RECT  5.88 1.31 6.05 1.415 ;
      RECT  3.74 1.205 4.46 1.335 ;
      RECT  4.33 1.335 4.46 1.415 ;
      RECT  3.74 1.335 3.865 1.44 ;
      RECT  4.33 1.415 5.32 1.585 ;
      RECT  5.88 1.415 6.51 1.585 ;
      RECT  2.14 1.205 2.86 1.33 ;
      RECT  2.14 1.33 2.265 1.44 ;
      RECT  2.735 1.33 2.86 1.44 ;
      RECT  0.55 1.215 1.25 1.305 ;
      RECT  0.55 1.305 0.65 1.41 ;
      RECT  1.15 1.305 1.25 1.44 ;
      RECT  0.065 1.41 0.65 1.5 ;
      RECT  1.15 1.44 2.265 1.56 ;
      RECT  2.735 1.44 3.865 1.565 ;
      RECT  0.065 1.5 0.185 1.61 ;
    END
    ANTENNADIFFAREA 1.376 ;
  END X
  OBS
      LAYER M1 ;
      RECT  6.28 0.21 7.11 0.23 ;
      RECT  6.28 0.23 8.53 0.35 ;
      RECT  6.28 0.35 6.45 0.44 ;
      RECT  8.41 0.35 8.53 0.45 ;
      RECT  4.17 0.44 6.45 0.48 ;
      RECT  0.065 0.39 0.185 0.48 ;
      RECT  0.065 0.48 6.45 0.61 ;
  END
END SEN_OAI31_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_0P5
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI31_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.91 ;
      RECT  0.35 0.91 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.845 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.155 1.41 1.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.595 0.05 0.725 0.385 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.19 1.25 0.665 ;
      RECT  0.95 0.665 1.25 0.755 ;
      RECT  0.95 0.755 1.05 1.44 ;
      RECT  0.83 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.095 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.19 0.445 0.485 ;
      RECT  0.34 0.485 1.0 0.575 ;
      RECT  0.88 0.19 1.0 0.485 ;
  END
END SEN_OAI31_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_0P75
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_0P75
  CLASS CORE ;
  FOREIGN SEN_OAI31_0P75 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0462 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.845 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0459 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.155 1.415 1.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.595 0.05 0.725 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.29 1.25 0.665 ;
      RECT  0.95 0.665 1.25 0.755 ;
      RECT  0.95 0.755 1.05 1.44 ;
      RECT  0.83 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.141 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.29 0.445 0.485 ;
      RECT  0.34 0.485 1.0 0.575 ;
      RECT  0.88 0.29 1.0 0.485 ;
  END
END SEN_OAI31_0P75
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_T_0P5
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_T_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI31_T_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.91 0.65 1.09 ;
      RECT  0.35 1.09 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0441 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.845 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0309 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.155 1.41 1.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.595 0.05 0.725 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.2 1.25 0.665 ;
      RECT  0.95 0.665 1.25 0.755 ;
      RECT  0.95 0.755 1.05 1.44 ;
      RECT  0.83 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.095 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.23 0.445 0.485 ;
      RECT  0.34 0.485 1.0 0.575 ;
      RECT  0.88 0.23 1.0 0.485 ;
  END
END SEN_OAI31_T_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_T_1
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_T_1
  CLASS CORE ;
  FOREIGN SEN_OAI31_T_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0882 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.945 0.71 1.05 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0882 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0882 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.905 ;
      RECT  1.55 0.905 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0612 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.305 1.41 0.435 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.915 1.41 2.045 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.33 0.05 0.46 0.385 ;
      RECT  0.85 0.05 0.98 0.385 ;
      RECT  1.37 0.05 1.5 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.945 0.29 2.05 1.11 ;
      RECT  1.75 1.11 2.05 1.2 ;
      RECT  1.585 1.2 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.208 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.075 0.375 0.195 0.475 ;
      RECT  0.075 0.475 1.805 0.595 ;
  END
END SEN_OAI31_T_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_T_2
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_T_2
  CLASS CORE ;
  FOREIGN SEN_OAI31_T_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 2.85 0.91 ;
      RECT  2.15 0.91 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1764 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 1.85 0.91 ;
      RECT  1.35 0.91 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1764 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.965 ;
      RECT  0.95 0.965 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1764 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.71 3.65 0.9 ;
      RECT  3.55 0.9 3.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1224 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.385 1.21 0.505 1.75 ;
      RECT  0.0 1.75 3.8 1.85 ;
      RECT  0.92 1.415 1.05 1.75 ;
      RECT  3.005 1.415 3.135 1.75 ;
      RECT  3.56 1.21 3.68 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      RECT  0.4 0.05 0.53 0.385 ;
      RECT  0.92 0.05 1.05 0.385 ;
      RECT  1.44 0.05 1.57 0.385 ;
      RECT  1.96 0.05 2.09 0.385 ;
      RECT  2.48 0.05 2.61 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.38 3.15 0.4 ;
      RECT  2.95 0.4 3.66 0.49 ;
      RECT  3.54 0.28 3.66 0.4 ;
      RECT  2.95 0.49 3.05 1.205 ;
      RECT  2.175 1.205 3.45 1.325 ;
      RECT  3.35 1.325 3.45 1.49 ;
    END
    ANTENNADIFFAREA 0.342 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.745 0.2 3.45 0.29 ;
      RECT  3.255 0.29 3.45 0.31 ;
      RECT  2.745 0.29 2.86 0.475 ;
      RECT  0.095 0.475 2.86 0.595 ;
      RECT  0.615 1.205 1.875 1.325 ;
      RECT  1.395 1.45 2.655 1.57 ;
  END
END SEN_OAI31_T_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_T_4
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_T_4
  CLASS CORE ;
  FOREIGN SEN_OAI31_T_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 4.65 0.91 ;
      RECT  3.95 0.91 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3528 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 2.85 0.91 ;
      RECT  2.15 0.91 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3528 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.25 0.91 ;
      RECT  0.55 0.91 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3528 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.51 6.25 0.71 ;
      RECT  5.55 0.71 6.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2448 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.365 1.415 0.495 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  0.885 1.415 1.015 1.75 ;
      RECT  1.405 1.415 1.535 1.75 ;
      RECT  5.335 1.415 5.465 1.75 ;
      RECT  5.855 1.415 5.985 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  0.625 0.05 0.755 0.385 ;
      RECT  1.145 0.05 1.275 0.385 ;
      RECT  1.665 0.05 1.795 0.385 ;
      RECT  2.185 0.05 2.315 0.385 ;
      RECT  2.705 0.05 2.835 0.385 ;
      RECT  3.235 0.05 3.365 0.385 ;
      RECT  3.775 0.05 3.905 0.385 ;
      RECT  4.295 0.05 4.425 0.385 ;
      RECT  4.815 0.05 4.945 0.385 ;
      RECT  0.11 0.05 0.23 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.34 0.44 6.03 0.56 ;
      RECT  5.34 0.56 5.46 1.11 ;
      RECT  5.34 1.11 6.25 1.205 ;
      RECT  3.495 1.205 6.25 1.325 ;
    END
    ANTENNADIFFAREA 0.716 ;
  END X
  OBS
      LAYER M1 ;
      RECT  5.08 0.225 6.29 0.345 ;
      RECT  5.08 0.345 5.2 0.475 ;
      RECT  0.32 0.475 5.2 0.595 ;
      RECT  0.06 1.205 3.375 1.325 ;
      RECT  1.88 1.445 4.99 1.565 ;
  END
END SEN_OAI31_T_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_T_8
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_T_8
  CLASS CORE ;
  FOREIGN SEN_OAI31_T_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.15 0.71 7.25 0.91 ;
      RECT  7.15 0.91 8.66 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7065 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.05 0.91 ;
      RECT  3.95 0.91 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7065 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 0.85 0.91 ;
      RECT  0.75 0.91 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7065 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  11.55 0.51 11.65 0.71 ;
      RECT  10.055 0.71 11.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4896 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.44 0.455 1.75 ;
      RECT  0.0 1.75 11.8 1.85 ;
      RECT  0.845 1.44 0.975 1.75 ;
      RECT  1.365 1.44 1.495 1.75 ;
      RECT  1.885 1.44 2.015 1.75 ;
      RECT  2.405 1.44 2.535 1.75 ;
      RECT  2.925 1.44 3.055 1.75 ;
      RECT  9.75 1.44 9.88 1.75 ;
      RECT  10.27 1.415 10.4 1.75 ;
      RECT  10.79 1.415 10.92 1.75 ;
      RECT  11.31 1.415 11.44 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.8 0.05 ;
      RECT  2.145 0.05 2.275 0.36 ;
      RECT  2.665 0.05 2.795 0.36 ;
      RECT  3.185 0.05 3.315 0.36 ;
      RECT  3.705 0.05 3.835 0.36 ;
      RECT  4.225 0.05 4.355 0.36 ;
      RECT  4.745 0.05 4.875 0.36 ;
      RECT  5.265 0.05 5.395 0.36 ;
      RECT  5.785 0.05 5.915 0.36 ;
      RECT  6.57 0.05 6.7 0.36 ;
      RECT  7.09 0.05 7.22 0.36 ;
      RECT  7.61 0.05 7.74 0.36 ;
      RECT  8.13 0.05 8.26 0.36 ;
      RECT  8.65 0.05 8.78 0.36 ;
      RECT  9.2 0.05 9.33 0.36 ;
      RECT  0.585 0.05 0.715 0.385 ;
      RECT  1.105 0.05 1.235 0.385 ;
      RECT  1.625 0.05 1.755 0.385 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  9.75 0.45 11.46 0.58 ;
      RECT  9.75 0.58 9.92 1.11 ;
      RECT  8.75 1.11 11.695 1.225 ;
      RECT  6.265 1.225 11.695 1.29 ;
      RECT  6.265 1.29 10.075 1.35 ;
    END
    ANTENNADIFFAREA 1.357 ;
  END X
  OBS
      LAYER M1 ;
      RECT  9.47 0.205 11.745 0.345 ;
      RECT  9.47 0.345 9.64 0.45 ;
      RECT  2.15 0.45 9.64 0.5 ;
      RECT  0.28 0.5 9.64 0.62 ;
      RECT  2.45 1.18 4.04 1.225 ;
      RECT  0.07 1.225 4.04 1.23 ;
      RECT  0.07 1.23 5.96 1.35 ;
      RECT  0.07 1.35 0.19 1.445 ;
      RECT  5.275 1.44 7.46 1.48 ;
      RECT  3.4 1.48 9.37 1.61 ;
  END
END SEN_OAI31_T_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_G_0P5
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_G_0P5
  CLASS CORE ;
  FOREIGN SEN_OAI31_G_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.92 ;
      RECT  0.35 0.92 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.835 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.06 1.41 0.19 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.155 1.41 1.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.595 0.05 0.725 0.385 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.21 1.25 0.655 ;
      RECT  0.95 0.655 1.25 0.745 ;
      RECT  0.95 0.745 1.05 1.44 ;
      RECT  0.83 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.098 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.21 0.445 0.475 ;
      RECT  0.34 0.475 1.0 0.565 ;
      RECT  0.88 0.21 1.0 0.475 ;
  END
END SEN_OAI31_G_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_G_1
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_G_1
  CLASS CORE ;
  FOREIGN SEN_OAI31_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.71 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.795 1.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.155 1.41 1.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.575 0.05 0.745 0.345 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.29 1.25 0.615 ;
      RECT  0.95 0.615 1.25 0.705 ;
      RECT  0.95 0.705 1.05 1.44 ;
      RECT  0.83 1.44 1.05 1.56 ;
    END
    ANTENNADIFFAREA 0.197 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.305 0.445 0.435 ;
      RECT  0.34 0.435 1.0 0.525 ;
      RECT  0.88 0.305 1.0 0.435 ;
  END
END SEN_OAI31_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_G_2
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_G_2
  CLASS CORE ;
  FOREIGN SEN_OAI31_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 1.85 0.9 ;
      RECT  1.15 0.9 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.9 ;
      RECT  0.95 0.9 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.9 ;
      RECT  0.35 0.9 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.51 2.45 0.96 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.415 0.455 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  2.135 1.4 2.265 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.585 0.05 0.715 0.385 ;
      RECT  1.105 0.05 1.235 0.385 ;
      RECT  1.615 0.05 1.745 0.385 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.47 2.25 1.11 ;
      RECT  1.35 1.11 2.52 1.29 ;
    END
    ANTENNADIFFAREA 0.408 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.4 0.17 2.52 0.26 ;
      RECT  1.88 0.26 2.52 0.38 ;
      RECT  1.88 0.38 2.0 0.475 ;
      RECT  0.28 0.475 2.0 0.595 ;
      RECT  0.07 1.205 1.26 1.325 ;
      RECT  0.07 1.325 0.19 1.425 ;
      RECT  0.8 1.44 1.79 1.56 ;
  END
END SEN_OAI31_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI31_G_4
#      Description : "3-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI31_G_4
  CLASS CORE ;
  FOREIGN SEN_OAI31_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 3.25 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A3
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.415 0.44 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.83 1.415 0.96 1.75 ;
      RECT  3.635 1.41 3.765 1.75 ;
      RECT  4.155 1.41 4.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.31 0.05 0.44 0.385 ;
      RECT  0.83 0.05 0.96 0.385 ;
      RECT  1.35 0.05 1.48 0.385 ;
      RECT  1.87 0.05 2.0 0.385 ;
      RECT  2.595 0.05 2.725 0.385 ;
      RECT  3.115 0.05 3.245 0.385 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.45 4.33 0.57 ;
      RECT  3.55 0.57 3.65 1.11 ;
      RECT  2.34 0.99 2.65 1.11 ;
      RECT  2.34 1.11 4.25 1.16 ;
      RECT  2.55 1.16 4.25 1.2 ;
      RECT  2.55 1.2 4.54 1.29 ;
      RECT  4.42 1.29 4.54 1.61 ;
    END
    ANTENNADIFFAREA 0.706 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.35 0.215 4.54 0.335 ;
      RECT  4.42 0.335 4.54 0.41 ;
      RECT  3.35 0.335 3.45 0.475 ;
      RECT  0.055 0.475 3.45 0.595 ;
      RECT  0.055 0.595 0.175 0.705 ;
      RECT  1.305 1.22 2.02 1.25 ;
      RECT  1.305 1.25 2.445 1.34 ;
      RECT  2.355 1.34 2.445 1.44 ;
      RECT  2.355 1.44 3.29 1.56 ;
      RECT  0.055 1.205 1.215 1.325 ;
      RECT  1.095 1.325 1.215 1.43 ;
      RECT  0.055 1.325 0.175 1.61 ;
      RECT  1.095 1.43 2.255 1.55 ;
      RECT  2.135 1.55 2.255 1.625 ;
  END
END SEN_OAI31_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI41_1
#      Description : "4-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3|A4)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI41_1
  CLASS CORE ;
  FOREIGN SEN_OAI41_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.945 0.69 1.06 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.057 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.695 0.685 0.85 0.88 ;
      RECT  0.75 0.88 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.057 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.58 0.88 ;
      RECT  0.35 0.88 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.057 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.685 0.26 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.057 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.815 1.52 0.935 ;
      RECT  1.35 0.935 1.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0501 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.41 0.195 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.41 1.41 1.54 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.305 0.05 0.475 0.325 ;
      RECT  0.825 0.05 0.995 0.325 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.29 1.52 0.625 ;
      RECT  1.15 0.625 1.52 0.715 ;
      RECT  1.15 0.715 1.25 1.43 ;
      RECT  1.13 1.43 1.25 1.625 ;
    END
    ANTENNADIFFAREA 0.183 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.315 0.19 0.415 ;
      RECT  0.07 0.415 1.23 0.535 ;
      RECT  1.11 0.315 1.23 0.415 ;
  END
END SEN_OAI41_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI41_2
#      Description : "4-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3|A4)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI41_2
  CLASS CORE ;
  FOREIGN SEN_OAI41_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.114 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.114 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.05 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.114 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.114 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.685 3.05 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1002 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.44 0.44 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  2.5 1.44 2.63 1.75 ;
      RECT  3.02 1.41 3.145 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.57 0.05 0.7 0.345 ;
      RECT  1.16 0.05 1.29 0.345 ;
      RECT  1.75 0.05 1.88 0.345 ;
      RECT  2.27 0.05 2.4 0.36 ;
      RECT  0.055 0.05 0.18 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.39 2.885 0.56 ;
      RECT  2.75 0.56 2.85 1.23 ;
      RECT  2.32 1.23 2.935 1.35 ;
      RECT  2.32 1.35 2.41 1.44 ;
      RECT  2.01 1.44 2.41 1.56 ;
    END
    ANTENNADIFFAREA 0.288 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.505 0.21 3.145 0.3 ;
      RECT  3.025 0.3 3.145 0.43 ;
      RECT  2.505 0.3 2.625 0.45 ;
      RECT  0.265 0.435 2.16 0.45 ;
      RECT  0.265 0.45 2.625 0.55 ;
      RECT  2.14 1.015 2.49 1.135 ;
      RECT  2.14 1.135 2.23 1.24 ;
      RECT  1.8 1.24 2.23 1.33 ;
      RECT  1.8 1.33 1.92 1.44 ;
      RECT  1.255 1.44 1.92 1.56 ;
      RECT  0.895 1.02 1.265 1.14 ;
      RECT  0.895 1.14 0.985 1.23 ;
      RECT  0.055 1.23 0.985 1.35 ;
      RECT  0.055 1.35 0.175 1.61 ;
      RECT  1.075 1.24 1.71 1.35 ;
      RECT  1.075 1.35 1.165 1.465 ;
      RECT  0.785 1.465 1.165 1.585 ;
  END
END SEN_OAI41_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAI41_4
#      Description : "4-input OR into 2-input NAND"
#      Equation    : X=!((A1|A2|A3|A4)&B)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAI41_4
  CLASS CORE ;
  FOREIGN SEN_OAI41_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.71 4.05 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2277 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.64 2.85 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2277 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.64 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2277 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2277 ;
  END A4
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.35 0.51 5.45 0.71 ;
      RECT  4.75 0.71 5.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2001 ;
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.45 0.455 1.75 ;
      RECT  0.0 1.75 5.6 1.85 ;
      RECT  0.845 1.45 0.975 1.75 ;
      RECT  4.32 1.39 4.445 1.75 ;
      RECT  4.835 1.39 4.965 1.75 ;
      RECT  5.38 1.21 5.5 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      RECT  0.305 0.05 0.475 0.32 ;
      RECT  0.825 0.05 0.995 0.32 ;
      RECT  3.515 0.05 3.685 0.32 ;
      RECT  4.035 0.05 4.205 0.32 ;
      RECT  1.435 0.05 1.605 0.335 ;
      RECT  1.955 0.05 2.125 0.335 ;
      RECT  2.475 0.05 2.645 0.335 ;
      RECT  2.995 0.05 3.165 0.335 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.415 5.26 0.535 ;
      RECT  4.55 0.535 4.65 1.11 ;
      RECT  3.65 1.11 5.25 1.205 ;
      RECT  3.23 1.205 5.25 1.29 ;
      RECT  3.23 1.29 3.74 1.325 ;
    END
    ANTENNADIFFAREA 0.576 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.32 0.215 5.53 0.325 ;
      RECT  4.32 0.325 4.44 0.41 ;
      RECT  3.28 0.27 3.4 0.41 ;
      RECT  3.28 0.41 4.44 0.44 ;
      RECT  0.07 0.31 0.19 0.41 ;
      RECT  0.07 0.41 1.275 0.44 ;
      RECT  1.155 0.265 1.275 0.41 ;
      RECT  0.07 0.44 4.44 0.53 ;
      RECT  1.72 0.27 1.84 0.44 ;
      RECT  2.24 0.27 2.36 0.44 ;
      RECT  2.76 0.265 2.88 0.44 ;
      RECT  0.07 1.24 1.89 1.36 ;
      RECT  0.07 1.36 0.19 1.46 ;
      RECT  2.45 1.24 3.14 1.36 ;
      RECT  3.02 1.36 3.14 1.44 ;
      RECT  3.02 1.44 4.23 1.56 ;
      RECT  1.41 1.45 2.93 1.56 ;
  END
END SEN_OAI41_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAO211_DG_1
#      Description : "One 2-input OR into 2-input AND into 2-input OR"
#      Equation    : X=((A1|A2)&B)|C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAO211_DG_1
  CLASS CORE ;
  FOREIGN SEN_OAO211_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.635 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.635 0.45 0.87 ;
      RECT  0.35 0.87 0.56 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.72 0.635 0.85 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.635 1.05 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.35 1.39 1.48 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.32 0.05 0.45 0.365 ;
      RECT  1.1 0.05 1.23 0.365 ;
      RECT  1.35 0.05 1.48 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.735 0.69 ;
      RECT  1.55 0.69 1.65 1.11 ;
      RECT  1.55 1.11 1.735 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.21 0.185 0.455 ;
      RECT  0.065 0.455 0.705 0.545 ;
      RECT  0.585 0.21 0.705 0.455 ;
      RECT  0.845 0.21 0.965 0.455 ;
      RECT  0.845 0.455 1.245 0.545 ;
      RECT  1.155 0.545 1.245 0.785 ;
      RECT  1.155 0.785 1.45 0.895 ;
      RECT  1.155 0.895 1.245 1.37 ;
      RECT  1.105 1.37 1.245 1.54 ;
      RECT  0.39 1.26 0.965 1.35 ;
      RECT  0.39 1.35 0.49 1.39 ;
      RECT  0.845 1.35 0.965 1.565 ;
      RECT  0.065 1.39 0.49 1.48 ;
      RECT  0.065 1.48 0.185 1.61 ;
  END
END SEN_OAO211_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAO211_DG_2
#      Description : "One 2-input OR into 2-input AND into 2-input OR"
#      Equation    : X=((A1|A2)&B)|C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAO211_DG_2
  CLASS CORE ;
  FOREIGN SEN_OAO211_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.635 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.545 0.89 ;
      RECT  0.35 0.89 0.45 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.5 0.85 0.71 ;
      RECT  0.655 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.13 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.49 1.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.53 1.44 0.645 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.3 1.42 1.43 1.75 ;
      RECT  1.83 1.41 1.94 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.33 0.05 0.44 0.365 ;
      RECT  1.18 0.05 1.35 0.38 ;
      RECT  1.83 0.05 1.94 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.85 0.69 ;
      RECT  1.75 0.69 1.85 1.11 ;
      RECT  1.55 1.11 1.85 1.29 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.55 0.215 0.72 0.385 ;
      RECT  0.55 0.385 0.64 0.455 ;
      RECT  0.08 0.23 0.17 0.455 ;
      RECT  0.08 0.455 0.64 0.545 ;
      RECT  1.355 0.785 1.66 0.895 ;
      RECT  1.355 0.895 1.445 1.24 ;
      RECT  0.83 0.215 1.045 0.385 ;
      RECT  0.955 0.385 1.045 1.24 ;
      RECT  0.955 1.24 1.445 1.33 ;
      RECT  1.055 1.33 1.155 1.53 ;
      RECT  0.34 1.24 0.825 1.33 ;
      RECT  0.34 1.33 0.43 1.405 ;
      RECT  0.735 1.33 0.825 1.415 ;
      RECT  0.065 1.405 0.43 1.495 ;
      RECT  0.735 1.415 0.905 1.585 ;
      RECT  0.065 1.495 0.185 1.585 ;
  END
END SEN_OAO211_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAO211_DG_4
#      Description : "One 2-input OR into 2-input AND into 2-input OR"
#      Equation    : X=((A1|A2)&B)|C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAO211_DG_4
  CLASS CORE ;
  FOREIGN SEN_OAO211_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.635 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.545 0.925 ;
      RECT  0.35 0.925 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.655 0.71 0.85 0.925 ;
      RECT  0.75 0.925 0.85 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.635 1.05 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.355 1.21 1.46 1.75 ;
      RECT  1.875 1.41 1.995 1.75 ;
      RECT  2.395 1.21 2.515 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.32 0.05 0.45 0.365 ;
      RECT  1.1 0.05 1.23 0.365 ;
      RECT  1.87 0.05 2.0 0.39 ;
      RECT  2.395 0.05 2.515 0.59 ;
      RECT  1.355 0.05 1.46 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 2.25 0.69 ;
      RECT  2.15 0.69 2.25 1.11 ;
      RECT  1.55 1.11 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.325 0.185 0.455 ;
      RECT  0.065 0.455 0.705 0.545 ;
      RECT  0.585 0.325 0.705 0.455 ;
      RECT  0.845 0.325 0.965 0.455 ;
      RECT  0.845 0.455 1.245 0.545 ;
      RECT  1.155 0.545 1.245 0.785 ;
      RECT  1.155 0.785 2.04 0.895 ;
      RECT  1.155 0.895 1.245 1.37 ;
      RECT  1.105 1.37 1.245 1.54 ;
      RECT  0.39 1.26 0.965 1.35 ;
      RECT  0.39 1.35 0.49 1.405 ;
      RECT  0.845 1.35 0.965 1.48 ;
      RECT  0.065 1.405 0.49 1.495 ;
      RECT  0.065 1.495 0.185 1.625 ;
  END
END SEN_OAO211_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAO211_DG_8
#      Description : "One 2-input OR into 2-input AND into 2-input OR"
#      Equation    : X=((A1|A2)&B)|C
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAO211_DG_8
  CLASS CORE ;
  FOREIGN SEN_OAO211_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 2.25 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.445 0.455 1.75 ;
      RECT  0.0 1.75 5.0 1.85 ;
      RECT  1.615 1.445 1.745 1.75 ;
      RECT  2.65 1.19 2.77 1.75 ;
      RECT  3.165 1.4 3.295 1.75 ;
      RECT  3.685 1.4 3.815 1.75 ;
      RECT  4.205 1.4 4.335 1.75 ;
      RECT  4.75 1.21 4.87 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      RECT  0.585 0.05 0.715 0.35 ;
      RECT  2.135 0.05 2.265 0.355 ;
      RECT  1.105 0.05 1.23 0.36 ;
      RECT  3.165 0.05 3.295 0.4 ;
      RECT  3.685 0.05 3.815 0.4 ;
      RECT  4.205 0.05 4.335 0.4 ;
      RECT  0.07 0.05 0.19 0.59 ;
      RECT  4.75 0.05 4.87 0.59 ;
      RECT  2.65 0.05 2.77 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.91 0.51 4.65 0.69 ;
      RECT  4.08 0.69 4.25 1.11 ;
      RECT  2.91 1.11 4.65 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.32 0.245 2.0 0.355 ;
      RECT  1.88 0.355 2.0 0.445 ;
      RECT  1.88 0.445 2.515 0.555 ;
      RECT  2.405 0.555 2.515 0.785 ;
      RECT  2.405 0.785 3.985 0.895 ;
      RECT  2.405 0.895 2.505 1.245 ;
      RECT  2.09 1.245 2.505 1.355 ;
      RECT  0.28 0.45 1.79 0.56 ;
      RECT  0.07 1.245 0.705 1.355 ;
      RECT  0.595 1.355 0.705 1.445 ;
      RECT  0.07 1.355 0.19 1.465 ;
      RECT  0.595 1.445 1.28 1.555 ;
      RECT  0.8 1.245 1.995 1.355 ;
      RECT  1.885 1.355 1.995 1.445 ;
      RECT  1.885 1.445 2.56 1.555 ;
  END
END SEN_OAO211_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_12
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_12
  CLASS CORE ;
  FOREIGN SEN_OAOI211_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 13 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.605 0.75 6.055 0.87 ;
      RECT  4.475 0.75 5.135 0.87 ;
      RECT  3.55 0.75 4.025 0.87 ;
      RECT  2.485 0.75 2.935 0.87 ;
      RECT  1.455 0.75 1.985 0.87 ;
      RECT  0.41 0.75 0.935 0.87 ;
      LAYER M2 ;
      RECT  0.45 0.75 6.055 0.85 ;
      LAYER V1 ;
      RECT  5.715 0.75 5.815 0.85 ;
      RECT  5.915 0.75 6.015 0.85 ;
      RECT  4.65 0.75 4.75 0.85 ;
      RECT  4.85 0.75 4.95 0.85 ;
      RECT  3.635 0.75 3.735 0.85 ;
      RECT  3.835 0.75 3.935 0.85 ;
      RECT  2.545 0.75 2.645 0.85 ;
      RECT  2.745 0.75 2.845 0.85 ;
      RECT  1.525 0.75 1.625 0.85 ;
      RECT  1.725 0.75 1.825 0.85 ;
      RECT  0.49 0.75 0.59 0.85 ;
      RECT  0.69 0.75 0.79 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7452 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.81 6.405 0.92 ;
      RECT  6.15 0.92 6.25 1.0 ;
      RECT  0.15 0.71 0.25 1.0 ;
      RECT  0.15 1.0 6.25 1.09 ;
      RECT  1.15 0.71 1.25 1.0 ;
      RECT  2.15 0.71 2.25 1.0 ;
      RECT  3.15 0.71 3.25 1.0 ;
      RECT  4.15 0.71 4.255 1.0 ;
      RECT  5.35 0.73 5.45 1.0 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7452 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.75 0.71 9.45 0.89 ;
      RECT  7.75 0.89 7.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7452 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.93 0.71 12.85 0.89 ;
      RECT  12.75 0.89 12.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7452 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 13.0 1.85 ;
      RECT  1.08 1.495 1.25 1.75 ;
      RECT  2.12 1.495 2.29 1.75 ;
      RECT  3.16 1.495 3.33 1.75 ;
      RECT  4.2 1.495 4.37 1.75 ;
      RECT  5.24 1.495 5.41 1.75 ;
      RECT  6.28 1.495 6.45 1.75 ;
      RECT  6.81 1.495 6.98 1.75 ;
      RECT  7.33 1.495 7.5 1.75 ;
      RECT  7.85 1.495 8.02 1.75 ;
      RECT  8.39 1.455 8.52 1.75 ;
      RECT  8.91 1.455 9.04 1.75 ;
      RECT  9.41 1.455 9.54 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 13.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
      RECT  11.85 1.75 11.95 1.85 ;
      RECT  12.45 1.75 12.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 13.0 0.05 ;
      RECT  4.2 0.05 4.37 0.305 ;
      RECT  4.72 0.05 4.89 0.305 ;
      RECT  5.24 0.05 5.41 0.305 ;
      RECT  5.76 0.05 5.93 0.305 ;
      RECT  6.285 0.05 6.455 0.32 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  2.66 0.05 2.79 0.36 ;
      RECT  3.18 0.05 3.31 0.36 ;
      RECT  3.7 0.05 3.83 0.36 ;
      RECT  9.97 0.05 10.08 0.36 ;
      RECT  10.47 0.05 10.6 0.36 ;
      RECT  10.99 0.05 11.12 0.36 ;
      RECT  11.51 0.05 11.64 0.36 ;
      RECT  12.03 0.05 12.16 0.36 ;
      RECT  12.55 0.05 12.68 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 13.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
      RECT  11.85 -0.05 11.95 0.05 ;
      RECT  12.45 -0.05 12.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.15 0.16 9.88 0.19 ;
      RECT  6.545 0.19 9.88 0.32 ;
      RECT  8.15 0.32 9.88 0.36 ;
      RECT  9.63 0.36 9.88 0.45 ;
      RECT  9.63 0.45 12.935 0.62 ;
      RECT  9.63 0.62 10.8 0.69 ;
      RECT  10.55 0.69 10.8 1.11 ;
      RECT  9.97 1.11 12.66 1.29 ;
    END
    ANTENNADIFFAREA 1.812 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.35 0.395 6.235 0.45 ;
      RECT  0.275 0.45 9.54 0.58 ;
      RECT  1.88 0.58 9.54 0.62 ;
      RECT  4.35 0.62 7.65 0.64 ;
      RECT  1.88 0.62 2.06 0.65 ;
      RECT  3.35 0.62 3.45 0.85 ;
      RECT  6.15 0.64 7.65 0.7 ;
      RECT  7.95 1.115 9.88 1.2 ;
      RECT  1.95 1.2 9.88 1.235 ;
      RECT  0.535 1.235 9.88 1.365 ;
      RECT  9.63 1.365 9.88 1.4 ;
      RECT  0.535 1.365 8.25 1.405 ;
      RECT  9.63 1.4 12.05 1.44 ;
      RECT  2.51 1.405 2.89 1.45 ;
      RECT  3.51 1.405 3.89 1.45 ;
      RECT  4.71 1.405 5.09 1.45 ;
      RECT  5.71 1.405 6.09 1.45 ;
      RECT  7.645 1.405 7.745 1.49 ;
      RECT  8.15 1.405 8.25 1.49 ;
      RECT  9.63 1.44 12.935 1.63 ;
      LAYER M2 ;
      RECT  1.88 0.55 6.54 0.65 ;
      RECT  2.51 1.35 8.29 1.45 ;
      LAYER V1 ;
      RECT  1.92 0.55 2.02 0.65 ;
      RECT  3.35 0.55 3.45 0.65 ;
      RECT  6.2 0.55 6.3 0.65 ;
      RECT  6.4 0.55 6.5 0.65 ;
      RECT  2.55 1.35 2.65 1.45 ;
      RECT  2.75 1.35 2.85 1.45 ;
      RECT  3.55 1.35 3.65 1.45 ;
      RECT  3.75 1.35 3.85 1.45 ;
      RECT  4.75 1.35 4.85 1.45 ;
      RECT  4.95 1.35 5.05 1.45 ;
      RECT  5.75 1.35 5.85 1.45 ;
      RECT  5.95 1.35 6.05 1.45 ;
      RECT  7.645 1.35 7.745 1.45 ;
      RECT  8.15 1.35 8.25 1.45 ;
  END
END SEN_OAOI211_12
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_8
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_8
  CLASS CORE ;
  FOREIGN SEN_OAOI211_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.43 0.75 3.88 0.87 ;
      RECT  2.495 0.75 2.945 0.87 ;
      RECT  1.495 0.75 1.945 0.87 ;
      RECT  0.53 0.75 1.0 0.87 ;
      LAYER M2 ;
      RECT  0.56 0.75 3.855 0.85 ;
      LAYER V1 ;
      RECT  3.515 0.75 3.615 0.85 ;
      RECT  3.715 0.75 3.815 0.85 ;
      RECT  2.57 0.75 2.67 0.85 ;
      RECT  2.77 0.75 2.87 0.85 ;
      RECT  1.555 0.75 1.655 0.85 ;
      RECT  1.755 0.75 1.855 0.85 ;
      RECT  0.64 0.75 0.74 0.85 ;
      RECT  0.84 0.75 0.94 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4968 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.96 ;
      RECT  0.15 0.96 4.25 1.05 ;
      RECT  1.15 0.71 1.25 0.96 ;
      RECT  2.15 0.71 2.25 0.96 ;
      RECT  3.15 0.71 3.25 0.96 ;
      RECT  4.15 0.71 4.25 0.96 ;
      RECT  0.15 1.05 0.25 1.105 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4968 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.25 0.89 ;
      RECT  6.15 0.89 6.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4968 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 8.65 0.89 ;
      RECT  8.55 0.89 8.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4968 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  3.18 1.44 3.31 1.75 ;
      RECT  4.22 1.44 4.35 1.75 ;
      RECT  4.71 1.44 4.84 1.75 ;
      RECT  5.23 1.44 5.36 1.75 ;
      RECT  5.75 1.44 5.88 1.75 ;
      RECT  6.27 1.44 6.395 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  2.66 0.05 2.79 0.36 ;
      RECT  3.18 0.05 3.31 0.36 ;
      RECT  3.7 0.05 3.83 0.36 ;
      RECT  4.22 0.05 4.34 0.36 ;
      RECT  6.79 0.05 6.92 0.36 ;
      RECT  7.31 0.05 7.44 0.36 ;
      RECT  7.83 0.05 7.96 0.36 ;
      RECT  8.35 0.05 8.48 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.43 0.19 6.685 0.34 ;
      RECT  5.15 0.34 6.685 0.36 ;
      RECT  6.515 0.36 6.685 0.45 ;
      RECT  6.515 0.45 8.735 0.58 ;
      RECT  8.615 0.36 8.735 0.45 ;
      RECT  6.515 0.58 7.25 0.69 ;
      RECT  7.08 0.69 7.25 1.11 ;
      RECT  6.75 1.11 8.46 1.29 ;
    END
    ANTENNADIFFAREA 1.211 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.325 0.45 5.05 0.47 ;
      RECT  0.325 0.47 6.425 0.6 ;
      RECT  0.325 0.6 5.05 0.62 ;
      RECT  4.43 1.055 4.6 1.175 ;
      RECT  0.585 1.175 4.6 1.18 ;
      RECT  0.585 1.18 6.66 1.35 ;
      RECT  6.49 1.35 6.66 1.415 ;
      RECT  6.49 1.415 8.74 1.585 ;
  END
END SEN_OAOI211_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_G_8
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_G_8
  CLASS CORE ;
  FOREIGN SEN_OAOI211_G_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.43 0.75 3.88 0.895 ;
      RECT  2.495 0.75 2.945 0.895 ;
      RECT  1.495 0.75 1.945 0.895 ;
      RECT  0.425 0.75 0.915 0.895 ;
      LAYER M2 ;
      RECT  0.425 0.75 3.855 0.85 ;
      LAYER V1 ;
      RECT  3.515 0.75 3.615 0.85 ;
      RECT  3.715 0.75 3.815 0.85 ;
      RECT  2.57 0.75 2.67 0.85 ;
      RECT  2.77 0.75 2.87 0.85 ;
      RECT  1.555 0.75 1.655 0.85 ;
      RECT  1.755 0.75 1.855 0.85 ;
      RECT  0.465 0.75 0.565 0.85 ;
      RECT  0.665 0.75 0.765 0.85 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 0.985 ;
      RECT  0.15 0.985 4.25 1.075 ;
      RECT  1.15 0.71 1.25 0.985 ;
      RECT  2.15 0.71 2.25 0.985 ;
      RECT  3.15 0.71 3.25 0.985 ;
      RECT  4.15 0.71 4.25 0.985 ;
      RECT  0.15 1.075 0.25 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.25 0.89 ;
      RECT  6.15 0.89 6.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.35 0.71 8.65 0.89 ;
      RECT  8.55 0.89 8.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 8.8 1.85 ;
      RECT  1.1 1.44 1.23 1.75 ;
      RECT  2.14 1.44 2.27 1.75 ;
      RECT  3.18 1.44 3.31 1.75 ;
      RECT  4.22 1.44 4.35 1.75 ;
      RECT  4.71 1.44 4.84 1.75 ;
      RECT  5.23 1.44 5.36 1.75 ;
      RECT  5.75 1.44 5.88 1.75 ;
      RECT  6.27 1.44 6.4 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  2.66 0.05 2.79 0.36 ;
      RECT  3.18 0.05 3.31 0.36 ;
      RECT  3.7 0.05 3.83 0.36 ;
      RECT  4.22 0.05 4.34 0.36 ;
      RECT  6.79 0.05 6.92 0.36 ;
      RECT  7.31 0.05 7.44 0.36 ;
      RECT  7.83 0.05 7.96 0.36 ;
      RECT  8.35 0.05 8.48 0.36 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.43 0.19 6.685 0.34 ;
      RECT  5.15 0.34 6.685 0.36 ;
      RECT  6.515 0.36 6.685 0.45 ;
      RECT  6.515 0.45 8.735 0.58 ;
      RECT  8.615 0.36 8.735 0.45 ;
      RECT  6.515 0.58 7.25 0.69 ;
      RECT  7.08 0.69 7.25 1.11 ;
      RECT  6.75 1.11 8.46 1.29 ;
    END
    ANTENNADIFFAREA 1.293 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.325 0.45 5.05 0.47 ;
      RECT  0.325 0.47 6.425 0.6 ;
      RECT  0.325 0.6 5.05 0.62 ;
      RECT  4.43 1.06 4.6 1.175 ;
      RECT  0.585 1.175 4.6 1.18 ;
      RECT  0.585 1.18 6.66 1.35 ;
      RECT  6.49 1.35 6.66 1.415 ;
      RECT  6.49 1.415 8.74 1.585 ;
  END
END SEN_OAOI211_G_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_0P5
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_0P5
  CLASS CORE ;
  FOREIGN SEN_OAOI211_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.635 0.25 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.545 0.91 ;
      RECT  0.35 0.91 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.655 0.71 0.85 0.91 ;
      RECT  0.75 0.91 0.85 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.635 1.05 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0312 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.58 1.44 0.71 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.32 0.05 0.45 0.365 ;
      RECT  1.12 0.05 1.25 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.845 0.21 0.965 0.455 ;
      RECT  0.845 0.455 1.25 0.545 ;
      RECT  1.15 0.545 1.25 1.37 ;
      RECT  1.105 1.37 1.25 1.54 ;
    END
    ANTENNADIFFAREA 0.092 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.21 0.185 0.455 ;
      RECT  0.065 0.455 0.705 0.545 ;
      RECT  0.585 0.21 0.705 0.455 ;
      RECT  0.39 1.26 0.965 1.35 ;
      RECT  0.39 1.35 0.49 1.38 ;
      RECT  0.845 1.35 0.965 1.51 ;
      RECT  0.065 1.38 0.49 1.47 ;
      RECT  0.065 1.47 0.185 1.6 ;
  END
END SEN_OAOI211_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_1
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_1
  CLASS CORE ;
  FOREIGN SEN_OAOI211_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.64 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0621 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.55 0.905 ;
      RECT  0.35 0.905 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0621 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.655 0.71 0.85 0.905 ;
      RECT  0.75 0.905 0.85 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0621 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.635 1.05 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0621 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.585 1.44 0.715 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.325 0.05 0.455 0.365 ;
      RECT  1.125 0.05 1.255 0.365 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.85 0.325 0.97 0.455 ;
      RECT  0.85 0.455 1.25 0.545 ;
      RECT  1.15 0.545 1.25 1.37 ;
      RECT  1.105 1.37 1.25 1.54 ;
    END
    ANTENNADIFFAREA 0.182 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.325 0.19 0.455 ;
      RECT  0.07 0.455 0.71 0.545 ;
      RECT  0.59 0.325 0.71 0.455 ;
      RECT  0.395 1.26 0.97 1.35 ;
      RECT  0.395 1.35 0.495 1.39 ;
      RECT  0.85 1.35 0.97 1.51 ;
      RECT  0.07 1.39 0.495 1.48 ;
      RECT  0.07 1.48 0.19 1.61 ;
  END
END SEN_OAOI211_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_2
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_2
  CLASS CORE ;
  FOREIGN SEN_OAOI211_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1242 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1242 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1242 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1242 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.445 0.455 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.615 1.445 1.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.585 0.05 0.715 0.355 ;
      RECT  2.14 0.05 2.27 0.355 ;
      RECT  1.105 0.05 1.23 0.36 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.32 0.245 2.05 0.355 ;
      RECT  1.885 0.355 2.05 0.445 ;
      RECT  1.885 0.445 2.52 0.555 ;
      RECT  2.4 0.335 2.52 0.445 ;
      RECT  2.15 0.555 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.346 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.45 1.79 0.56 ;
      RECT  0.07 1.245 0.705 1.355 ;
      RECT  0.595 1.355 0.705 1.445 ;
      RECT  0.07 1.355 0.19 1.465 ;
      RECT  0.595 1.445 1.28 1.555 ;
      RECT  0.8 1.245 1.995 1.355 ;
      RECT  1.885 1.355 1.995 1.39 ;
      RECT  1.885 1.39 2.52 1.5 ;
      RECT  2.4 1.5 2.52 1.61 ;
  END
END SEN_OAOI211_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_3
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_3
  CLASS CORE ;
  FOREIGN SEN_OAOI211_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1863 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1863 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.14 0.71 2.45 0.9 ;
      RECT  2.35 0.9 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1863 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.25 0.905 ;
      RECT  3.15 0.905 3.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1863 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.115 1.445 1.245 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  1.645 1.445 1.775 1.75 ;
      RECT  2.165 1.445 2.295 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.325 0.05 0.455 0.355 ;
      RECT  0.845 0.05 0.975 0.355 ;
      RECT  1.385 0.05 1.515 0.355 ;
      RECT  2.685 0.05 2.815 0.365 ;
      RECT  3.21 0.05 3.33 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.86 0.455 3.12 0.565 ;
      RECT  2.75 0.565 2.85 1.245 ;
      RECT  2.64 1.245 3.33 1.355 ;
      RECT  3.21 1.355 3.33 1.51 ;
    END
    ANTENNADIFFAREA 0.474 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.65 0.245 2.34 0.355 ;
      RECT  1.65 0.355 1.77 0.445 ;
      RECT  0.07 0.335 0.19 0.445 ;
      RECT  0.07 0.445 1.77 0.555 ;
      RECT  0.655 1.055 1.845 1.145 ;
      RECT  0.655 1.145 0.745 1.245 ;
      RECT  1.755 1.145 1.845 1.245 ;
      RECT  0.07 1.245 0.745 1.355 ;
      RECT  1.755 1.245 2.545 1.355 ;
      RECT  0.07 1.355 0.19 1.465 ;
      RECT  2.435 1.355 2.545 1.445 ;
      RECT  2.435 1.445 3.12 1.555 ;
      RECT  0.855 1.245 1.56 1.355 ;
      RECT  0.855 1.355 0.965 1.445 ;
      RECT  0.28 1.445 0.965 1.555 ;
  END
END SEN_OAOI211_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_4
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_4
  CLASS CORE ;
  FOREIGN SEN_OAOI211_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2484 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2484 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2484 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2484 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.445 0.435 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.835 1.445 0.955 1.75 ;
      RECT  2.595 1.445 2.715 1.75 ;
      RECT  3.115 1.445 3.235 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.315 0.05 0.435 0.355 ;
      RECT  0.835 0.05 0.955 0.355 ;
      RECT  1.355 0.05 1.475 0.355 ;
      RECT  3.635 0.05 3.755 0.355 ;
      RECT  4.155 0.05 4.275 0.355 ;
      RECT  1.875 0.05 1.995 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.29 0.22 3.49 0.33 ;
      RECT  3.35 0.33 3.49 0.445 ;
      RECT  3.35 0.445 4.52 0.555 ;
      RECT  4.43 0.385 4.52 0.445 ;
      RECT  3.55 0.555 3.65 1.11 ;
      RECT  3.55 1.11 4.26 1.29 ;
    END
    ANTENNADIFFAREA 0.626 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.055 0.415 0.175 0.49 ;
      RECT  0.055 0.49 3.26 0.6 ;
      RECT  2.57 0.475 2.74 0.49 ;
      RECT  3.09 0.475 3.26 0.49 ;
      RECT  2.325 0.99 2.45 1.245 ;
      RECT  1.33 1.245 3.46 1.355 ;
      RECT  3.35 1.355 3.46 1.44 ;
      RECT  3.35 1.44 4.535 1.555 ;
      RECT  4.415 1.555 4.535 1.61 ;
      RECT  0.055 1.245 1.21 1.355 ;
      RECT  1.1 1.355 1.21 1.445 ;
      RECT  0.055 1.355 0.175 1.6 ;
      RECT  1.1 1.445 2.28 1.555 ;
  END
END SEN_OAOI211_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_G_1
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_G_1
  CLASS CORE ;
  FOREIGN SEN_OAOI211_G_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.64 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.55 0.925 ;
      RECT  0.35 0.925 0.45 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.655 0.71 0.85 0.925 ;
      RECT  0.75 0.925 0.85 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.645 1.05 1.17 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.58 1.44 0.715 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  1.125 0.05 1.255 0.35 ;
      RECT  0.325 0.05 0.455 0.36 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.8 0.44 1.25 0.555 ;
      RECT  1.15 0.555 1.25 1.37 ;
      RECT  1.105 1.37 1.25 1.54 ;
    END
    ANTENNADIFFAREA 0.192 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.07 0.325 0.19 0.45 ;
      RECT  0.07 0.45 0.71 0.55 ;
      RECT  0.59 0.325 0.71 0.45 ;
      RECT  0.4 1.26 0.97 1.35 ;
      RECT  0.4 1.35 0.49 1.395 ;
      RECT  0.85 1.35 0.97 1.51 ;
      RECT  0.07 1.395 0.49 1.485 ;
      RECT  0.07 1.485 0.19 1.615 ;
  END
END SEN_OAOI211_G_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_G_2
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_G_2
  CLASS CORE ;
  FOREIGN SEN_OAOI211_G_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 1.85 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.35 0.71 2.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.445 0.455 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.615 1.445 1.745 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.585 0.05 0.715 0.355 ;
      RECT  2.14 0.05 2.265 0.355 ;
      RECT  1.105 0.05 1.23 0.36 ;
      RECT  0.07 0.05 0.19 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.32 0.245 2.05 0.355 ;
      RECT  1.88 0.355 2.05 0.445 ;
      RECT  1.88 0.445 2.52 0.555 ;
      RECT  2.4 0.335 2.52 0.445 ;
      RECT  2.15 0.555 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.37 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.28 0.45 1.79 0.565 ;
      RECT  0.07 1.245 0.705 1.355 ;
      RECT  0.595 1.355 0.705 1.445 ;
      RECT  0.07 1.355 0.19 1.465 ;
      RECT  0.595 1.445 1.28 1.555 ;
      RECT  0.8 1.24 2.0 1.355 ;
      RECT  1.88 1.355 2.0 1.4 ;
      RECT  1.88 1.4 2.52 1.51 ;
      RECT  2.4 1.51 2.52 1.62 ;
  END
END SEN_OAOI211_G_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OAOI211_G_4
#      Description : "One 2-input OR into 2-input AND into 2-input NOR"
#      Equation    : X=!(((A1|A2)&B)|C)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OAOI211_G_4
  CLASS CORE ;
  FOREIGN SEN_OAOI211_G_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.705 2.05 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.05 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A2
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.65 0.89 ;
      RECT  4.55 0.89 4.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.395 1.445 0.525 1.75 ;
      RECT  0.0 1.75 4.8 1.85 ;
      RECT  0.915 1.445 1.045 1.75 ;
      RECT  2.725 1.445 2.855 1.75 ;
      RECT  3.245 1.445 3.375 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      RECT  0.655 0.05 0.785 0.355 ;
      RECT  1.175 0.05 1.305 0.355 ;
      RECT  1.695 0.05 1.825 0.355 ;
      RECT  3.765 0.05 3.895 0.355 ;
      RECT  4.285 0.05 4.415 0.355 ;
      RECT  2.215 0.05 2.34 0.36 ;
      RECT  0.12 0.05 0.24 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.43 0.245 3.65 0.355 ;
      RECT  3.51 0.355 3.65 0.445 ;
      RECT  3.51 0.445 4.72 0.555 ;
      RECT  3.75 0.555 3.85 1.11 ;
      RECT  3.75 1.11 4.45 1.29 ;
    END
    ANTENNADIFFAREA 0.682 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.35 0.45 3.42 0.56 ;
      RECT  0.09 1.245 1.295 1.355 ;
      RECT  1.185 1.355 1.295 1.445 ;
      RECT  1.185 1.445 2.39 1.555 ;
      RECT  1.39 1.245 3.625 1.355 ;
      RECT  3.515 1.355 3.625 1.445 ;
      RECT  3.515 1.445 4.72 1.555 ;
  END
END SEN_OAOI211_G_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_1
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_1
  CLASS CORE ;
  FOREIGN SEN_OR2_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.495 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.55 0.89 0.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0558 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.64 1.41 0.77 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.64 0.05 0.77 0.35 ;
      RECT  0.075 0.05 0.205 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.31 1.05 1.3 ;
    END
    ANTENNADIFFAREA 0.194 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.345 0.33 0.465 0.44 ;
      RECT  0.345 0.44 0.845 0.56 ;
      RECT  0.755 0.56 0.845 1.21 ;
      RECT  0.46 1.21 0.845 1.3 ;
      RECT  0.46 1.3 0.55 1.41 ;
      RECT  0.08 1.41 0.55 1.5 ;
      RECT  0.08 1.5 0.2 1.63 ;
  END
END SEN_OR2_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_12
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_12
  CLASS CORE ;
  FOREIGN SEN_OR2_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.615 ;
      RECT  0.35 0.615 1.85 0.715 ;
      RECT  0.35 0.715 0.45 0.895 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4572 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.31 2.65 0.51 ;
      RECT  2.55 0.51 3.595 0.69 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4572 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.68 1.45 2.79 1.75 ;
      RECT  0.0 1.75 8.2 1.85 ;
      RECT  3.18 1.45 3.31 1.75 ;
      RECT  3.7 1.41 3.83 1.75 ;
      RECT  4.22 1.41 4.35 1.75 ;
      RECT  4.745 1.21 4.865 1.75 ;
      RECT  5.26 1.41 5.39 1.75 ;
      RECT  5.78 1.41 5.91 1.75 ;
      RECT  6.32 1.41 6.45 1.75 ;
      RECT  6.88 1.41 7.01 1.75 ;
      RECT  7.44 1.41 7.57 1.75 ;
      RECT  8.0 1.21 8.12 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      RECT  0.84 0.05 0.97 0.345 ;
      RECT  1.36 0.05 1.53 0.345 ;
      RECT  3.96 0.05 4.09 0.385 ;
      RECT  0.275 0.05 0.405 0.39 ;
      RECT  3.42 0.05 3.55 0.39 ;
      RECT  4.48 0.05 4.61 0.39 ;
      RECT  5.26 0.05 5.39 0.39 ;
      RECT  5.78 0.05 5.91 0.39 ;
      RECT  6.32 0.05 6.45 0.39 ;
      RECT  6.88 0.05 7.01 0.39 ;
      RECT  7.44 0.05 7.57 0.39 ;
      RECT  4.745 0.05 4.865 0.59 ;
      RECT  7.995 0.05 8.115 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.2 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.98 0.51 7.875 0.63 ;
      RECT  5.55 0.63 7.875 0.69 ;
      RECT  7.01 0.69 7.26 1.11 ;
      RECT  5.005 1.11 7.875 1.29 ;
    END
    ANTENNADIFFAREA 1.296 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.705 0.19 3.825 0.475 ;
      RECT  3.705 0.475 4.345 0.565 ;
      RECT  4.225 0.19 4.345 0.475 ;
      RECT  4.225 0.565 4.345 0.75 ;
      RECT  4.225 0.75 5.385 0.8 ;
      RECT  0.585 0.19 0.705 0.435 ;
      RECT  0.585 0.435 2.12 0.525 ;
      RECT  1.105 0.19 1.225 0.435 ;
      RECT  2.0 0.525 2.12 0.8 ;
      RECT  2.0 0.8 6.88 0.905 ;
      RECT  2.0 0.905 5.995 1.0 ;
      RECT  2.0 1.0 4.36 1.05 ;
      RECT  2.0 1.05 2.25 1.08 ;
      RECT  1.625 1.08 2.25 1.15 ;
      RECT  0.065 1.15 2.25 1.28 ;
      RECT  0.065 1.28 0.185 1.37 ;
      RECT  2.34 1.16 4.63 1.28 ;
      RECT  2.34 1.28 3.595 1.36 ;
      RECT  2.34 1.36 2.59 1.39 ;
      RECT  0.275 1.39 2.59 1.51 ;
      RECT  1.345 1.51 2.59 1.59 ;
  END
END SEN_OR2_12
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_2
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_2
  CLASS CORE ;
  FOREIGN SEN_OR2_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0906 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0906 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.84 1.45 0.97 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.29 1.425 1.42 1.75 ;
      RECT  1.815 1.21 1.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.855 0.05 0.985 0.35 ;
      RECT  1.255 0.05 1.385 0.35 ;
      RECT  0.235 0.05 0.365 0.39 ;
      RECT  1.815 0.05 1.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.5 1.66 1.3 ;
    END
    ANTENNADIFFAREA 0.224 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.55 0.44 1.445 0.56 ;
      RECT  1.355 0.56 1.445 0.965 ;
      RECT  0.55 0.56 0.66 1.04 ;
      RECT  0.27 1.04 0.66 1.15 ;
      RECT  1.105 1.02 1.225 1.24 ;
      RECT  0.065 1.24 1.225 1.36 ;
      RECT  0.065 1.36 0.185 1.46 ;
  END
END SEN_OR2_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_3
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_3
  CLASS CORE ;
  FOREIGN SEN_OR2_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.31 0.65 0.71 ;
      RECT  0.15 0.71 0.65 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1251 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.45 0.71 ;
      RECT  1.15 0.71 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1251 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.11 1.41 1.235 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.63 1.21 1.75 1.75 ;
      RECT  2.145 1.41 2.275 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  2.07 0.05 2.2 0.39 ;
      RECT  0.24 0.05 0.36 0.57 ;
      RECT  1.13 0.05 1.25 0.59 ;
      RECT  1.54 0.05 1.66 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 2.45 0.69 ;
      RECT  2.35 0.69 2.45 1.11 ;
      RECT  1.9 1.11 2.53 1.29 ;
    END
    ANTENNADIFFAREA 0.394 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.715 0.79 2.24 0.895 ;
      RECT  1.715 0.895 1.805 1.01 ;
      RECT  0.85 0.315 0.97 1.01 ;
      RECT  0.75 1.01 1.805 1.1 ;
      RECT  0.75 1.1 0.84 1.21 ;
      RECT  0.07 1.21 0.84 1.33 ;
      RECT  0.07 1.33 0.19 1.43 ;
      RECT  0.93 1.21 1.515 1.32 ;
      RECT  0.93 1.32 1.02 1.42 ;
      RECT  0.33 1.42 1.02 1.53 ;
      RECT  0.33 1.53 0.45 1.63 ;
  END
END SEN_OR2_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_4
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_4
  CLASS CORE ;
  FOREIGN SEN_OR2_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.49 0.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1596 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.655 0.89 ;
      RECT  1.35 0.89 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1596 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.125 1.41 1.255 1.75 ;
      RECT  0.0 1.75 3.0 1.85 ;
      RECT  1.715 1.21 1.835 1.75 ;
      RECT  2.29 1.41 2.42 1.75 ;
      RECT  2.815 1.21 2.935 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      RECT  0.235 0.05 0.365 0.39 ;
      RECT  0.865 0.05 0.995 0.39 ;
      RECT  1.125 0.05 1.255 0.39 ;
      RECT  1.71 0.05 1.84 0.39 ;
      RECT  2.29 0.05 2.42 0.39 ;
      RECT  2.815 0.05 2.935 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.01 0.51 2.66 0.69 ;
      RECT  2.55 0.69 2.66 1.11 ;
      RECT  1.95 1.11 2.66 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.61 0.19 0.73 0.5 ;
      RECT  0.61 0.5 1.905 0.59 ;
      RECT  1.39 0.19 1.51 0.5 ;
      RECT  1.815 0.59 1.905 0.79 ;
      RECT  0.61 0.59 0.73 1.21 ;
      RECT  1.815 0.79 2.44 0.89 ;
      RECT  0.09 1.21 0.73 1.3 ;
      RECT  0.09 1.3 0.21 1.43 ;
      RECT  0.87 1.21 1.56 1.31 ;
      RECT  0.87 1.31 0.99 1.39 ;
      RECT  0.35 1.39 0.99 1.49 ;
      RECT  0.35 1.49 0.47 1.61 ;
  END
END SEN_OR2_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_6
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_6
  CLASS CORE ;
  FOREIGN SEN_OR2_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.31 0.45 0.5 ;
      RECT  0.35 0.5 0.85 0.69 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2286 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.295 1.85 0.51 ;
      RECT  1.75 0.51 2.25 0.69 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2286 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.62 1.45 1.75 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  2.14 1.45 2.27 1.75 ;
      RECT  2.665 1.21 2.785 1.75 ;
      RECT  3.18 1.4 3.31 1.75 ;
      RECT  3.7 1.4 3.83 1.75 ;
      RECT  4.22 1.41 4.345 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  0.82 0.05 0.95 0.39 ;
      RECT  1.38 0.05 1.51 0.39 ;
      RECT  2.12 0.05 2.25 0.39 ;
      RECT  3.18 0.05 3.31 0.39 ;
      RECT  3.7 0.05 3.83 0.39 ;
      RECT  2.66 0.05 2.79 0.395 ;
      RECT  4.22 0.05 4.345 0.395 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.92 0.51 4.25 0.69 ;
      RECT  3.92 0.69 4.05 1.11 ;
      RECT  2.92 1.11 4.25 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.405 0.195 2.525 0.795 ;
      RECT  2.405 0.795 3.83 0.895 ;
      RECT  2.405 0.895 2.525 1.01 ;
      RECT  1.1 0.195 1.22 1.01 ;
      RECT  1.1 1.01 2.525 1.1 ;
      RECT  1.1 1.1 1.22 1.21 ;
      RECT  0.06 1.21 1.22 1.32 ;
      RECT  0.06 1.32 0.18 1.59 ;
      RECT  1.365 1.24 2.55 1.36 ;
      RECT  1.365 1.36 1.485 1.44 ;
      RECT  0.295 1.44 1.485 1.56 ;
  END
END SEN_OR2_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_8
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_8
  CLASS CORE ;
  FOREIGN SEN_OR2_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.31 2.05 0.51 ;
      RECT  1.95 0.51 2.755 0.69 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3024 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.51 1.45 0.69 ;
      RECT  1.35 0.69 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3024 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.325 1.255 0.445 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  0.845 1.255 0.965 1.75 ;
      RECT  1.365 1.255 1.485 1.75 ;
      RECT  3.435 1.21 3.555 1.75 ;
      RECT  3.95 1.41 4.08 1.75 ;
      RECT  4.47 1.41 4.6 1.75 ;
      RECT  5.015 1.41 5.145 1.75 ;
      RECT  5.59 1.21 5.71 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  0.625 0.05 0.795 0.24 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  2.64 0.05 2.77 0.39 ;
      RECT  3.95 0.05 4.08 0.39 ;
      RECT  4.47 0.05 4.6 0.39 ;
      RECT  5.015 0.05 5.145 0.39 ;
      RECT  3.34 0.05 3.46 0.59 ;
      RECT  5.59 0.05 5.71 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.695 0.51 5.46 0.69 ;
      RECT  5.09 0.69 5.26 1.11 ;
      RECT  3.695 1.11 5.46 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.925 0.22 3.045 0.79 ;
      RECT  2.925 0.79 4.93 0.91 ;
      RECT  2.925 0.91 4.275 0.96 ;
      RECT  2.925 0.96 3.095 1.2 ;
      RECT  0.325 0.2 0.445 0.33 ;
      RECT  0.325 0.33 1.77 0.42 ;
      RECT  1.65 0.42 1.77 0.79 ;
      RECT  1.65 0.79 2.0 0.895 ;
      RECT  1.885 0.895 2.0 1.2 ;
      RECT  1.885 1.2 3.095 1.35 ;
      RECT  0.065 1.01 1.77 1.16 ;
      RECT  0.065 1.16 0.185 1.23 ;
      RECT  1.6 1.16 1.77 1.44 ;
      RECT  1.6 1.44 3.33 1.59 ;
  END
END SEN_OR2_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_DG_1
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_DG_1
  CLASS CORE ;
  FOREIGN SEN_OR2_DG_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.305 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.525 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0279 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.635 1.39 0.765 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.615 0.05 0.785 0.345 ;
      RECT  0.075 0.05 0.205 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.45 1.05 1.29 ;
    END
    ANTENNADIFFAREA 0.189 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.2 0.46 0.435 ;
      RECT  0.34 0.435 0.72 0.545 ;
      RECT  0.63 0.545 0.72 0.755 ;
      RECT  0.63 0.755 0.86 0.925 ;
      RECT  0.63 0.925 0.72 1.19 ;
      RECT  0.385 1.19 0.72 1.295 ;
      RECT  0.385 1.295 0.485 1.395 ;
      RECT  0.08 1.395 0.485 1.515 ;
      RECT  0.08 1.515 0.2 1.615 ;
  END
END SEN_OR2_DG_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_DG_2
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_DG_2
  CLASS CORE ;
  FOREIGN SEN_OR2_DG_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.305 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.525 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.605 1.42 0.785 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.2 1.21 1.32 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.575 0.05 0.745 0.345 ;
      RECT  1.175 0.05 1.345 0.345 ;
      RECT  0.055 0.05 0.225 0.355 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.915 0.51 1.25 0.69 ;
      RECT  1.15 0.69 1.25 1.0 ;
      RECT  0.95 1.0 1.25 1.1 ;
      RECT  0.95 1.1 1.05 1.3 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.26 0.46 0.435 ;
      RECT  0.34 0.435 0.72 0.545 ;
      RECT  0.63 0.545 0.72 0.795 ;
      RECT  0.63 0.795 1.04 0.885 ;
      RECT  0.63 0.885 0.72 1.205 ;
      RECT  0.385 1.205 0.72 1.31 ;
      RECT  0.385 1.31 0.485 1.41 ;
      RECT  0.08 1.41 0.485 1.53 ;
      RECT  0.08 1.53 0.2 1.63 ;
  END
END SEN_OR2_DG_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_DG_3
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_DG_3
  CLASS CORE ;
  FOREIGN SEN_OR2_DG_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.305 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.505 0.89 ;
      RECT  0.35 0.89 0.45 1.12 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.048 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.585 1.44 0.755 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.14 1.24 1.31 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.55 0.05 0.72 0.345 ;
      RECT  0.055 0.05 0.2 0.37 ;
      RECT  1.16 0.05 1.29 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.88 0.51 1.545 0.69 ;
      RECT  1.35 0.69 1.45 1.015 ;
      RECT  1.35 1.015 1.54 1.05 ;
      RECT  0.88 1.05 1.54 1.15 ;
      RECT  1.425 1.15 1.54 1.19 ;
    END
    ANTENNADIFFAREA 0.356 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.265 0.435 0.685 0.545 ;
      RECT  0.595 0.545 0.685 0.795 ;
      RECT  0.595 0.795 1.24 0.885 ;
      RECT  0.595 0.885 0.685 1.25 ;
      RECT  0.35 1.25 0.685 1.34 ;
      RECT  0.35 1.34 0.44 1.395 ;
      RECT  0.055 1.395 0.44 1.485 ;
      RECT  0.055 1.485 0.175 1.615 ;
  END
END SEN_OR2_DG_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_DG_4
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_DG_4
  CLASS CORE ;
  FOREIGN SEN_OR2_DG_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.14 0.71 0.255 1.305 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.52 0.925 ;
      RECT  0.35 0.925 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.57 1.405 0.7 1.75 ;
      RECT  0.0 1.75 1.8 1.85 ;
      RECT  1.095 1.25 1.215 1.75 ;
      RECT  1.61 1.41 1.74 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      RECT  0.55 0.05 0.72 0.345 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  1.61 0.05 1.74 0.39 ;
      RECT  1.09 0.05 1.22 0.41 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.81 0.51 1.65 0.69 ;
      RECT  1.55 0.69 1.65 1.04 ;
      RECT  0.835 1.04 1.65 1.16 ;
      RECT  0.835 1.16 0.955 1.27 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.265 0.435 0.72 0.545 ;
      RECT  0.63 0.545 0.72 0.79 ;
      RECT  0.63 0.79 1.44 0.89 ;
      RECT  0.63 0.89 0.72 1.21 ;
      RECT  0.36 1.21 0.72 1.315 ;
      RECT  0.36 1.315 0.47 1.395 ;
      RECT  0.055 1.395 0.47 1.505 ;
      RECT  0.055 1.505 0.175 1.615 ;
  END
END SEN_OR2_DG_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_DG_6
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_DG_6
  CLASS CORE ;
  FOREIGN SEN_OR2_DG_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.725 0.71 0.945 0.905 ;
      RECT  0.725 0.905 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.71 0.49 0.905 ;
      RECT  0.145 0.905 0.265 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.096 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.31 1.39 0.44 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.515 1.245 1.685 1.75 ;
      RECT  2.035 1.24 2.205 1.75 ;
      RECT  2.555 1.24 2.725 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.55 0.05 0.72 0.345 ;
      RECT  1.215 0.05 1.345 0.37 ;
      RECT  1.8 0.05 1.92 0.385 ;
      RECT  2.32 0.05 2.44 0.385 ;
      RECT  0.055 0.05 0.18 0.39 ;
      RECT  2.87 0.05 2.99 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.495 0.51 2.725 0.69 ;
      RECT  2.52 0.69 2.65 1.05 ;
      RECT  1.235 1.05 3.01 1.15 ;
    END
    ANTENNADIFFAREA 0.702 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.265 0.435 1.145 0.545 ;
      RECT  1.05 0.545 1.145 0.79 ;
      RECT  1.05 0.79 2.405 0.89 ;
      RECT  1.05 0.89 1.145 1.24 ;
      RECT  0.785 1.24 1.145 1.36 ;
      RECT  0.055 1.18 0.695 1.28 ;
      RECT  0.055 1.28 0.175 1.375 ;
      RECT  0.575 1.28 0.695 1.465 ;
      RECT  0.575 1.465 1.265 1.585 ;
  END
END SEN_OR2_DG_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_DG_8
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_DG_8
  CLASS CORE ;
  FOREIGN SEN_OR2_DG_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.73 0.71 0.985 0.905 ;
      RECT  0.73 0.905 0.85 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.14 0.71 0.535 0.905 ;
      RECT  0.14 0.905 0.26 1.11 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.315 1.44 0.485 1.75 ;
      RECT  0.0 1.75 3.6 1.85 ;
      RECT  1.57 1.245 1.74 1.75 ;
      RECT  2.09 1.24 2.26 1.75 ;
      RECT  2.61 1.24 2.78 1.75 ;
      RECT  3.13 1.24 3.3 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      RECT  1.095 0.05 1.265 0.34 ;
      RECT  0.575 0.05 0.745 0.355 ;
      RECT  3.13 0.05 3.3 0.375 ;
      RECT  1.575 0.05 1.725 0.385 ;
      RECT  2.09 0.05 2.26 0.385 ;
      RECT  2.61 0.05 2.78 0.39 ;
      RECT  0.08 0.05 0.2 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.31 0.51 3.535 0.69 ;
      RECT  2.88 0.69 3.05 1.025 ;
      RECT  2.88 1.025 3.535 1.04 ;
      RECT  1.295 1.04 3.535 1.15 ;
      RECT  3.415 1.15 3.535 1.245 ;
    END
    ANTENNADIFFAREA 0.968 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.29 0.445 1.205 0.555 ;
      RECT  1.11 0.555 1.205 0.79 ;
      RECT  1.11 0.79 2.735 0.89 ;
      RECT  1.11 0.89 1.205 1.24 ;
      RECT  0.81 1.24 1.205 1.36 ;
      RECT  0.08 1.25 0.72 1.35 ;
      RECT  0.6 1.35 0.72 1.465 ;
      RECT  0.08 1.35 0.2 1.47 ;
      RECT  0.6 1.465 1.29 1.585 ;
  END
END SEN_OR2_DG_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_10
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_10
  CLASS CORE ;
  FOREIGN SEN_OR2_10 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.71 ;
      RECT  0.15 0.71 1.69 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5256 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.51 2.85 0.71 ;
      RECT  2.75 0.71 4.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5256 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.66 1.27 2.83 1.75 ;
      RECT  0.0 1.75 7.6 1.85 ;
      RECT  3.18 1.27 3.35 1.75 ;
      RECT  3.7 1.27 3.87 1.75 ;
      RECT  4.22 1.27 4.39 1.75 ;
      RECT  4.74 1.27 4.91 1.75 ;
      RECT  5.26 1.27 5.43 1.75 ;
      RECT  5.78 1.27 5.95 1.75 ;
      RECT  6.3 1.27 6.47 1.75 ;
      RECT  6.82 1.27 6.99 1.75 ;
      RECT  7.385 1.21 7.505 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      RECT  2.165 0.05 2.335 0.325 ;
      RECT  4.22 0.05 4.39 0.335 ;
      RECT  0.57 0.05 0.745 0.34 ;
      RECT  1.095 0.05 1.265 0.345 ;
      RECT  1.615 0.05 1.785 0.345 ;
      RECT  3.18 0.05 3.35 0.35 ;
      RECT  3.7 0.05 3.87 0.35 ;
      RECT  4.76 0.05 4.89 0.4 ;
      RECT  5.28 0.05 5.41 0.4 ;
      RECT  5.8 0.05 5.93 0.4 ;
      RECT  6.32 0.05 6.45 0.4 ;
      RECT  6.84 0.05 6.97 0.4 ;
      RECT  7.385 0.05 7.505 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  5.01 0.51 7.25 0.69 ;
      RECT  6.83 0.69 7.05 1.02 ;
      RECT  4.975 1.02 7.275 1.18 ;
    END
    ANTENNADIFFAREA 1.08 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.43 0.145 3.08 0.315 ;
      RECT  2.43 0.315 2.6 0.415 ;
      RECT  2.94 0.315 3.08 0.445 ;
      RECT  1.885 0.415 2.6 0.445 ;
      RECT  0.34 0.365 0.46 0.445 ;
      RECT  0.34 0.445 2.6 0.585 ;
      RECT  2.94 0.445 4.64 0.585 ;
      RECT  2.135 0.585 2.305 1.015 ;
      RECT  4.49 0.585 4.64 0.785 ;
      RECT  4.49 0.785 6.675 0.915 ;
      RECT  0.08 1.015 2.305 1.165 ;
      RECT  0.08 1.165 0.2 1.235 ;
      RECT  2.41 1.02 4.675 1.18 ;
      RECT  2.41 1.18 2.56 1.425 ;
      RECT  0.29 1.425 2.56 1.575 ;
  END
END SEN_OR2_10
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_16
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_16
  CLASS CORE ;
  FOREIGN SEN_OR2_16 0 0 ;
  ORIGIN 0 0 ;
  SIZE 12.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.51 0.25 0.71 ;
      RECT  0.145 0.71 3.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8856 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.51 4.25 0.71 ;
      RECT  4.15 0.71 7.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.8856 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  4.19 1.27 4.36 1.75 ;
      RECT  0.0 1.75 12.2 1.85 ;
      RECT  4.71 1.27 4.88 1.75 ;
      RECT  5.23 1.27 5.4 1.75 ;
      RECT  5.75 1.27 5.92 1.75 ;
      RECT  6.27 1.27 6.44 1.75 ;
      RECT  6.79 1.27 6.96 1.75 ;
      RECT  7.31 1.27 7.48 1.75 ;
      RECT  7.83 1.27 8.0 1.75 ;
      RECT  8.35 1.27 8.52 1.75 ;
      RECT  8.87 1.27 9.04 1.75 ;
      RECT  9.39 1.27 9.56 1.75 ;
      RECT  9.91 1.27 10.08 1.75 ;
      RECT  10.43 1.27 10.6 1.75 ;
      RECT  10.95 1.27 11.12 1.75 ;
      RECT  11.47 1.27 11.64 1.75 ;
      RECT  12.01 1.41 12.14 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 12.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 12.2 0.05 ;
      RECT  5.23 0.05 5.4 0.335 ;
      RECT  5.75 0.05 5.92 0.335 ;
      RECT  6.27 0.05 6.44 0.335 ;
      RECT  6.79 0.05 6.96 0.335 ;
      RECT  7.31 0.05 7.48 0.335 ;
      RECT  0.56 0.05 0.71 0.345 ;
      RECT  1.07 0.05 1.24 0.345 ;
      RECT  1.59 0.05 1.76 0.345 ;
      RECT  2.11 0.05 2.28 0.345 ;
      RECT  2.63 0.05 2.8 0.345 ;
      RECT  3.15 0.05 3.32 0.35 ;
      RECT  4.67 0.05 4.84 0.35 ;
      RECT  12.01 0.05 12.14 0.39 ;
      RECT  8.37 0.05 8.5 0.4 ;
      RECT  8.89 0.05 9.02 0.4 ;
      RECT  9.41 0.05 9.54 0.4 ;
      RECT  9.93 0.05 10.06 0.4 ;
      RECT  10.45 0.05 10.58 0.4 ;
      RECT  10.97 0.05 11.1 0.4 ;
      RECT  11.49 0.05 11.62 0.4 ;
      RECT  7.855 0.05 7.975 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 12.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  8.1 0.505 11.875 0.69 ;
      RECT  10.525 0.69 10.85 1.02 ;
      RECT  8.09 1.02 11.925 1.18 ;
    END
    ANTENNADIFFAREA 1.728 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.42 0.14 4.58 0.28 ;
      RECT  4.44 0.28 4.58 0.44 ;
      RECT  3.42 0.28 3.57 0.45 ;
      RECT  4.44 0.44 7.73 0.58 ;
      RECT  0.315 0.2 0.46 0.385 ;
      RECT  0.37 0.385 0.46 0.45 ;
      RECT  0.37 0.45 3.57 0.585 ;
      RECT  7.58 0.58 7.73 0.785 ;
      RECT  3.42 0.585 3.57 1.015 ;
      RECT  7.58 0.785 10.39 0.895 ;
      RECT  0.06 1.015 3.85 1.165 ;
      RECT  0.06 1.165 0.175 1.21 ;
      RECT  3.94 1.02 7.745 1.18 ;
      RECT  3.94 1.18 4.09 1.425 ;
      RECT  0.265 1.425 4.09 1.575 ;
  END
END SEN_OR2_16
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_1P5
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_1P5
  CLASS CORE ;
  FOREIGN SEN_OR2_1P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.084 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.945 0.505 1.05 0.705 ;
      RECT  0.945 0.705 1.25 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.084 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.85 1.27 1.02 1.75 ;
      RECT  0.0 1.75 2.2 1.85 ;
      RECT  1.395 1.215 1.515 1.75 ;
      RECT  1.935 1.225 2.055 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      RECT  0.825 0.05 0.995 0.185 ;
      RECT  1.37 0.05 1.54 0.335 ;
      RECT  0.31 0.05 0.485 0.34 ;
      RECT  1.93 0.05 2.06 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.655 0.29 1.775 0.51 ;
      RECT  1.655 0.51 2.05 0.69 ;
      RECT  1.95 0.69 2.05 1.045 ;
      RECT  1.66 1.045 2.05 1.135 ;
      RECT  1.66 1.135 1.77 1.345 ;
    END
    ANTENNADIFFAREA 0.162 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.6 0.275 1.255 0.375 ;
      RECT  0.6 0.375 0.725 0.445 ;
      RECT  1.14 0.375 1.255 0.445 ;
      RECT  0.08 0.26 0.2 0.445 ;
      RECT  0.08 0.445 0.725 0.535 ;
      RECT  1.14 0.445 1.48 0.535 ;
      RECT  0.35 0.535 0.725 0.54 ;
      RECT  1.39 0.535 1.48 0.81 ;
      RECT  0.35 0.54 0.45 1.315 ;
      RECT  1.39 0.81 1.74 0.92 ;
      RECT  0.6 1.05 1.25 1.15 ;
      RECT  1.14 1.15 1.25 1.385 ;
      RECT  0.6 1.15 0.72 1.405 ;
      RECT  0.08 1.405 0.72 1.515 ;
      RECT  0.08 1.515 0.2 1.625 ;
  END
END SEN_OR2_1P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_24
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_24
  CLASS CORE ;
  FOREIGN SEN_OR2_24 0 0 ;
  ORIGIN 0 0 ;
  SIZE 17.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.145 0.51 0.25 0.71 ;
      RECT  0.145 0.71 4.31 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3104 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.75 0.705 10.45 0.905 ;
      RECT  10.35 0.905 10.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.3104 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  5.75 1.285 5.92 1.75 ;
      RECT  0.0 1.75 17.4 1.85 ;
      RECT  6.27 1.285 6.44 1.75 ;
      RECT  6.79 1.285 6.96 1.75 ;
      RECT  7.31 1.285 7.48 1.75 ;
      RECT  7.83 1.285 8.0 1.75 ;
      RECT  8.35 1.285 8.52 1.75 ;
      RECT  8.87 1.285 9.04 1.75 ;
      RECT  9.39 1.285 9.56 1.75 ;
      RECT  9.93 1.45 10.06 1.75 ;
      RECT  10.45 1.45 10.58 1.75 ;
      RECT  10.975 1.19 11.095 1.75 ;
      RECT  11.495 1.4 11.625 1.75 ;
      RECT  12.015 1.4 12.145 1.75 ;
      RECT  12.535 1.4 12.665 1.75 ;
      RECT  13.055 1.4 13.185 1.75 ;
      RECT  13.575 1.4 13.705 1.75 ;
      RECT  14.095 1.4 14.225 1.75 ;
      RECT  14.615 1.4 14.745 1.75 ;
      RECT  15.135 1.4 15.265 1.75 ;
      RECT  15.655 1.4 15.785 1.75 ;
      RECT  16.175 1.4 16.305 1.75 ;
      RECT  16.695 1.4 16.825 1.75 ;
      RECT  17.215 1.41 17.34 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 17.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
      RECT  9.25 1.75 9.35 1.85 ;
      RECT  9.85 1.75 9.95 1.85 ;
      RECT  10.45 1.75 10.55 1.85 ;
      RECT  11.05 1.75 11.15 1.85 ;
      RECT  11.65 1.75 11.75 1.85 ;
      RECT  12.25 1.75 12.35 1.85 ;
      RECT  12.85 1.75 12.95 1.85 ;
      RECT  13.45 1.75 13.55 1.85 ;
      RECT  14.05 1.75 14.15 1.85 ;
      RECT  14.65 1.75 14.75 1.85 ;
      RECT  15.25 1.75 15.35 1.85 ;
      RECT  15.85 1.75 15.95 1.85 ;
      RECT  16.45 1.75 16.55 1.85 ;
      RECT  17.05 1.75 17.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 17.4 0.05 ;
      RECT  6.27 0.05 6.44 0.335 ;
      RECT  6.79 0.05 6.96 0.335 ;
      RECT  7.31 0.05 7.48 0.335 ;
      RECT  7.83 0.05 8.0 0.335 ;
      RECT  8.35 0.05 8.52 0.335 ;
      RECT  8.87 0.05 9.04 0.335 ;
      RECT  9.39 0.05 9.56 0.335 ;
      RECT  9.91 0.05 10.08 0.335 ;
      RECT  10.43 0.05 10.6 0.34 ;
      RECT  12.515 0.05 12.685 0.345 ;
      RECT  14.075 0.05 14.245 0.345 ;
      RECT  14.595 0.05 14.765 0.345 ;
      RECT  15.115 0.05 15.285 0.345 ;
      RECT  15.635 0.05 15.805 0.345 ;
      RECT  16.155 0.05 16.325 0.345 ;
      RECT  16.675 0.05 16.845 0.345 ;
      RECT  0.81 0.05 0.98 0.35 ;
      RECT  1.33 0.05 1.5 0.35 ;
      RECT  1.85 0.05 2.02 0.35 ;
      RECT  2.37 0.05 2.54 0.35 ;
      RECT  2.89 0.05 3.06 0.35 ;
      RECT  3.41 0.05 3.58 0.35 ;
      RECT  3.93 0.05 4.1 0.35 ;
      RECT  4.45 0.05 4.62 0.35 ;
      RECT  4.97 0.05 5.14 0.35 ;
      RECT  5.62 0.05 5.79 0.35 ;
      RECT  11.475 0.05 11.645 0.35 ;
      RECT  13.555 0.05 13.725 0.35 ;
      RECT  11.995 0.05 12.165 0.355 ;
      RECT  13.035 0.05 13.205 0.355 ;
      RECT  0.285 0.05 0.415 0.39 ;
      RECT  17.215 0.05 17.34 0.39 ;
      RECT  10.98 0.05 11.09 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 17.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
      RECT  9.25 -0.05 9.35 0.05 ;
      RECT  9.85 -0.05 9.95 0.05 ;
      RECT  10.45 -0.05 10.55 0.05 ;
      RECT  11.05 -0.05 11.15 0.05 ;
      RECT  11.65 -0.05 11.75 0.05 ;
      RECT  12.25 -0.05 12.35 0.05 ;
      RECT  12.85 -0.05 12.95 0.05 ;
      RECT  13.45 -0.05 13.55 0.05 ;
      RECT  14.05 -0.05 14.15 0.05 ;
      RECT  14.65 -0.05 14.75 0.05 ;
      RECT  15.25 -0.05 15.35 0.05 ;
      RECT  15.85 -0.05 15.95 0.05 ;
      RECT  16.45 -0.05 16.55 0.05 ;
      RECT  17.05 -0.05 17.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  11.215 0.455 17.13 0.57 ;
      RECT  11.215 0.57 16.65 0.625 ;
      RECT  13.305 0.625 15.05 0.69 ;
      RECT  13.95 0.69 14.45 1.055 ;
      RECT  13.35 1.055 17.095 1.11 ;
      RECT  11.215 1.11 17.095 1.29 ;
    END
    ANTENNADIFFAREA 2.592 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.56 0.44 10.85 0.615 ;
      RECT  0.56 0.615 4.87 0.62 ;
      RECT  10.655 0.615 10.85 0.735 ;
      RECT  4.61 0.62 4.87 1.015 ;
      RECT  10.655 0.735 13.14 0.78 ;
      RECT  10.655 0.78 13.38 0.895 ;
      RECT  0.055 1.015 5.365 1.21 ;
      RECT  15.23 0.75 16.855 0.895 ;
      RECT  5.455 1.0 9.845 1.195 ;
      RECT  9.745 1.195 9.845 1.24 ;
      RECT  5.455 1.195 5.65 1.405 ;
      RECT  9.745 1.24 10.86 1.36 ;
      RECT  0.275 1.405 5.65 1.6 ;
      LAYER M2 ;
      RECT  12.76 0.75 15.645 0.85 ;
      LAYER V1 ;
      RECT  12.8 0.75 12.9 0.85 ;
      RECT  13.0 0.75 13.1 0.85 ;
      RECT  15.27 0.75 15.37 0.85 ;
      RECT  15.495 0.75 15.595 0.85 ;
  END
END SEN_OR2_24
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_2P5
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_2P5
  CLASS CORE ;
  FOREIGN SEN_OR2_2P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.495 0.25 0.705 ;
      RECT  0.15 0.705 0.505 0.91 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1404 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.505 1.25 0.705 ;
      RECT  1.15 0.705 1.48 0.71 ;
      RECT  0.95 0.71 1.48 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1404 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.095 1.27 1.265 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.64 1.21 1.76 1.75 ;
      RECT  2.155 1.41 2.285 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.07 0.05 1.24 0.19 ;
      RECT  0.55 0.05 0.725 0.345 ;
      RECT  1.615 0.05 1.785 0.35 ;
      RECT  2.135 0.05 2.305 0.35 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.42 0.205 2.535 0.445 ;
      RECT  1.85 0.445 2.535 0.555 ;
      RECT  2.35 0.555 2.45 1.11 ;
      RECT  1.905 1.11 2.45 1.115 ;
      RECT  1.905 1.115 2.535 1.29 ;
    END
    ANTENNADIFFAREA 0.3 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.28 1.5 0.37 ;
      RECT  0.845 0.37 0.955 0.435 ;
      RECT  1.375 0.37 1.5 0.45 ;
      RECT  0.32 0.205 0.455 0.4 ;
      RECT  0.365 0.4 0.455 0.435 ;
      RECT  0.365 0.435 0.955 0.535 ;
      RECT  1.375 0.45 1.725 0.54 ;
      RECT  0.63 0.535 0.725 1.135 ;
      RECT  1.63 0.54 1.725 0.78 ;
      RECT  1.63 0.78 2.25 0.89 ;
      RECT  0.06 1.135 0.725 1.235 ;
      RECT  0.06 1.235 0.18 1.34 ;
      RECT  0.865 1.07 1.495 1.16 ;
      RECT  1.385 1.16 1.495 1.35 ;
      RECT  0.865 1.16 0.975 1.445 ;
      RECT  0.27 1.445 0.975 1.555 ;
  END
END SEN_OR2_2P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OR2_5
#      Description : "2-Input OR"
#      Equation    : X=A1|A2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR2_5
  CLASS CORE ;
  FOREIGN SEN_OR2_5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 0.705 ;
      RECT  0.15 0.705 0.98 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2805 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.505 1.85 0.71 ;
      RECT  1.75 0.71 2.505 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2805 ;
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.66 1.26 1.83 1.75 ;
      RECT  0.0 1.75 4.2 1.85 ;
      RECT  2.18 1.26 2.35 1.75 ;
      RECT  2.7 1.26 2.87 1.75 ;
      RECT  3.22 1.27 3.39 1.75 ;
      RECT  3.74 1.27 3.91 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      RECT  1.635 0.05 1.805 0.215 ;
      RECT  2.18 0.05 2.35 0.365 ;
      RECT  0.595 0.05 0.725 0.38 ;
      RECT  1.115 0.05 1.245 0.385 ;
      RECT  2.72 0.05 2.85 0.39 ;
      RECT  3.24 0.05 3.37 0.39 ;
      RECT  3.76 0.05 3.89 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.505 4.145 0.69 ;
      RECT  3.94 0.69 4.05 1.0 ;
      RECT  3.94 1.0 4.145 1.065 ;
      RECT  2.935 1.065 4.145 1.18 ;
    END
    ANTENNADIFFAREA 0.574 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.38 0.315 2.065 0.415 ;
      RECT  1.38 0.415 1.49 0.475 ;
      RECT  1.94 0.415 2.065 0.485 ;
      RECT  0.345 0.29 0.455 0.475 ;
      RECT  0.345 0.475 1.49 0.585 ;
      RECT  1.94 0.485 2.735 0.605 ;
      RECT  1.135 0.585 1.265 1.04 ;
      RECT  2.625 0.605 2.735 0.785 ;
      RECT  2.625 0.785 3.77 0.895 ;
      RECT  0.08 1.04 1.265 1.155 ;
      RECT  0.08 1.155 0.2 1.26 ;
      RECT  1.38 1.04 2.635 1.16 ;
      RECT  1.38 1.16 1.5 1.44 ;
      RECT  0.29 1.44 1.5 1.56 ;
  END
END SEN_OR2_5
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3_1
#      Description : "3-Input OR"
#      Equation    : X=A1|A2|A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3_1
  CLASS CORE ;
  FOREIGN SEN_OR3_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.65 0.89 ;
      RECT  0.35 0.89 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.74 0.51 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.865 1.41 0.995 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.31 0.05 0.48 0.21 ;
      RECT  0.85 0.05 1.02 0.21 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.3 0.69 ;
      RECT  1.15 0.69 1.25 1.29 ;
    END
    ANTENNADIFFAREA 0.173 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.2 0.185 0.3 ;
      RECT  0.065 0.3 1.06 0.42 ;
      RECT  0.97 0.42 1.06 1.21 ;
      RECT  0.625 1.21 1.06 1.3 ;
      RECT  0.625 1.3 0.725 1.41 ;
      RECT  0.065 1.41 0.725 1.51 ;
      RECT  0.065 1.51 0.185 1.63 ;
  END
END SEN_OR3_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3_2
#      Description : "3-Input OR"
#      Equation    : X=A1|A2|A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3_2
  CLASS CORE ;
  FOREIGN SEN_OR3_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.51 1.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.36 1.415 1.475 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.885 1.21 2.005 1.75 ;
      RECT  2.405 1.21 2.525 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  0.57 0.05 0.74 0.21 ;
      RECT  1.125 0.05 1.295 0.21 ;
      RECT  2.4 0.05 2.53 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  1.86 0.05 1.98 0.605 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.5 2.45 0.69 ;
      RECT  2.35 0.69 2.45 1.0 ;
      RECT  2.15 1.0 2.45 1.1 ;
      RECT  2.15 1.1 2.25 1.3 ;
    END
    ANTENNADIFFAREA 0.216 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.29 0.3 1.77 0.42 ;
      RECT  1.68 0.42 1.77 0.785 ;
      RECT  0.55 0.42 0.65 1.21 ;
      RECT  1.68 0.785 2.26 0.895 ;
      RECT  0.285 1.21 0.65 1.33 ;
      RECT  0.81 1.21 1.775 1.32 ;
      RECT  0.065 1.34 0.185 1.44 ;
      RECT  0.065 1.44 1.27 1.56 ;
  END
END SEN_OR3_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3_4
#      Description : "3-Input OR"
#      Equation    : X=A1|A2|A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3_4
  CLASS CORE ;
  FOREIGN SEN_OR3_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2253 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2253 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 2.65 0.71 ;
      RECT  2.55 0.71 3.05 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2253 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.28 1.22 2.52 1.325 ;
      RECT  2.42 1.325 2.52 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  2.85 1.255 2.97 1.75 ;
      RECT  3.37 1.21 3.49 1.75 ;
      RECT  3.885 1.44 4.015 1.75 ;
      RECT  4.41 1.21 4.53 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  2.715 0.05 2.845 0.24 ;
      RECT  3.885 0.05 4.015 0.35 ;
      RECT  0.46 0.05 0.59 0.375 ;
      RECT  1.17 0.05 1.3 0.375 ;
      RECT  1.82 0.05 1.95 0.375 ;
      RECT  3.37 0.05 3.49 0.59 ;
      RECT  4.41 0.05 4.53 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.6 0.51 4.255 0.69 ;
      RECT  4.15 0.69 4.255 1.11 ;
      RECT  3.63 1.11 4.255 1.29 ;
    END
    ANTENNADIFFAREA 0.432 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.145 0.33 3.28 0.42 ;
      RECT  2.145 0.42 2.26 0.47 ;
      RECT  3.16 0.42 3.28 0.785 ;
      RECT  0.065 0.37 0.185 0.47 ;
      RECT  0.065 0.47 2.26 0.59 ;
      RECT  0.955 0.59 1.045 1.23 ;
      RECT  3.16 0.785 4.04 0.895 ;
      RECT  0.285 1.23 1.045 1.35 ;
      RECT  2.03 1.01 3.27 1.13 ;
      RECT  2.03 1.13 2.13 1.205 ;
      RECT  1.34 1.205 2.13 1.31 ;
      RECT  0.065 1.36 0.185 1.465 ;
      RECT  0.065 1.465 2.31 1.585 ;
  END
END SEN_OR3_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3_6
#      Description : "3-Input OR"
#      Equation    : X=A1|A2|A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3_6
  CLASS CORE ;
  FOREIGN SEN_OR3_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 1.05 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3276 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.64 2.65 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3276 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.35 0.64 4.05 0.89 ;
      RECT  3.35 0.89 3.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3276 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  3.17 1.435 3.3 1.75 ;
      RECT  0.0 1.75 6.4 1.85 ;
      RECT  3.69 1.435 3.82 1.75 ;
      RECT  4.43 1.21 4.55 1.75 ;
      RECT  5.095 1.405 5.225 1.75 ;
      RECT  5.615 1.405 5.745 1.75 ;
      RECT  6.17 1.21 6.29 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 6.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      RECT  1.85 0.05 2.02 0.305 ;
      RECT  2.37 0.05 2.54 0.305 ;
      RECT  2.89 0.05 3.06 0.305 ;
      RECT  3.41 0.05 3.58 0.305 ;
      RECT  3.93 0.05 4.1 0.305 ;
      RECT  0.57 0.05 0.7 0.36 ;
      RECT  1.16 0.05 1.29 0.36 ;
      RECT  0.05 0.05 0.18 0.39 ;
      RECT  5.095 0.05 5.225 0.39 ;
      RECT  5.615 0.05 5.745 0.39 ;
      RECT  4.52 0.05 4.64 0.57 ;
      RECT  6.18 0.05 6.3 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 6.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.51 6.05 0.69 ;
      RECT  5.92 0.69 6.05 1.11 ;
      RECT  4.75 1.11 6.05 1.29 ;
    END
    ANTENNADIFFAREA 0.648 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.4 0.395 4.375 0.45 ;
      RECT  0.275 0.45 4.375 0.525 ;
      RECT  0.275 0.525 1.53 0.57 ;
      RECT  4.245 0.525 4.375 0.785 ;
      RECT  1.4 0.57 1.53 1.215 ;
      RECT  4.245 0.785 5.81 0.895 ;
      RECT  0.29 1.215 1.53 1.345 ;
      RECT  1.82 1.215 4.13 1.345 ;
      RECT  0.055 1.37 0.175 1.445 ;
      RECT  0.055 1.445 2.83 1.575 ;
  END
END SEN_OR3_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3_3
#      Description : "3-Input OR"
#      Equation    : X=A1|A2|A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3_3
  CLASS CORE ;
  FOREIGN SEN_OR3_3 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.65 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1656 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.45 0.89 ;
      RECT  0.95 0.89 1.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1656 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.7 2.05 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1656 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.88 1.42 2.01 1.75 ;
      RECT  0.0 1.75 3.4 1.85 ;
      RECT  2.405 1.19 2.525 1.75 ;
      RECT  2.92 1.41 3.05 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.4 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      RECT  0.82 0.05 0.99 0.315 ;
      RECT  1.34 0.05 1.51 0.315 ;
      RECT  0.3 0.05 0.47 0.32 ;
      RECT  1.87 0.05 2.04 0.32 ;
      RECT  2.92 0.05 3.05 0.39 ;
      RECT  2.405 0.05 2.525 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.4 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.665 0.51 3.305 0.69 ;
      RECT  3.15 0.69 3.25 1.11 ;
      RECT  2.665 1.11 3.305 1.29 ;
    END
    ANTENNADIFFAREA 0.389 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.305 0.185 0.41 ;
      RECT  0.065 0.41 2.275 0.525 ;
      RECT  2.155 0.325 2.275 0.41 ;
      RECT  2.155 0.525 2.275 0.78 ;
      RECT  0.755 0.525 0.845 1.245 ;
      RECT  2.155 0.78 3.06 0.9 ;
      RECT  0.065 1.245 0.845 1.355 ;
      RECT  0.065 1.355 0.185 1.465 ;
      RECT  1.055 1.21 2.315 1.33 ;
      RECT  0.275 1.455 1.535 1.575 ;
  END
END SEN_OR3_3
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3_8
#      Description : "3-Input OR"
#      Equation    : X=A1|A2|A3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3_8
  CLASS CORE ;
  FOREIGN SEN_OR3_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 1.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.64 3.45 0.89 ;
      RECT  2.15 0.89 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.55 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4482 ;
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  3.95 1.44 4.08 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  4.47 1.44 4.6 1.75 ;
      RECT  4.99 1.44 5.12 1.75 ;
      RECT  5.51 1.44 5.64 1.75 ;
      RECT  6.035 1.19 6.155 1.75 ;
      RECT  6.55 1.41 6.68 1.75 ;
      RECT  7.07 1.41 7.2 1.75 ;
      RECT  7.59 1.41 7.72 1.75 ;
      RECT  8.14 1.21 8.26 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  2.12 0.05 2.29 0.31 ;
      RECT  2.64 0.05 2.81 0.31 ;
      RECT  3.16 0.05 3.33 0.31 ;
      RECT  3.68 0.05 3.85 0.31 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.755 0.36 ;
      RECT  4.22 0.05 4.35 0.36 ;
      RECT  4.47 0.05 4.6 0.36 ;
      RECT  4.99 0.05 5.12 0.36 ;
      RECT  5.51 0.05 5.64 0.36 ;
      RECT  6.55 0.05 6.68 0.39 ;
      RECT  7.07 0.05 7.2 0.39 ;
      RECT  7.59 0.05 7.72 0.39 ;
      RECT  0.065 0.05 0.185 0.59 ;
      RECT  8.14 0.05 8.26 0.59 ;
      RECT  6.035 0.05 6.155 0.61 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  6.295 0.51 8.05 0.69 ;
      RECT  7.675 0.69 7.85 1.11 ;
      RECT  6.295 1.11 8.05 1.29 ;
    END
    ANTENNADIFFAREA 0.864 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.885 0.24 2.005 0.4 ;
      RECT  1.885 0.4 4.085 0.45 ;
      RECT  2.405 0.24 2.525 0.4 ;
      RECT  2.925 0.24 3.045 0.4 ;
      RECT  3.445 0.24 3.565 0.4 ;
      RECT  3.965 0.21 4.085 0.4 ;
      RECT  0.275 0.45 5.92 0.53 ;
      RECT  0.275 0.53 1.99 0.57 ;
      RECT  3.705 0.53 5.92 0.57 ;
      RECT  1.82 0.57 1.99 1.0 ;
      RECT  5.81 0.57 5.92 0.79 ;
      RECT  5.81 0.79 7.565 0.895 ;
      RECT  0.34 1.0 1.99 1.17 ;
      RECT  2.355 1.0 4.205 1.17 ;
      RECT  4.035 1.17 4.205 1.18 ;
      RECT  4.035 1.18 5.945 1.35 ;
      RECT  0.065 1.315 3.825 1.485 ;
  END
END SEN_OR3_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3B_0P5
#      Description : "3-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3B_0P5
  CLASS CORE ;
  FOREIGN SEN_OR3B_0P5 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.51 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0324 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.545 0.51 0.655 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0234 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.61 1.39 0.74 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.2 1.54 1.33 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.085 0.05 0.215 0.39 ;
      RECT  0.61 0.05 0.74 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.19 1.28 0.41 ;
      RECT  1.15 0.41 1.25 1.36 ;
      RECT  0.9 1.36 1.25 1.45 ;
      RECT  0.9 1.45 1.02 1.58 ;
    END
    ANTENNADIFFAREA 0.108 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.355 0.19 0.475 0.385 ;
      RECT  0.355 0.385 0.455 1.18 ;
      RECT  0.355 1.18 1.06 1.27 ;
      RECT  0.96 0.81 1.06 1.18 ;
      RECT  0.355 1.27 0.455 1.39 ;
      RECT  0.095 1.39 0.455 1.49 ;
      RECT  0.095 1.49 0.215 1.61 ;
  END
END SEN_OR3B_0P5
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3B_1
#      Description : "3-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3B_1
  CLASS CORE ;
  FOREIGN SEN_OR3B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.7 0.65 0.925 ;
      RECT  0.55 0.925 0.65 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  0.0 1.75 1.4 1.85 ;
      RECT  1.195 1.41 1.325 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.58 0.05 0.71 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.31 1.25 0.6 ;
      RECT  1.15 0.6 1.345 0.69 ;
      RECT  1.245 0.69 1.345 1.11 ;
      RECT  0.95 1.11 1.345 1.29 ;
    END
    ANTENNADIFFAREA 0.255 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.34 0.345 0.445 0.5 ;
      RECT  0.34 0.5 1.04 0.59 ;
      RECT  0.94 0.59 1.04 0.785 ;
      RECT  0.34 0.59 0.43 1.41 ;
      RECT  0.94 0.785 1.14 0.895 ;
      RECT  0.065 1.41 0.43 1.53 ;
      RECT  0.065 1.53 0.185 1.63 ;
  END
END SEN_OR3B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3B_12
#      Description : "3-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3B_12
  CLASS CORE ;
  FOREIGN SEN_OR3B_12 0 0 ;
  ORIGIN 0 0 ;
  SIZE 10 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.71 9.65 0.78 ;
      RECT  6.965 0.78 9.65 0.895 ;
      RECT  9.55 0.895 9.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7776 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 0.695 ;
      RECT  0.15 0.695 1.345 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.381 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.95 0.71 3.25 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.381 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.99 1.455 2.12 1.75 ;
      RECT  0.0 1.75 10.0 1.85 ;
      RECT  2.51 1.455 2.64 1.75 ;
      RECT  3.03 1.455 3.16 1.75 ;
      RECT  3.55 1.41 3.68 1.75 ;
      RECT  4.07 1.41 4.2 1.75 ;
      RECT  4.59 1.41 4.72 1.75 ;
      RECT  5.11 1.41 5.24 1.75 ;
      RECT  5.63 1.41 5.76 1.75 ;
      RECT  6.15 1.43 6.28 1.75 ;
      RECT  6.67 1.43 6.8 1.75 ;
      RECT  7.19 1.41 7.32 1.75 ;
      RECT  7.71 1.41 7.84 1.75 ;
      RECT  8.23 1.41 8.36 1.75 ;
      RECT  8.75 1.41 8.88 1.75 ;
      RECT  9.27 1.41 9.4 1.75 ;
      RECT  9.805 1.21 9.925 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 10.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 10.0 0.05 ;
      RECT  0.69 0.05 0.82 0.345 ;
      RECT  1.21 0.05 1.34 0.345 ;
      RECT  1.73 0.05 1.86 0.345 ;
      RECT  2.25 0.05 2.38 0.345 ;
      RECT  2.77 0.05 2.9 0.345 ;
      RECT  3.29 0.05 3.415 0.345 ;
      RECT  6.945 0.05 7.06 0.345 ;
      RECT  7.45 0.05 7.58 0.345 ;
      RECT  7.97 0.05 8.1 0.345 ;
      RECT  8.49 0.05 8.62 0.345 ;
      RECT  9.01 0.05 9.14 0.345 ;
      RECT  9.53 0.05 9.66 0.345 ;
      RECT  0.145 0.05 0.275 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 10.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.765 0.51 6.05 0.535 ;
      RECT  3.765 0.535 6.535 0.69 ;
      RECT  5.385 0.69 6.535 0.73 ;
      RECT  5.855 0.73 6.535 0.77 ;
      RECT  6.285 0.77 6.535 1.11 ;
      RECT  3.75 1.11 9.45 1.18 ;
      RECT  3.75 1.18 9.705 1.29 ;
      RECT  5.855 1.29 7.09 1.34 ;
    END
    ANTENNADIFFAREA 2.016 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.505 0.19 6.855 0.325 ;
      RECT  5.075 0.325 6.855 0.345 ;
      RECT  5.595 0.345 6.855 0.39 ;
      RECT  6.115 0.39 6.855 0.425 ;
      RECT  6.625 0.425 6.855 0.435 ;
      RECT  6.625 0.435 9.915 0.555 ;
      RECT  9.795 0.335 9.915 0.435 ;
      RECT  6.625 0.555 8.9 0.585 ;
      RECT  6.625 0.585 7.875 0.635 ;
      RECT  6.625 0.635 7.355 0.665 ;
      RECT  0.385 0.435 3.675 0.555 ;
      RECT  1.365 0.555 3.675 0.585 ;
      RECT  3.525 0.585 3.675 0.785 ;
      RECT  1.47 0.585 1.62 1.215 ;
      RECT  3.525 0.785 5.1 0.82 ;
      RECT  3.525 0.82 5.765 0.86 ;
      RECT  3.525 0.86 6.065 0.95 ;
      RECT  0.385 1.215 1.62 1.34 ;
      RECT  1.735 1.235 3.465 1.365 ;
      RECT  1.735 1.365 1.865 1.46 ;
      RECT  0.125 1.46 1.865 1.59 ;
  END
END SEN_OR3B_12
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3B_2
#      Description : "3-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3B_2
  CLASS CORE ;
  FOREIGN SEN_OR3B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.71 2.45 0.89 ;
      RECT  2.35 0.89 2.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 2.6 1.85 ;
      RECT  1.355 1.2 1.46 1.75 ;
      RECT  1.87 1.41 2.0 1.75 ;
      RECT  2.4 1.21 2.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.6 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      RECT  1.08 0.05 1.25 0.335 ;
      RECT  0.58 0.05 0.71 0.345 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  2.135 0.05 2.265 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.6 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.72 0.69 ;
      RECT  1.55 0.69 1.65 1.11 ;
      RECT  1.55 1.11 2.25 1.29 ;
    END
    ANTENNADIFFAREA 0.34 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.355 0.2 1.475 0.305 ;
      RECT  1.355 0.305 1.995 0.395 ;
      RECT  1.875 0.395 1.995 0.48 ;
      RECT  1.875 0.48 2.52 0.59 ;
      RECT  2.4 0.37 2.52 0.48 ;
      RECT  0.285 0.435 1.25 0.54 ;
      RECT  1.16 0.54 1.25 0.79 ;
      RECT  1.16 0.79 1.46 0.9 ;
      RECT  1.16 0.9 1.25 1.24 ;
      RECT  0.805 1.24 1.25 1.36 ;
      RECT  0.065 1.21 0.705 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.585 1.3 0.705 1.45 ;
      RECT  0.585 1.45 1.25 1.57 ;
  END
END SEN_OR3B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3B_4
#      Description : "3-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3B_4
  CLASS CORE ;
  FOREIGN SEN_OR3B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.86 0.71 4.45 0.89 ;
      RECT  4.35 0.89 4.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2139 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2139 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 4.6 1.85 ;
      RECT  0.84 1.41 0.97 1.75 ;
      RECT  2.345 0.99 2.47 1.75 ;
      RECT  2.865 1.415 2.985 1.75 ;
      RECT  3.385 1.415 3.505 1.75 ;
      RECT  3.905 1.415 4.025 1.75 ;
      RECT  4.425 1.4 4.545 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      RECT  0.58 0.05 0.71 0.345 ;
      RECT  1.1 0.05 1.23 0.345 ;
      RECT  1.62 0.05 1.75 0.345 ;
      RECT  2.14 0.05 2.255 0.345 ;
      RECT  3.64 0.05 3.77 0.38 ;
      RECT  4.16 0.05 4.29 0.38 ;
      RECT  0.06 0.05 0.19 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.605 0.51 3.25 0.69 ;
      RECT  3.15 0.69 3.25 1.11 ;
      RECT  2.605 1.11 4.26 1.29 ;
      RECT  4.15 1.29 4.285 1.49 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.345 0.275 3.505 0.395 ;
      RECT  3.385 0.395 3.505 0.47 ;
      RECT  2.345 0.395 2.465 0.685 ;
      RECT  3.385 0.47 4.545 0.59 ;
      RECT  4.425 0.19 4.545 0.47 ;
      RECT  0.285 0.435 2.24 0.54 ;
      RECT  2.15 0.54 2.24 0.785 ;
      RECT  2.15 0.785 3.04 0.895 ;
      RECT  2.15 0.895 2.24 1.21 ;
      RECT  1.325 1.21 2.24 1.315 ;
      RECT  0.065 1.21 1.225 1.32 ;
      RECT  0.065 1.32 0.185 1.43 ;
      RECT  1.105 1.32 1.225 1.48 ;
      RECT  1.105 1.48 2.255 1.59 ;
      RECT  2.145 1.405 2.255 1.48 ;
  END
END SEN_OR3B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OR3B_8
#      Description : "3-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR3B_8
  CLASS CORE ;
  FOREIGN SEN_OR3B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.51 0.45 0.71 ;
      RECT  0.35 0.71 1.05 0.905 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.258 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.45 0.9 ;
      RECT  1.55 0.9 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.258 ;
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.615 1.44 1.745 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  2.135 1.44 2.265 1.75 ;
      RECT  2.655 1.41 2.785 1.75 ;
      RECT  3.175 1.41 3.305 1.75 ;
      RECT  3.695 1.41 3.825 1.75 ;
      RECT  4.215 1.41 4.345 1.75 ;
      RECT  4.735 1.41 4.865 1.75 ;
      RECT  5.255 1.41 5.385 1.75 ;
      RECT  5.775 1.41 5.905 1.75 ;
      RECT  6.295 1.45 6.425 1.75 ;
      RECT  6.815 1.41 6.94 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  4.995 0.05 5.125 0.36 ;
      RECT  1.095 0.05 1.225 0.38 ;
      RECT  1.615 0.05 1.745 0.38 ;
      RECT  2.235 0.05 2.365 0.38 ;
      RECT  5.515 0.05 5.645 0.39 ;
      RECT  6.035 0.05 6.165 0.39 ;
      RECT  6.555 0.05 6.685 0.39 ;
      RECT  0.56 0.05 0.68 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.87 0.51 4.625 0.63 ;
      RECT  2.87 0.63 4.51 0.69 ;
      RECT  4.34 0.69 4.51 1.11 ;
      RECT  2.75 1.11 6.25 1.245 ;
      RECT  2.75 1.245 6.73 1.29 ;
      RECT  6.145 1.29 6.73 1.36 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.61 0.215 4.885 0.335 ;
      RECT  4.19 0.335 4.885 0.365 ;
      RECT  4.735 0.365 4.885 0.45 ;
      RECT  4.735 0.45 5.43 0.48 ;
      RECT  4.735 0.48 6.945 0.6 ;
      RECT  6.82 0.2 6.945 0.48 ;
      RECT  0.79 0.47 2.75 0.59 ;
      RECT  2.63 0.59 2.75 0.78 ;
      RECT  1.145 0.59 1.255 1.225 ;
      RECT  2.63 0.78 4.23 0.895 ;
      RECT  0.06 1.225 1.255 1.345 ;
      RECT  0.06 1.345 0.18 1.61 ;
      RECT  1.36 1.22 2.57 1.34 ;
      RECT  1.36 1.34 1.48 1.435 ;
      RECT  0.27 1.435 1.48 1.56 ;
  END
END SEN_OR3B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4_1
#      Description : "4-Input OR"
#      Equation    : X=A1|A2|A3|A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4_1
  CLASS CORE ;
  FOREIGN SEN_OR4_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.51 0.91 ;
      RECT  0.35 0.91 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.51 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0534 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.665 1.41 0.795 1.75 ;
      RECT  0.0 1.75 2.0 1.85 ;
      RECT  1.285 1.41 1.415 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  0.58 0.05 0.71 0.39 ;
      RECT  1.285 0.05 1.415 0.39 ;
      RECT  1.805 0.05 1.935 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.78 0.495 1.05 0.675 ;
      RECT  0.95 0.675 1.05 1.44 ;
      RECT  0.95 1.44 1.175 1.56 ;
    END
    ANTENNADIFFAREA 0.183 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.325 0.31 0.445 0.5 ;
      RECT  0.325 0.5 0.69 0.59 ;
      RECT  0.6 0.59 0.69 0.765 ;
      RECT  0.6 0.765 0.855 0.935 ;
      RECT  0.6 0.935 0.69 1.21 ;
      RECT  0.355 1.21 0.69 1.3 ;
      RECT  0.355 1.3 0.445 1.41 ;
      RECT  0.065 1.41 0.445 1.5 ;
      RECT  0.065 1.5 0.185 1.63 ;
      RECT  1.55 0.31 1.66 0.5 ;
      RECT  1.145 0.5 1.66 0.59 ;
      RECT  1.145 0.59 1.245 1.21 ;
      RECT  1.145 1.21 1.93 1.3 ;
      RECT  1.81 1.3 1.93 1.43 ;
  END
END SEN_OR4_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4_2
#      Description : "4-Input OR"
#      Equation    : X=A1|A2|A3|A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4_2
  CLASS CORE ;
  FOREIGN SEN_OR4_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  3.75 0.89 3.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1068 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.41 0.45 1.75 ;
      RECT  0.0 1.75 4.0 1.85 ;
      RECT  1.615 1.41 1.745 1.75 ;
      RECT  2.195 1.41 2.325 1.75 ;
      RECT  3.535 1.41 3.665 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      RECT  0.555 0.05 0.735 0.34 ;
      RECT  1.075 0.05 1.255 0.34 ;
      RECT  2.72 0.05 2.9 0.34 ;
      RECT  3.25 0.05 3.43 0.34 ;
      RECT  2.2 0.05 2.32 0.36 ;
      RECT  0.06 0.05 0.19 0.385 ;
      RECT  3.795 0.05 3.925 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.51 1.85 0.69 ;
      RECT  1.75 0.69 1.85 1.11 ;
      RECT  1.35 1.11 2.65 1.29 ;
    END
    ANTENNADIFFAREA 0.477 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.355 0.2 2.06 0.29 ;
      RECT  1.355 0.29 1.475 0.42 ;
      RECT  1.94 0.29 2.06 0.45 ;
      RECT  1.94 0.45 2.61 0.57 ;
      RECT  0.3 0.43 1.25 0.53 ;
      RECT  1.155 0.53 1.25 0.785 ;
      RECT  1.155 0.785 1.64 0.895 ;
      RECT  1.155 0.895 1.25 1.21 ;
      RECT  0.79 1.21 1.25 1.33 ;
      RECT  2.76 0.43 3.71 0.53 ;
      RECT  2.76 0.53 2.85 0.785 ;
      RECT  2.15 0.785 2.85 0.895 ;
      RECT  2.75 0.895 2.85 1.21 ;
      RECT  2.75 1.21 3.165 1.33 ;
      RECT  0.065 1.21 0.7 1.3 ;
      RECT  0.065 1.3 0.185 1.43 ;
      RECT  0.585 1.3 0.7 1.44 ;
      RECT  0.585 1.44 1.28 1.56 ;
      RECT  3.28 1.21 3.92 1.3 ;
      RECT  3.8 1.3 3.92 1.43 ;
      RECT  3.28 1.3 3.4 1.45 ;
      RECT  2.71 1.45 3.4 1.56 ;
  END
END SEN_OR4_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4_4
#      Description : "4-Input OR"
#      Equation    : X=A1|A2|A3|A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4_4
  CLASS CORE ;
  FOREIGN SEN_OR4_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.85 0.89 ;
      RECT  1.35 0.89 1.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2139 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.35 0.89 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2139 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.15 0.71 5.65 0.89 ;
      RECT  5.55 0.89 5.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2139 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.15 0.71 6.65 0.89 ;
      RECT  6.55 0.89 6.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2139 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.32 1.42 0.45 1.75 ;
      RECT  0.0 1.75 7.0 1.85 ;
      RECT  0.84 1.42 0.97 1.75 ;
      RECT  2.395 1.21 2.515 1.75 ;
      RECT  2.91 1.41 3.04 1.75 ;
      RECT  3.43 1.41 3.56 1.75 ;
      RECT  3.95 1.41 4.08 1.75 ;
      RECT  4.475 1.21 4.595 1.75 ;
      RECT  6.02 1.42 6.15 1.75 ;
      RECT  6.54 1.42 6.67 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.0 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      RECT  0.84 0.05 0.97 0.38 ;
      RECT  1.36 0.05 1.49 0.38 ;
      RECT  1.935 0.05 2.065 0.38 ;
      RECT  3.69 0.05 3.82 0.38 ;
      RECT  4.21 0.05 4.34 0.38 ;
      RECT  4.94 0.05 5.06 0.38 ;
      RECT  5.5 0.05 5.63 0.38 ;
      RECT  6.02 0.05 6.15 0.38 ;
      RECT  6.64 0.05 6.76 0.39 ;
      RECT  0.24 0.05 0.36 0.585 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.0 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.51 3.32 0.69 ;
      RECT  3.15 0.69 3.32 1.11 ;
      RECT  2.63 1.11 4.36 1.29 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.395 0.2 3.56 0.32 ;
      RECT  2.395 0.32 2.515 0.39 ;
      RECT  3.43 0.32 3.56 0.47 ;
      RECT  3.43 0.47 4.62 0.59 ;
      RECT  0.53 0.47 2.25 0.59 ;
      RECT  2.15 0.59 2.25 0.785 ;
      RECT  2.15 0.785 3.06 0.895 ;
      RECT  2.15 0.895 2.25 1.21 ;
      RECT  1.34 1.21 2.25 1.33 ;
      RECT  4.75 0.47 6.46 0.59 ;
      RECT  4.75 0.59 4.85 0.79 ;
      RECT  3.74 0.79 4.85 0.89 ;
      RECT  4.75 0.89 4.85 1.21 ;
      RECT  4.75 1.21 5.675 1.33 ;
      RECT  0.065 1.21 1.225 1.33 ;
      RECT  0.065 1.33 0.185 1.43 ;
      RECT  1.105 1.33 1.225 1.48 ;
      RECT  1.105 1.48 2.265 1.6 ;
      RECT  2.145 1.43 2.265 1.48 ;
      RECT  5.765 1.21 6.925 1.33 ;
      RECT  6.805 1.33 6.925 1.45 ;
      RECT  5.765 1.33 5.885 1.48 ;
      RECT  4.725 1.43 4.845 1.48 ;
      RECT  4.725 1.48 5.885 1.6 ;
  END
END SEN_OR4_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4_6
#      Description : "4-Input OR"
#      Equation    : X=A1|A2|A3|A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4_6
  CLASS CORE ;
  FOREIGN SEN_OR4_6 0 0 ;
  ORIGIN 0 0 ;
  SIZE 9 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.45 0.89 ;
      RECT  1.75 0.89 1.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.55 0.71 1.25 0.89 ;
      RECT  1.15 0.89 1.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.71 7.25 0.89 ;
      RECT  6.75 0.89 6.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  7.95 0.71 8.45 0.89 ;
      RECT  8.35 0.89 8.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 9.0 1.85 ;
      RECT  0.58 1.415 0.71 1.75 ;
      RECT  1.1 1.415 1.23 1.75 ;
      RECT  2.915 1.21 3.035 1.75 ;
      RECT  3.43 1.41 3.56 1.75 ;
      RECT  3.95 1.41 4.08 1.75 ;
      RECT  4.47 1.41 4.6 1.75 ;
      RECT  4.99 1.41 5.12 1.75 ;
      RECT  5.51 1.41 5.64 1.75 ;
      RECT  6.03 1.41 6.16 1.75 ;
      RECT  7.775 1.415 7.905 1.75 ;
      RECT  8.295 1.415 8.425 1.75 ;
      RECT  8.815 1.41 8.94 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 9.0 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
      RECT  8.65 1.75 8.75 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  1.1 0.05 1.23 0.36 ;
      RECT  1.62 0.05 1.75 0.36 ;
      RECT  2.14 0.05 2.27 0.36 ;
      RECT  2.66 0.05 2.79 0.36 ;
      RECT  6.215 0.05 6.345 0.36 ;
      RECT  6.735 0.05 6.865 0.36 ;
      RECT  7.255 0.05 7.385 0.36 ;
      RECT  7.775 0.05 7.905 0.36 ;
      RECT  8.295 0.05 8.425 0.36 ;
      RECT  8.815 0.05 8.94 0.39 ;
      RECT  4.73 0.05 4.86 0.41 ;
      RECT  5.25 0.05 5.38 0.41 ;
      RECT  5.77 0.05 5.9 0.41 ;
      RECT  0.065 0.05 0.185 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 9.0 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
      RECT  8.65 -0.05 8.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.15 0.51 4.32 0.69 ;
      RECT  4.12 0.69 4.25 1.11 ;
      RECT  3.15 1.11 5.895 1.29 ;
      RECT  3.15 1.29 3.26 1.49 ;
      RECT  3.75 1.29 3.85 1.49 ;
      RECT  4.75 1.29 4.85 1.49 ;
      RECT  5.75 1.29 5.895 1.49 ;
    END
    ANTENNADIFFAREA 1.008 ;
  END X
  OBS
      LAYER M1 ;
      RECT  2.915 0.215 4.595 0.345 ;
      RECT  2.915 0.345 3.035 0.43 ;
      RECT  4.465 0.345 4.595 0.545 ;
      RECT  4.465 0.545 6.155 0.675 ;
      RECT  6.035 0.48 6.155 0.545 ;
      RECT  0.275 0.46 2.785 0.58 ;
      RECT  2.665 0.58 2.785 0.785 ;
      RECT  2.665 0.785 4.02 0.895 ;
      RECT  2.665 0.895 2.785 1.19 ;
      RECT  1.6 1.19 2.785 1.31 ;
      RECT  6.245 0.46 8.73 0.58 ;
      RECT  6.245 0.58 6.34 0.785 ;
      RECT  4.945 0.785 6.34 0.895 ;
      RECT  6.22 0.895 6.34 1.205 ;
      RECT  6.22 1.205 7.43 1.325 ;
      RECT  7.52 1.195 8.73 1.315 ;
      RECT  7.52 1.315 7.64 1.435 ;
      RECT  6.43 1.435 7.64 1.555 ;
      RECT  0.275 1.205 1.485 1.325 ;
      RECT  1.365 1.325 1.485 1.43 ;
      RECT  1.365 1.43 2.575 1.55 ;
  END
END SEN_OR4_6
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4_8
#      Description : "4-Input OR"
#      Equation    : X=A1|A2|A3|A4
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4_8
  CLASS CORE ;
  FOREIGN SEN_OR4_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 11.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.655 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.396 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.675 1.65 0.89 ;
      RECT  0.75 0.89 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.396 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  8.55 0.67 9.45 0.89 ;
      RECT  8.55 0.89 8.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.396 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  10.35 0.71 11.65 0.89 ;
      RECT  11.55 0.89 11.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.396 ;
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.345 1.43 0.475 1.75 ;
      RECT  0.0 1.75 11.8 1.85 ;
      RECT  0.865 1.43 0.995 1.75 ;
      RECT  1.385 1.43 1.515 1.75 ;
      RECT  3.41 0.99 3.52 1.75 ;
      RECT  3.91 1.41 4.04 1.75 ;
      RECT  4.43 1.41 4.56 1.75 ;
      RECT  4.95 1.41 5.08 1.75 ;
      RECT  5.47 1.41 5.6 1.75 ;
      RECT  5.99 1.41 6.12 1.75 ;
      RECT  6.51 1.41 6.64 1.75 ;
      RECT  7.03 1.41 7.16 1.75 ;
      RECT  7.55 1.41 7.68 1.75 ;
      RECT  9.895 1.255 10.015 1.75 ;
      RECT  10.415 1.255 10.535 1.75 ;
      RECT  10.935 1.255 11.055 1.75 ;
      RECT  11.48 1.21 11.6 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 11.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
      RECT  5.85 1.75 5.95 1.85 ;
      RECT  6.45 1.75 6.55 1.85 ;
      RECT  7.05 1.75 7.15 1.85 ;
      RECT  7.65 1.75 7.75 1.85 ;
      RECT  8.25 1.75 8.35 1.85 ;
      RECT  8.85 1.75 8.95 1.85 ;
      RECT  9.45 1.75 9.55 1.85 ;
      RECT  10.05 1.75 10.15 1.85 ;
      RECT  10.65 1.75 10.75 1.85 ;
      RECT  11.25 1.75 11.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 11.8 0.05 ;
      RECT  0.585 0.05 0.755 0.315 ;
      RECT  1.105 0.05 1.275 0.315 ;
      RECT  1.625 0.05 1.795 0.315 ;
      RECT  2.145 0.05 2.315 0.315 ;
      RECT  2.665 0.05 2.835 0.315 ;
      RECT  3.185 0.05 3.355 0.315 ;
      RECT  8.31 0.05 8.48 0.32 ;
      RECT  8.83 0.05 9.0 0.32 ;
      RECT  9.35 0.05 9.52 0.32 ;
      RECT  9.87 0.05 10.04 0.32 ;
      RECT  10.39 0.05 10.56 0.32 ;
      RECT  10.91 0.05 11.08 0.32 ;
      RECT  6.25 0.05 6.38 0.38 ;
      RECT  6.77 0.05 6.9 0.38 ;
      RECT  7.29 0.05 7.42 0.38 ;
      RECT  7.81 0.05 7.94 0.38 ;
      RECT  3.73 0.05 3.84 0.385 ;
      RECT  0.065 0.05 0.185 0.585 ;
      RECT  11.48 0.05 11.6 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 11.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
      RECT  5.85 -0.05 5.95 0.05 ;
      RECT  6.45 -0.05 6.55 0.05 ;
      RECT  7.05 -0.05 7.15 0.05 ;
      RECT  7.65 -0.05 7.75 0.05 ;
      RECT  8.25 -0.05 8.35 0.05 ;
      RECT  8.85 -0.05 8.95 0.05 ;
      RECT  9.45 -0.05 9.55 0.05 ;
      RECT  10.05 -0.05 10.15 0.05 ;
      RECT  10.65 -0.05 10.75 0.05 ;
      RECT  11.25 -0.05 11.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.51 5.88 0.69 ;
      RECT  5.71 0.69 5.88 1.11 ;
      RECT  3.655 1.11 7.935 1.29 ;
      RECT  7.815 1.02 7.935 1.11 ;
    END
    ANTENNADIFFAREA 1.361 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.93 0.205 6.145 0.375 ;
      RECT  5.975 0.375 6.145 0.47 ;
      RECT  3.93 0.375 4.035 0.69 ;
      RECT  5.975 0.47 8.195 0.64 ;
      RECT  7.555 0.32 7.675 0.47 ;
      RECT  8.075 0.27 8.195 0.47 ;
      RECT  8.285 0.42 11.37 0.55 ;
      RECT  8.285 0.55 8.375 0.82 ;
      RECT  6.55 0.82 8.375 0.93 ;
      RECT  8.26 0.93 8.375 1.2 ;
      RECT  8.26 1.2 9.47 1.33 ;
      RECT  3.15 0.78 4.975 0.9 ;
      RECT  3.15 0.9 3.255 1.18 ;
      RECT  0.275 0.405 3.64 0.535 ;
      RECT  1.9 0.535 2.03 1.18 ;
      RECT  1.9 1.18 3.255 1.305 ;
      RECT  9.585 0.995 11.32 1.165 ;
      RECT  9.585 1.165 9.755 1.425 ;
      RECT  8.0 1.425 9.755 1.595 ;
      RECT  0.065 1.18 1.81 1.34 ;
      RECT  0.065 1.34 0.185 1.4 ;
      RECT  1.615 1.34 1.81 1.415 ;
      RECT  1.615 1.415 3.32 1.585 ;
  END
END SEN_OR4_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4B_1
#      Description : "4-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2|B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4B_1
  CLASS CORE ;
  FOREIGN SEN_OR4B_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.6 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.07 0.925 ;
      RECT  0.95 0.925 1.05 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0648 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.7 0.25 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.52 0.7 0.65 1.6 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.7 0.85 1.3 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0564 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.845 1.41 0.975 1.75 ;
      RECT  0.0 1.75 1.6 1.85 ;
      RECT  1.39 1.41 1.52 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.6 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      RECT  0.32 0.05 0.45 0.39 ;
      RECT  0.85 0.05 0.98 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.6 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.31 1.505 0.6 ;
      RECT  1.35 0.6 1.54 0.69 ;
      RECT  1.44 0.69 1.54 1.11 ;
      RECT  1.145 1.11 1.54 1.29 ;
      RECT  1.145 1.29 1.25 1.5 ;
    END
    ANTENNADIFFAREA 0.205 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.32 0.185 0.5 ;
      RECT  0.065 0.5 1.25 0.59 ;
      RECT  0.585 0.32 0.705 0.5 ;
      RECT  1.16 0.59 1.25 0.8 ;
      RECT  0.34 0.59 0.43 1.41 ;
      RECT  1.16 0.8 1.35 0.9 ;
      RECT  0.065 1.41 0.43 1.5 ;
      RECT  0.065 1.5 0.185 1.63 ;
  END
END SEN_OR4B_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4B_2
#      Description : "4-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2|B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4B_2
  CLASS CORE ;
  FOREIGN SEN_OR4B_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 3.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.55 0.7 3.05 0.89 ;
      RECT  2.95 0.89 3.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1296 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.5 0.25 0.71 ;
      RECT  0.15 0.71 0.45 0.89 ;
      RECT  0.15 0.89 0.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.71 1.05 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.71 1.65 0.89 ;
      RECT  1.55 0.89 1.65 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1128 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.395 1.41 1.525 1.75 ;
      RECT  0.0 1.75 3.2 1.85 ;
      RECT  1.92 1.21 2.04 1.75 ;
      RECT  2.46 1.21 2.58 1.75 ;
      RECT  3.0 1.21 3.12 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 3.2 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      RECT  0.085 0.05 0.215 0.39 ;
      RECT  0.625 0.05 0.755 0.39 ;
      RECT  1.155 0.05 1.285 0.39 ;
      RECT  1.68 0.05 1.81 0.39 ;
      RECT  2.735 0.05 2.865 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 3.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.4 0.69 ;
      RECT  2.31 0.69 2.4 0.71 ;
      RECT  2.31 0.71 2.45 1.0 ;
      RECT  2.15 1.0 2.85 1.1 ;
      RECT  2.15 1.1 2.3 1.3 ;
      RECT  2.745 1.1 2.85 1.3 ;
    END
    ANTENNADIFFAREA 0.336 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.96 0.16 2.615 0.25 ;
      RECT  1.96 0.25 2.08 0.39 ;
      RECT  2.495 0.25 2.615 0.5 ;
      RECT  2.495 0.5 3.12 0.59 ;
      RECT  3.0 0.37 3.12 0.5 ;
      RECT  0.37 0.32 0.49 0.5 ;
      RECT  0.37 0.5 2.05 0.59 ;
      RECT  0.89 0.32 1.01 0.5 ;
      RECT  1.42 0.32 1.55 0.5 ;
      RECT  1.95 0.59 2.05 0.785 ;
      RECT  0.555 0.59 0.645 1.01 ;
      RECT  1.95 0.785 2.2 0.89 ;
      RECT  0.37 1.01 0.645 1.1 ;
      RECT  0.37 1.1 0.49 1.24 ;
      RECT  0.865 1.21 1.78 1.31 ;
      RECT  1.66 1.31 1.78 1.43 ;
      RECT  0.07 1.45 1.305 1.55 ;
  END
END SEN_OR4B_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4B_4
#      Description : "4-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2|B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4B_4
  CLASS CORE ;
  FOREIGN SEN_OR4B_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 5.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.95 0.7 5.45 0.89 ;
      RECT  5.35 0.89 5.45 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2592 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.85 0.89 ;
      RECT  0.75 0.89 0.85 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2253 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2253 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.71 3.25 0.89 ;
      RECT  3.15 0.89 3.25 1.1 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2253 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.43 1.41 2.56 1.75 ;
      RECT  0.0 1.75 5.8 1.85 ;
      RECT  2.92 1.41 3.11 1.75 ;
      RECT  3.5 1.21 3.62 1.75 ;
      RECT  4.035 1.41 4.165 1.75 ;
      RECT  4.555 1.41 4.685 1.75 ;
      RECT  5.075 1.41 5.205 1.75 ;
      RECT  5.61 1.21 5.73 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 5.8 1.85 ;
      LAYER V1 ;
      RECT  0.45 1.75 0.55 1.85 ;
      RECT  1.05 1.75 1.15 1.85 ;
      RECT  1.65 1.75 1.75 1.85 ;
      RECT  2.25 1.75 2.35 1.85 ;
      RECT  2.85 1.75 2.95 1.85 ;
      RECT  3.45 1.75 3.55 1.85 ;
      RECT  4.05 1.75 4.15 1.85 ;
      RECT  4.65 1.75 4.75 1.85 ;
      RECT  5.25 1.75 5.35 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      RECT  0.42 0.05 0.55 0.39 ;
      RECT  1.105 0.05 1.235 0.39 ;
      RECT  1.81 0.05 1.935 0.39 ;
      RECT  2.555 0.05 2.685 0.39 ;
      RECT  3.21 0.05 3.34 0.39 ;
      RECT  4.815 0.05 4.945 0.39 ;
      RECT  5.335 0.05 5.465 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 5.8 0.05 ;
      LAYER V1 ;
      RECT  0.45 -0.05 0.55 0.05 ;
      RECT  1.05 -0.05 1.15 0.05 ;
      RECT  1.65 -0.05 1.75 0.05 ;
      RECT  2.25 -0.05 2.35 0.05 ;
      RECT  2.85 -0.05 2.95 0.05 ;
      RECT  3.45 -0.05 3.55 0.05 ;
      RECT  4.05 -0.05 4.15 0.05 ;
      RECT  4.65 -0.05 4.75 0.05 ;
      RECT  5.25 -0.05 5.35 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  3.75 0.51 4.46 0.69 ;
      RECT  4.35 0.69 4.46 1.11 ;
      RECT  3.75 1.11 5.25 1.21 ;
      RECT  3.75 1.21 5.5 1.29 ;
      RECT  5.075 1.29 5.5 1.31 ;
    END
    ANTENNADIFFAREA 0.672 ;
  END X
  OBS
      LAYER M1 ;
      RECT  3.47 0.24 4.68 0.34 ;
      RECT  4.56 0.34 4.68 0.48 ;
      RECT  4.56 0.48 5.73 0.59 ;
      RECT  5.61 0.37 5.73 0.48 ;
      RECT  0.075 0.37 0.195 0.48 ;
      RECT  0.075 0.48 3.6 0.59 ;
      RECT  3.48 0.59 3.6 0.79 ;
      RECT  1.08 0.59 1.22 1.21 ;
      RECT  3.48 0.79 4.24 0.89 ;
      RECT  0.3 1.21 1.22 1.32 ;
      RECT  1.33 1.21 3.39 1.32 ;
      RECT  0.085 1.33 0.2 1.45 ;
      RECT  0.085 1.45 2.34 1.55 ;
  END
END SEN_OR4B_4
#-----------------------------------------------------------------------
#      Cell        : SEN_OR4B_8
#      Description : "4-Input OR (A inverted input)"
#      Equation    : X=!A|B1|B2|B3
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR4B_8
  CLASS CORE ;
  FOREIGN SEN_OR4B_8 0 0 ;
  ORIGIN 0 0 ;
  SIZE 8.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.75 0.71 8.25 0.89 ;
      RECT  8.15 0.89 8.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.5184 ;
  END A
  PIN B1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.61 1.0 0.72 ;
      RECT  0.35 0.72 0.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2943 ;
  END B1
  PIN B2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.55 0.65 2.45 0.89 ;
      RECT  1.55 0.89 1.65 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2943 ;
  END B2
  PIN B3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.75 0.67 3.65 0.89 ;
      RECT  2.75 0.89 2.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2943 ;
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  2.92 1.415 3.05 1.75 ;
      RECT  0.0 1.75 8.4 1.85 ;
      RECT  3.44 1.415 3.57 1.75 ;
      RECT  4.015 1.21 4.135 1.75 ;
      RECT  4.57 1.41 4.7 1.75 ;
      RECT  5.09 1.41 5.22 1.75 ;
      RECT  5.61 1.41 5.74 1.75 ;
      RECT  6.13 1.41 6.26 1.75 ;
      RECT  6.65 1.41 6.78 1.75 ;
      RECT  7.17 1.41 7.3 1.75 ;
      RECT  7.69 1.41 7.82 1.75 ;
      RECT  8.215 1.21 8.335 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 8.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
      RECT  8.05 1.75 8.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      RECT  0.3 0.05 0.47 0.32 ;
      RECT  0.82 0.05 0.99 0.32 ;
      RECT  1.34 0.05 1.51 0.32 ;
      RECT  1.86 0.05 2.03 0.32 ;
      RECT  2.38 0.05 2.55 0.32 ;
      RECT  2.9 0.05 3.07 0.32 ;
      RECT  3.42 0.05 3.59 0.32 ;
      RECT  6.39 0.05 6.52 0.38 ;
      RECT  6.91 0.05 7.04 0.4 ;
      RECT  7.43 0.05 7.56 0.4 ;
      RECT  7.95 0.05 8.08 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 8.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
      RECT  8.05 -0.05 8.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  4.15 0.51 6.035 0.645 ;
      RECT  4.15 0.645 5.91 0.69 ;
      RECT  5.74 0.69 5.91 1.11 ;
      RECT  4.265 1.11 8.06 1.29 ;
    END
    ANTENNADIFFAREA 1.344 ;
  END X
  OBS
      LAYER M1 ;
      RECT  4.005 0.24 6.29 0.37 ;
      RECT  5.59 0.37 6.29 0.395 ;
      RECT  6.135 0.395 6.29 0.47 ;
      RECT  6.135 0.47 6.815 0.51 ;
      RECT  6.135 0.51 8.335 0.62 ;
      RECT  8.215 0.4 8.335 0.51 ;
      RECT  0.065 0.25 0.185 0.41 ;
      RECT  0.065 0.41 3.89 0.5 ;
      RECT  0.585 0.25 0.705 0.41 ;
      RECT  1.105 0.25 1.225 0.41 ;
      RECT  1.625 0.25 1.745 0.41 ;
      RECT  2.145 0.25 2.265 0.41 ;
      RECT  2.665 0.25 2.785 0.41 ;
      RECT  1.1 0.5 3.89 0.54 ;
      RECT  3.76 0.54 3.89 0.785 ;
      RECT  1.1 0.54 1.23 1.255 ;
      RECT  3.76 0.785 5.645 0.915 ;
      RECT  0.06 1.255 1.23 1.385 ;
      RECT  0.06 1.385 0.185 1.475 ;
      RECT  1.575 1.195 3.875 1.325 ;
      RECT  0.275 1.48 2.575 1.61 ;
  END
END SEN_OR4B_8
#-----------------------------------------------------------------------
#      Cell        : SEN_OR5_1
#      Description : "5-Input OR"
#      Equation    : X=A1|A2|A3|A4|A5
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR5_1
  CLASS CORE ;
  FOREIGN SEN_OR5_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 2.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.51 0.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0552 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.35 0.71 0.545 0.81 ;
      RECT  0.35 0.81 0.45 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0552 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.75 0.675 0.85 0.91 ;
      RECT  0.55 0.91 0.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0552 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.51 2.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0483 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.75 0.71 2.05 0.89 ;
      RECT  1.95 0.89 2.05 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0483 ;
  END A5
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.975 1.41 1.105 1.75 ;
      RECT  0.0 1.75 2.4 1.85 ;
      RECT  1.64 1.41 1.77 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 2.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      RECT  0.58 0.05 0.71 0.36 ;
      RECT  0.06 0.05 0.19 0.39 ;
      RECT  2.175 0.05 2.305 0.39 ;
      RECT  1.64 0.05 1.77 0.4 ;
      LAYER M2 ;
      RECT  0.0 -0.05 2.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  1.12 0.51 1.45 0.69 ;
      RECT  1.35 0.69 1.45 1.37 ;
      RECT  1.35 1.37 1.49 1.54 ;
    END
    ANTENNADIFFAREA 0.187 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.845 0.28 0.965 0.445 ;
      RECT  0.845 0.445 1.03 0.45 ;
      RECT  0.34 0.28 0.445 0.45 ;
      RECT  0.34 0.45 1.03 0.54 ;
      RECT  0.94 0.54 1.03 0.81 ;
      RECT  0.94 0.81 1.26 0.92 ;
      RECT  0.94 0.92 1.03 1.22 ;
      RECT  0.795 1.22 1.03 1.31 ;
      RECT  0.795 1.31 0.885 1.46 ;
      RECT  0.065 1.33 0.185 1.46 ;
      RECT  0.065 1.46 0.885 1.55 ;
      RECT  1.92 0.29 2.04 0.5 ;
      RECT  1.55 0.5 2.04 0.59 ;
      RECT  1.55 0.59 1.66 1.18 ;
      RECT  1.55 1.18 2.3 1.3 ;
      RECT  2.18 1.3 2.3 1.4 ;
  END
END SEN_OR5_1
#-----------------------------------------------------------------------
#      Cell        : SEN_OR5_2
#      Description : "5-Input OR"
#      Equation    : X=A1|A2|A3|A4|A5
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR5_2
  CLASS CORE ;
  FOREIGN SEN_OR5_2 0 0 ;
  ORIGIN 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.71 0.25 1.29 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1104 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.15 0.51 1.25 0.71 ;
      RECT  0.75 0.71 1.25 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1104 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  1.35 0.51 1.65 0.69 ;
      RECT  1.35 0.69 1.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1104 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.55 0.71 3.85 0.89 ;
      RECT  3.75 0.89 3.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  3.95 0.71 4.25 0.89 ;
      RECT  4.15 0.89 4.25 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0966 ;
  END A5
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  1.37 1.4 1.5 1.75 ;
      RECT  0.0 1.75 4.4 1.85 ;
      RECT  1.895 1.21 2.015 1.75 ;
      RECT  2.41 1.41 2.54 1.75 ;
      RECT  2.94 1.19 3.055 1.75 ;
      RECT  3.96 1.4 4.09 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 4.4 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      RECT  1.09 0.05 1.26 0.24 ;
      RECT  2.67 0.05 2.8 0.36 ;
      RECT  3.705 0.05 3.825 0.385 ;
      RECT  4.225 0.05 4.345 0.39 ;
      RECT  3.18 0.05 3.31 0.405 ;
      RECT  1.62 0.05 1.79 0.415 ;
      RECT  0.58 0.05 0.71 0.44 ;
      RECT  0.06 0.05 0.19 0.51 ;
      LAYER M2 ;
      RECT  0.0 -0.05 4.4 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  2.15 0.49 2.275 0.67 ;
      RECT  2.15 0.67 2.45 0.76 ;
      RECT  2.35 0.76 2.45 1.11 ;
      RECT  2.15 1.11 2.85 1.29 ;
    END
    ANTENNADIFFAREA 0.316 ;
  END X
  OBS
      LAYER M1 ;
      RECT  1.895 0.215 2.535 0.335 ;
      RECT  1.895 0.335 2.015 0.435 ;
      RECT  2.415 0.335 2.535 0.46 ;
      RECT  2.415 0.46 3.105 0.58 ;
      RECT  3.445 0.27 3.565 0.49 ;
      RECT  3.35 0.49 4.085 0.58 ;
      RECT  3.965 0.27 4.085 0.49 ;
      RECT  3.35 0.58 3.44 0.81 ;
      RECT  2.655 0.81 3.44 0.92 ;
      RECT  3.35 0.92 3.44 1.1 ;
      RECT  3.35 1.1 3.615 1.22 ;
      RECT  1.54 0.85 2.23 0.96 ;
      RECT  1.54 0.96 1.63 0.98 ;
      RECT  0.845 0.33 1.53 0.42 ;
      RECT  0.845 0.42 0.965 0.53 ;
      RECT  0.34 0.37 0.445 0.53 ;
      RECT  0.34 0.53 0.965 0.62 ;
      RECT  0.34 0.62 0.445 0.98 ;
      RECT  0.34 0.98 1.63 1.07 ;
      RECT  0.34 1.07 0.445 1.23 ;
      RECT  0.795 1.18 1.805 1.3 ;
      RECT  3.705 1.22 4.345 1.31 ;
      RECT  3.705 1.31 3.825 1.44 ;
      RECT  4.225 1.31 4.345 1.61 ;
      RECT  3.185 1.34 3.305 1.44 ;
      RECT  3.185 1.44 3.825 1.56 ;
      RECT  0.065 1.39 0.185 1.48 ;
      RECT  0.065 1.48 1.245 1.61 ;
      RECT  1.125 1.39 1.245 1.48 ;
  END
END SEN_OR5_2
#-----------------------------------------------------------------------
#      Cell        : SEN_OR5_4
#      Description : "5-Input OR"
#      Equation    : X=A1|A2|A3|A4|A5
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_OR5_4
  CLASS CORE ;
  FOREIGN SEN_OR5_4 0 0 ;
  ORIGIN 0 0 ;
  SIZE 7.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN A1
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  6.95 0.71 7.45 0.89 ;
      RECT  7.35 0.89 7.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2214 ;
  END A1
  PIN A2
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  5.95 0.71 6.45 0.89 ;
      RECT  6.35 0.89 6.45 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2214 ;
  END A2
  PIN A3
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.75 0.71 5.25 0.89 ;
      RECT  4.75 0.89 4.85 1.09 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2214 ;
  END A3
  PIN A4
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  2.95 0.51 3.05 0.71 ;
      RECT  2.95 0.71 3.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1929 ;
  END A4
  PIN A5
    DIRECTION INPUT ;
    PORT
      LAYER M1 ;
      RECT  4.35 0.51 4.45 0.71 ;
      RECT  3.75 0.71 4.45 0.89 ;
    END
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1929 ;
  END A5
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.065 1.21 0.185 1.75 ;
      RECT  0.0 1.75 7.8 1.85 ;
      RECT  0.58 1.41 0.71 1.75 ;
      RECT  1.1 1.41 1.23 1.75 ;
      RECT  1.62 1.41 1.75 1.75 ;
      RECT  2.145 1.18 2.265 1.75 ;
      RECT  3.76 1.415 3.87 1.75 ;
      RECT  4.265 1.21 4.385 1.75 ;
      RECT  4.78 1.44 4.91 1.75 ;
      RECT  5.3 1.43 5.43 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 7.8 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
      RECT  1.45 1.75 1.55 1.85 ;
      RECT  2.05 1.75 2.15 1.85 ;
      RECT  2.65 1.75 2.75 1.85 ;
      RECT  3.25 1.75 3.35 1.85 ;
      RECT  3.85 1.75 3.95 1.85 ;
      RECT  4.45 1.75 4.55 1.85 ;
      RECT  5.05 1.75 5.15 1.85 ;
      RECT  5.65 1.75 5.75 1.85 ;
      RECT  6.25 1.75 6.35 1.85 ;
      RECT  6.85 1.75 6.95 1.85 ;
      RECT  7.45 1.75 7.55 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      RECT  2.65 0.05 2.82 0.2 ;
      RECT  3.19 0.05 3.36 0.2 ;
      RECT  3.72 0.05 3.89 0.32 ;
      RECT  4.76 0.05 4.93 0.32 ;
      RECT  5.325 0.05 5.455 0.36 ;
      RECT  5.715 0.05 5.845 0.36 ;
      RECT  6.255 0.05 6.385 0.36 ;
      RECT  6.8 0.05 6.93 0.36 ;
      RECT  4.26 0.05 4.39 0.39 ;
      RECT  1.36 0.05 1.49 0.4 ;
      RECT  1.88 0.05 2.01 0.4 ;
      RECT  7.37 0.05 7.49 0.59 ;
      LAYER M2 ;
      RECT  0.0 -0.05 7.8 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
      RECT  1.45 -0.05 1.55 0.05 ;
      RECT  2.05 -0.05 2.15 0.05 ;
      RECT  2.65 -0.05 2.75 0.05 ;
      RECT  3.25 -0.05 3.35 0.05 ;
      RECT  3.85 -0.05 3.95 0.05 ;
      RECT  4.45 -0.05 4.55 0.05 ;
      RECT  5.05 -0.05 5.15 0.05 ;
      RECT  5.65 -0.05 5.75 0.05 ;
      RECT  6.25 -0.05 6.35 0.05 ;
      RECT  6.85 -0.05 6.95 0.05 ;
      RECT  7.45 -0.05 7.55 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.34 0.51 1.05 0.69 ;
      RECT  0.34 0.69 0.45 1.11 ;
      RECT  0.34 1.11 2.05 1.29 ;
    END
    ANTENNADIFFAREA 0.632 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.065 0.2 1.25 0.32 ;
      RECT  0.065 0.32 0.185 0.42 ;
      RECT  1.14 0.32 1.25 0.49 ;
      RECT  1.14 0.49 2.265 0.61 ;
      RECT  2.145 0.39 2.265 0.49 ;
      RECT  2.405 0.29 3.63 0.41 ;
      RECT  3.54 0.41 4.17 0.52 ;
      RECT  2.405 0.41 2.525 0.74 ;
      RECT  1.47 0.74 2.73 0.84 ;
      RECT  2.64 0.84 2.73 1.1 ;
      RECT  2.64 1.1 3.31 1.205 ;
      RECT  3.195 1.01 3.31 1.1 ;
      RECT  4.54 0.29 4.645 0.41 ;
      RECT  4.54 0.41 5.19 0.45 ;
      RECT  4.54 0.45 7.235 0.565 ;
      RECT  6.75 0.565 7.235 0.57 ;
      RECT  4.54 0.565 4.63 0.98 ;
      RECT  6.75 0.57 6.86 1.24 ;
      RECT  3.4 0.98 4.63 1.085 ;
      RECT  3.4 1.085 3.49 1.295 ;
      RECT  6.75 1.24 7.48 1.36 ;
      RECT  0.56 0.805 1.245 0.915 ;
      RECT  1.155 0.915 1.245 0.93 ;
      RECT  1.155 0.93 2.51 1.02 ;
      RECT  2.42 1.02 2.51 1.295 ;
      RECT  2.42 1.295 3.49 1.385 ;
      RECT  5.44 1.005 6.13 1.125 ;
      RECT  6.01 1.125 6.13 1.205 ;
      RECT  6.01 1.205 6.65 1.325 ;
      RECT  6.53 1.325 6.65 1.46 ;
      RECT  6.53 1.46 7.74 1.58 ;
      RECT  3.58 1.205 4.175 1.325 ;
      RECT  3.58 1.325 3.67 1.48 ;
      RECT  2.355 1.48 3.67 1.6 ;
      RECT  4.475 1.22 5.615 1.34 ;
      RECT  5.525 1.34 5.615 1.415 ;
      RECT  5.525 1.415 6.44 1.535 ;
  END
END SEN_OR5_4
#-----------------------------------------------------------------------
#      Cell        : SEN_TIE0_1
#      Description : "Tie low"
#      Equation    : X=0
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_TIE0_1
  CLASS CORE TIELOW ;
  FOREIGN SEN_TIE0_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.435 1.41 0.565 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.985 1.405 1.115 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.985 0.05 1.115 0.39 ;
      RECT  0.425 0.05 0.545 0.605 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.31 0.25 1.09 ;
    END
    ANTENNADIFFAREA 0.084 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.72 0.23 0.84 0.525 ;
      RECT  0.72 0.525 1.08 0.635 ;
      RECT  0.38 1.165 0.84 1.275 ;
      RECT  0.72 1.275 0.84 1.58 ;
  END
END SEN_TIE0_1
#-----------------------------------------------------------------------
#      Cell        : SEN_TIE1_1
#      Description : "Tie high"
#      Equation    : X=1
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_TIE1_1
  CLASS CORE TIEHIGH ;
  FOREIGN SEN_TIE1_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 1.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.085 1.41 0.215 1.75 ;
      RECT  0.0 1.75 1.2 1.85 ;
      RECT  0.64 1.21 0.76 1.75 ;
      LAYER M2 ;
      RECT  0.0 1.75 1.2 1.85 ;
      LAYER V1 ;
      RECT  0.25 1.75 0.35 1.85 ;
      RECT  0.85 1.75 0.95 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      RECT  0.085 0.05 0.215 0.39 ;
      RECT  0.645 0.05 0.775 0.39 ;
      LAYER M2 ;
      RECT  0.0 -0.05 1.2 0.05 ;
      LAYER V1 ;
      RECT  0.25 -0.05 0.35 0.05 ;
      RECT  0.85 -0.05 0.95 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION OUTPUT ;
    PORT
      LAYER M1 ;
      RECT  0.95 0.71 1.05 1.49 ;
    END
    ANTENNADIFFAREA 0.123 ;
  END X
  OBS
      LAYER M1 ;
      RECT  0.36 0.22 0.48 0.525 ;
      RECT  0.36 0.525 0.8 0.635 ;
      RECT  0.125 1.165 0.475 1.275 ;
      RECT  0.365 1.275 0.475 1.59 ;
  END
END SEN_TIE1_1
#-----------------------------------------------------------------------
#      Cell        : SEN_TIEDIN_1
#      Description : "Antenna diode with N+/Pwell Diode"
#      Equation    : X=tristate(enable=0,data=0)
#      Version     : 5.6
#      Created     : 2007/10/29 19:10:27
#
MACRO SEN_TIEDIN_1
  CLASS CORE ANTENNACELL ;
  FOREIGN SEN_TIEDIN_1 0 0 ;
  ORIGIN 0 0 ;
  SIZE 0.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE cp65_dst ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 1.75 0.4 1.85 ;
      LAYER M2 ;
      RECT  0.0 1.75 0.4 1.85 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
      RECT  0.0 -0.05 0.4 0.05 ;
      LAYER M2 ;
      RECT  0.0 -0.05 0.4 0.05 ;
    END
  END VSS
  PIN X
    DIRECTION INOUT ;
    PORT
      LAYER M1 ;
      RECT  0.15 0.265 0.25 1.09 ;
    END
    ANTENNADIFFAREA 0.144 ;
  END X
END SEN_TIEDIN_1

END LIBRARY
