
module ShiftLR ( Z, X, S, LEFT, LOG );
  output [31:0] Z;
  input [31:0] X;
  input [4:0] S;
  input LEFT, LOG;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222;

  SEN_AN2_4 U224 ( .A1(n81), .A2(n40), .X(n220) );
  SEN_OAI21_G_1 U225 ( .A1(n40), .A2(n34), .B(n148), .X(n87) );
  SEN_EO2_G_2 U226 ( .A1(n188), .A2(S[3]), .X(n108) );
  SEN_ND2_G_1 U227 ( .A1(LEFT), .A2(n187), .X(n188) );
  SEN_EO2_DG_2 U228 ( .A1(S[2]), .A2(n190), .X(n66) );
  SEN_ND2_0P8 U229 ( .A1(n108), .A2(n66), .X(n111) );
  SEN_INV_2 U230 ( .A(n66), .X(n46) );
  SEN_INV_S_2 U231 ( .A(n111), .X(n45) );
  SEN_OAI221_1 U232 ( .A1(n20), .A2(n111), .B1(n120), .B2(n97), .C(n109), .X(
        n104) );
  SEN_OAI221_1 U233 ( .A1(n23), .A2(n111), .B1(n112), .B2(n97), .C(n109), .X(
        n100) );
  SEN_BUF_1 U234 ( .A(n66), .X(n197) );
  SEN_AOI22_0P75 U235 ( .A1(n51), .A2(n104), .B1(n48), .B2(n100), .X(n110) );
  SEN_AOI22_0P5 U236 ( .A1(n51), .A2(n100), .B1(n48), .B2(n93), .X(n102) );
  SEN_AOI22_0P75 U237 ( .A1(n47), .A2(n93), .B1(n50), .B2(n100), .X(n99) );
  SEN_INV_5 U238 ( .A(n108), .X(n44) );
  SEN_OA22_DG_2 U239 ( .A1(n3), .A2(n66), .B1(n73), .B2(n46), .X(n63) );
  SEN_ND2_0P8 U240 ( .A1(n81), .A2(n44), .X(n109) );
  SEN_ND2_S_0P5 U241 ( .A1(n43), .A2(n81), .X(n124) );
  SEN_OA21B_1 U242 ( .A1(n94), .A2(n66), .B(n81), .X(n80) );
  SEN_AOI22_0P5 U243 ( .A1(n51), .A2(n82), .B1(n48), .B2(n81), .X(n89) );
  SEN_ND2_G_4 U244 ( .A1(n209), .A2(n210), .X(n160) );
  SEN_ND2_G_1 U245 ( .A1(n211), .A2(S[4]), .X(n210) );
  SEN_ND2_S_2 U246 ( .A1(n186), .A2(n208), .X(n209) );
  SEN_ND2_3 U247 ( .A1(n46), .A2(n108), .X(n97) );
  SEN_AO21B_1 U248 ( .A1(n160), .A2(X[23]), .B(n148), .X(n126) );
  SEN_ND3_S_0P5 U249 ( .A1(n221), .A2(n222), .A3(n155), .X(n146) );
  SEN_OR3_1 U250 ( .A1(n204), .A2(n205), .A3(n193), .X(n143) );
  SEN_ND2B_V1_4 U251 ( .A(S[2]), .B(n189), .X(n187) );
  SEN_OAI21_S_1 U252 ( .A1(S[3]), .A2(n187), .B(LEFT), .X(n186) );
  SEN_NR2_T_6 U253 ( .A1(S[1]), .A2(S[0]), .X(n189) );
  SEN_INV_2 U254 ( .A(n192), .X(n216) );
  SEN_AO21B_1 U255 ( .A1(n160), .A2(X[21]), .B(n148), .X(n137) );
  SEN_OA22_1 U256 ( .A1(n68), .A2(n57), .B1(n75), .B2(n49), .X(n71) );
  SEN_INV_S_1 U257 ( .A(n150), .X(n2) );
  SEN_ND3_S_0P5 U258 ( .A1(n214), .A2(n215), .A3(n144), .X(n135) );
  SEN_INV_S_1 U259 ( .A(n135), .X(n8) );
  SEN_INV_S_1 U260 ( .A(n123), .X(n6) );
  SEN_NR3_1 U261 ( .A1(LOG), .A2(LEFT), .A3(n25), .X(n81) );
  SEN_NR2_1 U262 ( .A1(n206), .A2(n207), .X(n149) );
  SEN_OA2BB2_1 U263 ( .A1(n158), .A2(n49), .B1(n60), .B2(n49), .X(n53) );
  SEN_OR2_DG_1 U264 ( .A1(n44), .A2(n160), .X(n192) );
  SEN_INV_5 U265 ( .A(n220), .X(n148) );
  SEN_OR2_1 U266 ( .A1(n212), .A2(n213), .X(n193) );
  SEN_OR2_1 U267 ( .A1(n218), .A2(n217), .X(n194) );
  SEN_ND2_2 U268 ( .A1(n46), .A2(n44), .X(n106) );
  SEN_INV_S_1 U269 ( .A(n50), .X(n195) );
  SEN_INV_S_0P5 U270 ( .A(n47), .X(n196) );
  SEN_INV_1 U271 ( .A(n79), .X(n47) );
  SEN_OA21_2 U272 ( .A1(S[3]), .A2(n187), .B(LEFT), .X(n211) );
  SEN_OAI222_0P75 U273 ( .A1(n19), .A2(n111), .B1(n112), .B2(n156), .C1(n163), 
        .C2(n197), .X(n154) );
  SEN_AOI222_0P5 U274 ( .A1(n216), .A2(X[26]), .B1(n86), .B2(X[10]), .C1(n164), 
        .C2(n44), .X(n76) );
  SEN_AOI222_0P5 U275 ( .A1(n216), .A2(X[28]), .B1(n86), .B2(X[12]), .C1(n141), 
        .C2(n44), .X(n69) );
  SEN_AOI222_0P5 U276 ( .A1(n216), .A2(X[30]), .B1(n86), .B2(X[14]), .C1(n133), 
        .C2(n44), .X(n163) );
  SEN_NR2_G_0P5 U277 ( .A1(n97), .A2(n40), .X(n171) );
  SEN_OAI221_0P5 U278 ( .A1(n36), .A2(n173), .B1(n25), .B2(n174), .C(n185), 
        .X(n184) );
  SEN_OAI21_0P5 U279 ( .A1(n40), .A2(n25), .B(n24), .X(n107) );
  SEN_NR2_G_1 U280 ( .A1(n219), .A2(n194), .X(n73) );
  SEN_AN2_S_1 U281 ( .A1(n161), .A2(n44), .X(n219) );
  SEN_NR2B_V1_1 U282 ( .A(LEFT), .B(n189), .X(n190) );
  SEN_OR2_1 U283 ( .A1(n13), .A2(n111), .X(n198) );
  SEN_OR2_1 U284 ( .A1(n120), .A2(n156), .X(n199) );
  SEN_OR2_DG_1 U285 ( .A1(n69), .A2(n66), .X(n200) );
  SEN_ND3_1 U286 ( .A1(n198), .A2(n199), .A3(n200), .X(n158) );
  SEN_AN2_S_0P5 U287 ( .A1(n216), .A2(X[25]), .X(n201) );
  SEN_AN2_DG_1 U288 ( .A1(n86), .A2(X[9]), .X(n202) );
  SEN_AN2_S_0P5 U289 ( .A1(n87), .A2(n44), .X(n203) );
  SEN_NR3_G_1 U290 ( .A1(n201), .A2(n202), .A3(n203), .X(n65) );
  SEN_OA22_DG_1 U291 ( .A1(n28), .A2(n66), .B1(n65), .B2(n46), .X(n72) );
  SEN_NR2_1 U292 ( .A1(n117), .A2(n106), .X(n204) );
  SEN_NR2_S_0P5 U293 ( .A1(n5), .A2(n97), .X(n205) );
  SEN_AOI22_1 U294 ( .A1(n51), .A2(n143), .B1(n48), .B2(n135), .X(n142) );
  SEN_OAI211_1 U295 ( .A1(n120), .A2(n111), .B1(n124), .B2(n140), .X(n131) );
  SEN_OAI221_0P5 U296 ( .A1(n152), .A2(n90), .B1(n2), .B2(n91), .C(n157), .X(
        Z[12]) );
  SEN_OAI221_0P5 U297 ( .A1(n4), .A2(n79), .B1(n2), .B2(n78), .C(n145), .X(
        Z[15]) );
  SEN_OAI221_0P5 U298 ( .A1(n2), .A2(n196), .B1(n152), .B2(n78), .C(n153), .X(
        Z[13]) );
  SEN_AN2_1 U299 ( .A1(n51), .A2(n150), .X(n206) );
  SEN_AN2_DG_1 U300 ( .A1(n48), .A2(n143), .X(n207) );
  SEN_INV_1 U301 ( .A(n90), .X(n51) );
  SEN_OAI222_1 U302 ( .A1(n10), .A2(n111), .B1(n105), .B2(n156), .C1(n159), 
        .C2(n197), .X(n150) );
  SEN_INV_1 U303 ( .A(n91), .X(n48) );
  SEN_INV_S_1 U304 ( .A(S[4]), .X(n208) );
  SEN_AOI21B_0P5 U305 ( .A1(n160), .A2(X[27]), .B(n148), .X(n105) );
  SEN_ND2_S_0P8 U306 ( .A1(n160), .A2(n44), .X(n173) );
  SEN_INV_10 U307 ( .A(n160), .X(n40) );
  SEN_AN2_1 U308 ( .A1(n43), .A2(n101), .X(n212) );
  SEN_AN2_S_0P5 U309 ( .A1(n45), .A2(n137), .X(n213) );
  SEN_INV_S_1 U310 ( .A(n143), .X(n4) );
  SEN_INV_2 U311 ( .A(n156), .X(n43) );
  SEN_OAI221_1 U312 ( .A1(n21), .A2(n111), .B1(n117), .B2(n97), .C(n109), .X(
        n114) );
  SEN_OR2_DG_1 U313 ( .A1(n105), .A2(n106), .X(n214) );
  SEN_OR2_DG_1 U314 ( .A1(n10), .A2(n97), .X(n215) );
  SEN_INV_0P5 U315 ( .A(n161), .X(n10) );
  SEN_NR2_T_1 U316 ( .A1(n40), .A2(n44), .X(n86) );
  SEN_OAI211_1 U317 ( .A1(n117), .A2(n111), .B1(n124), .B2(n136), .X(n123) );
  SEN_INV_S_0P5 U318 ( .A(n97), .X(n41) );
  SEN_INV_0P5 U319 ( .A(n114), .X(n7) );
  SEN_INV_1 U320 ( .A(n82), .X(n22) );
  SEN_AOI22_T_0P5 U321 ( .A1(n47), .A2(n82), .B1(n50), .B2(n93), .X(n92) );
  SEN_OAI22_S_1 U322 ( .A1(n53), .A2(n52), .B1(S[0]), .B2(n54), .X(Z[9]) );
  SEN_OAI21_S_0P5 U323 ( .A1(n23), .A2(n97), .B(n98), .X(n82) );
  SEN_OAI21_S_0P5 U324 ( .A1(n20), .A2(n97), .B(n98), .X(n93) );
  SEN_OAI221_1 U325 ( .A1(n112), .A2(n106), .B1(n19), .B2(n97), .C(n147), .X(
        n139) );
  SEN_OAI221_1 U326 ( .A1(n34), .A2(n167), .B1(n28), .B2(n46), .C(n180), .X(
        n179) );
  SEN_AOI22_1 U327 ( .A1(n49), .A2(n84), .B1(n57), .B2(n179), .X(n127) );
  SEN_AN2_S_0P5 U328 ( .A1(n216), .A2(X[27]), .X(n217) );
  SEN_AN2_S_0P5 U329 ( .A1(n86), .A2(X[11]), .X(n218) );
  SEN_OA22_DG_1 U330 ( .A1(n159), .A2(n46), .B1(n73), .B2(n66), .X(n56) );
  SEN_AOI222_0P5 U331 ( .A1(n216), .A2(X[24]), .B1(n86), .B2(X[8]), .C1(n129), 
        .C2(n44), .X(n70) );
  SEN_AOI222_1 U332 ( .A1(n169), .A2(X[25]), .B1(n170), .B2(X[9]), .C1(X[1]), 
        .C2(n171), .X(n180) );
  SEN_OA222_1 U333 ( .A1(n5), .A2(n111), .B1(n117), .B2(n156), .C1(n64), .C2(
        n66), .X(n152) );
  SEN_AOI22_0P5 U334 ( .A1(n47), .A2(n100), .B1(n50), .B2(n104), .X(n103) );
  SEN_ND2_T_0P5 U335 ( .A1(n41), .A2(n40), .X(n167) );
  SEN_AOI22_0P5 U336 ( .A1(n51), .A2(n119), .B1(n48), .B2(n104), .X(n118) );
  SEN_AOI22_0P5 U337 ( .A1(n51), .A2(n116), .B1(n48), .B2(n114), .X(n115) );
  SEN_INV_S_1 U338 ( .A(n154), .X(n16) );
  SEN_INV_1 U339 ( .A(n121), .X(n20) );
  SEN_INV_S_0P5 U340 ( .A(n146), .X(n12) );
  SEN_AOI22_S_1 U341 ( .A1(n47), .A2(n154), .B1(n50), .B2(n158), .X(n157) );
  SEN_AOI22_0P5 U342 ( .A1(n43), .A2(n121), .B1(n45), .B2(n141), .X(n155) );
  SEN_AOI222_0P5 U343 ( .A1(n216), .A2(X[31]), .B1(n86), .B2(X[15]), .C1(n126), 
        .C2(n44), .X(n159) );
  SEN_AOI222_0P5 U344 ( .A1(n216), .A2(X[29]), .B1(n86), .B2(X[13]), .C1(n137), 
        .C2(n44), .X(n64) );
  SEN_INV_1 U345 ( .A(n181), .X(n28) );
  SEN_OAI21_G_0P5 U346 ( .A1(n127), .A2(n52), .B(n165), .X(Z[0]) );
  SEN_OAI22_S_1 U347 ( .A1(n54), .A2(n52), .B1(S[0]), .B2(n55), .X(Z[8]) );
  SEN_OAI22_S_1 U348 ( .A1(n62), .A2(n52), .B1(S[0]), .B2(n67), .X(Z[5]) );
  SEN_OAI22_S_1 U349 ( .A1(n59), .A2(n52), .B1(S[0]), .B2(n62), .X(Z[6]) );
  SEN_OAI22_S_1 U350 ( .A1(n55), .A2(n52), .B1(S[0]), .B2(n59), .X(Z[7]) );
  SEN_OAI22_S_1 U351 ( .A1(n67), .A2(n52), .B1(S[0]), .B2(n71), .X(Z[4]) );
  SEN_AOI21B_0P5 U352 ( .A1(n160), .A2(X[24]), .B(n148), .X(n120) );
  SEN_OR2_DG_1 U353 ( .A1(n120), .A2(n106), .X(n221) );
  SEN_OR2_DG_1 U354 ( .A1(n13), .A2(n97), .X(n222) );
  SEN_AOI22_S_1 U355 ( .A1(n51), .A2(n146), .B1(n48), .B2(n139), .X(n145) );
  SEN_AOI22_0P75 U356 ( .A1(n51), .A2(n123), .B1(n48), .B2(n116), .X(n122) );
  SEN_AOI22_0P75 U357 ( .A1(n51), .A2(n131), .B1(n48), .B2(n119), .X(n130) );
  SEN_INV_S_0P5 U358 ( .A(n104), .X(n15) );
  SEN_INV_S_0P5 U359 ( .A(n131), .X(n14) );
  SEN_INV_1 U360 ( .A(n113), .X(n23) );
  SEN_INV_S_0P5 U361 ( .A(n116), .X(n9) );
  SEN_INV_S_0P5 U362 ( .A(n119), .X(n18) );
  SEN_INV_S_0P5 U363 ( .A(n87), .X(n5) );
  SEN_AOI22_0P5 U364 ( .A1(n43), .A2(n107), .B1(n45), .B2(n126), .X(n144) );
  SEN_OAI22_T_0P5 U365 ( .A1(n162), .A2(n52), .B1(S[0]), .B2(n53), .X(Z[10])
         );
  SEN_OAI22_T_0P5 U366 ( .A1(n83), .A2(n52), .B1(S[0]), .B2(n127), .X(Z[1]) );
  SEN_OAI22_T_0P5 U367 ( .A1(n74), .A2(n52), .B1(S[0]), .B2(n83), .X(Z[2]) );
  SEN_OAI22_T_0P5 U368 ( .A1(n71), .A2(n52), .B1(S[0]), .B2(n74), .X(Z[3]) );
  SEN_INV_4 U369 ( .A(X[31]), .X(n25) );
  SEN_AOI22_S_1 U370 ( .A1(n51), .A2(n154), .B1(n48), .B2(n146), .X(n153) );
  SEN_AOI22_S_1 U371 ( .A1(n51), .A2(n135), .B1(n48), .B2(n123), .X(n134) );
  SEN_AOI22_S_1 U372 ( .A1(n51), .A2(n139), .B1(n48), .B2(n131), .X(n138) );
  SEN_INV_S_0P5 U373 ( .A(n164), .X(n19) );
  SEN_INV_S_0P5 U374 ( .A(n129), .X(n13) );
  SEN_INV_S_1 U375 ( .A(n139), .X(n17) );
  SEN_ND2_G_1 U376 ( .A1(n49), .A2(n52), .X(n79) );
  SEN_NR2_S_0P5 U377 ( .A1(n106), .A2(n160), .X(n169) );
  SEN_OAI21_S_0P5 U378 ( .A1(n40), .A2(n31), .B(n148), .X(n121) );
  SEN_AOI22_0P5 U379 ( .A1(n43), .A2(n113), .B1(n45), .B2(n133), .X(n147) );
  SEN_OAI21_S_0P5 U380 ( .A1(n40), .A2(n27), .B(n148), .X(n113) );
  SEN_AOI22_0P5 U381 ( .A1(n42), .A2(n121), .B1(n41), .B2(n141), .X(n140) );
  SEN_AOI22_0P5 U382 ( .A1(n42), .A2(n101), .B1(n41), .B2(n137), .X(n136) );
  SEN_OAI211_1 U383 ( .A1(n112), .A2(n111), .B1(n124), .B2(n132), .X(n119) );
  SEN_AOI22_0P5 U384 ( .A1(n42), .A2(n113), .B1(n41), .B2(n133), .X(n132) );
  SEN_OAI211_1 U385 ( .A1(n105), .A2(n111), .B1(n124), .B2(n125), .X(n116) );
  SEN_AOI22_0P5 U386 ( .A1(n42), .A2(n107), .B1(n41), .B2(n126), .X(n125) );
  SEN_ND2_S_0P5 U387 ( .A1(n81), .A2(n97), .X(n98) );
  SEN_OAI21_S_0P5 U388 ( .A1(n40), .A2(n29), .B(n148), .X(n101) );
  SEN_AOI21B_0P5 U389 ( .A1(n107), .A2(n108), .B(n109), .X(n94) );
  SEN_OA22_1 U390 ( .A1(n152), .A2(n57), .B1(n56), .B2(n49), .X(n162) );
  SEN_OA22_DG_1 U391 ( .A1(n26), .A2(n66), .B1(n76), .B2(n46), .X(n68) );
  SEN_OA22_DG_1 U392 ( .A1(n30), .A2(n66), .B1(n70), .B2(n46), .X(n75) );
  SEN_OA22_DG_1 U393 ( .A1(n61), .A2(n57), .B1(n68), .B2(n49), .X(n62) );
  SEN_OA22_DG_1 U394 ( .A1(n58), .A2(n57), .B1(n63), .B2(n49), .X(n59) );
  SEN_OA22_DG_1 U395 ( .A1(n63), .A2(n57), .B1(n72), .B2(n49), .X(n67) );
  SEN_OA22_DG_1 U396 ( .A1(n64), .A2(n46), .B1(n65), .B2(n66), .X(n58) );
  SEN_OA22_DG_1 U397 ( .A1(n163), .A2(n46), .B1(n76), .B2(n66), .X(n60) );
  SEN_AOI21B_0P5 U398 ( .A1(n160), .A2(X[26]), .B(n148), .X(n112) );
  SEN_AOI21B_0P5 U399 ( .A1(n160), .A2(X[25]), .B(n148), .X(n117) );
  SEN_INV_S_0P5 U400 ( .A(n158), .X(n11) );
  SEN_EO2_1 U401 ( .A1(n191), .A2(S[1]), .X(n57) );
  SEN_INV_S_1 U402 ( .A(S[0]), .X(n52) );
  SEN_AO21B_1 U403 ( .A1(n160), .A2(X[20]), .B(n148), .X(n141) );
  SEN_INV_1 U404 ( .A(n172), .X(n26) );
  SEN_AOI22_0P5 U405 ( .A1(X[6]), .A2(n86), .B1(X[22]), .B2(n216), .X(n175) );
  SEN_INV_1 U406 ( .A(n184), .X(n3) );
  SEN_AOI22_0P5 U407 ( .A1(X[7]), .A2(n86), .B1(X[23]), .B2(n216), .X(n185) );
  SEN_INV_1 U408 ( .A(n177), .X(n30) );
  SEN_AOI22_0P5 U409 ( .A1(X[4]), .A2(n86), .B1(X[20]), .B2(n216), .X(n178) );
  SEN_AOI22_0P5 U410 ( .A1(X[5]), .A2(n86), .B1(X[21]), .B2(n216), .X(n182) );
  SEN_AOI22_0P5 U411 ( .A1(n50), .A2(n166), .B1(n47), .B2(n128), .X(n165) );
  SEN_OAI221_0P5 U412 ( .A1(n35), .A2(n167), .B1(n30), .B2(n46), .C(n176), .X(
        n166) );
  SEN_INV_S_1 U413 ( .A(n106), .X(n42) );
  SEN_NR2_1 U414 ( .A1(n106), .A2(n40), .X(n170) );
  SEN_AOI21B_1 U415 ( .A1(n101), .A2(n41), .B(n98), .X(n88) );
  SEN_INV_S_1 U416 ( .A(n78), .X(n50) );
  SEN_OAI221_1 U417 ( .A1(n88), .A2(n79), .B1(n95), .B2(n78), .C(n96), .X(
        Z[27]) );
  SEN_AOI22_1 U418 ( .A1(n51), .A2(n93), .B1(n48), .B2(n82), .X(n96) );
  SEN_OAI221_1 U419 ( .A1(n95), .A2(n79), .B1(n7), .B2(n78), .C(n102), .X(
        Z[25]) );
  SEN_ND2_G_1 U420 ( .A1(n44), .A2(n40), .X(n174) );
  SEN_OAI221_1 U421 ( .A1(n7), .A2(n79), .B1(n9), .B2(n78), .C(n110), .X(Z[23]) );
  SEN_OAI221_1 U422 ( .A1(n12), .A2(n79), .B1(n16), .B2(n78), .C(n149), .X(
        Z[14]) );
  SEN_OAI221_1 U423 ( .A1(n17), .A2(n79), .B1(n12), .B2(n78), .C(n142), .X(
        Z[16]) );
  SEN_OAI221_1 U424 ( .A1(n8), .A2(n79), .B1(n4), .B2(n78), .C(n138), .X(Z[17]) );
  SEN_OAI221_1 U425 ( .A1(n15), .A2(n79), .B1(n18), .B2(n78), .C(n115), .X(
        Z[22]) );
  SEN_OAI221_1 U426 ( .A1(n14), .A2(n79), .B1(n17), .B2(n78), .C(n134), .X(
        Z[18]) );
  SEN_OAI221_1 U427 ( .A1(n6), .A2(n79), .B1(n8), .B2(n78), .C(n130), .X(Z[19]) );
  SEN_OAI221_1 U428 ( .A1(n18), .A2(n79), .B1(n14), .B2(n78), .C(n122), .X(
        Z[20]) );
  SEN_OAI221_1 U429 ( .A1(n9), .A2(n79), .B1(n6), .B2(n78), .C(n118), .X(Z[21]) );
  SEN_INV_1 U430 ( .A(n101), .X(n21) );
  SEN_ND2_G_1 U431 ( .A1(n57), .A2(n52), .X(n78) );
  SEN_OAI222_1 U432 ( .A1(n22), .A2(n195), .B1(n24), .B2(n79), .C1(n77), .C2(
        n52), .X(Z[30]) );
  SEN_OA2BB2_1 U433 ( .A1(n128), .A2(n57), .B1(n75), .B2(n57), .X(n83) );
  SEN_OA2BB2_1 U434 ( .A1(n84), .A2(n57), .B1(n72), .B2(n57), .X(n74) );
  SEN_INV_S_1 U435 ( .A(n81), .X(n24) );
  SEN_OAI221_1 U436 ( .A1(n7), .A2(n90), .B1(n95), .B2(n91), .C(n103), .X(
        Z[24]) );
  SEN_OAI221_1 U437 ( .A1(n95), .A2(n90), .B1(n88), .B2(n91), .C(n99), .X(
        Z[26]) );
  SEN_OAI221_1 U438 ( .A1(n88), .A2(n90), .B1(n80), .B2(n91), .C(n92), .X(
        Z[28]) );
  SEN_ND2_S_0P5 U439 ( .A1(n44), .A2(n66), .X(n156) );
  SEN_OA21B_1 U440 ( .A1(n80), .A2(n49), .B(n81), .X(n77) );
  SEN_OA222_0P5 U441 ( .A1(n105), .A2(n97), .B1(n24), .B2(n106), .C1(n94), 
        .C2(n46), .X(n95) );
  SEN_INV_S_1 U442 ( .A(n57), .X(n49) );
  SEN_OAI21_G_1 U443 ( .A1(n40), .A2(n35), .B(n148), .X(n129) );
  SEN_OAI21_G_1 U444 ( .A1(n40), .A2(n33), .B(n148), .X(n164) );
  SEN_OAI21_G_1 U445 ( .A1(n40), .A2(n32), .B(n148), .X(n161) );
  SEN_OAI221_1 U446 ( .A1(n80), .A2(n79), .B1(n88), .B2(n78), .C(n89), .X(
        Z[29]) );
  SEN_OA22_DG_1 U447 ( .A1(n60), .A2(n57), .B1(n61), .B2(n49), .X(n55) );
  SEN_OA22_DG_1 U448 ( .A1(n56), .A2(n57), .B1(n58), .B2(n49), .X(n54) );
  SEN_OA22_1 U449 ( .A1(n69), .A2(n46), .B1(n70), .B2(n66), .X(n61) );
  SEN_ND2_G_1 U450 ( .A1(n57), .A2(S[0]), .X(n90) );
  SEN_OAI221_1 U451 ( .A1(n33), .A2(n167), .B1(n26), .B2(n46), .C(n168), .X(
        n128) );
  SEN_AOI222_1 U452 ( .A1(n169), .A2(X[26]), .B1(n170), .B2(X[10]), .C1(X[2]), 
        .C2(n171), .X(n168) );
  SEN_ND2_G_1 U453 ( .A1(S[0]), .A2(n49), .X(n91) );
  SEN_OAI222_1 U454 ( .A1(n16), .A2(n91), .B1(n11), .B2(n90), .C1(S[0]), .C2(
        n162), .X(Z[11]) );
  SEN_OAI221_1 U455 ( .A1(n32), .A2(n167), .B1(n3), .B2(n46), .C(n183), .X(n84) );
  SEN_AOI222_1 U456 ( .A1(n169), .A2(X[27]), .B1(n170), .B2(X[11]), .C1(X[3]), 
        .C2(n171), .X(n183) );
  SEN_AO21B_1 U457 ( .A1(n160), .A2(X[22]), .B(n148), .X(n133) );
  SEN_OAI21_G_1 U458 ( .A1(S[0]), .A2(n77), .B(n24), .X(Z[31]) );
  SEN_AOI222_1 U459 ( .A1(n169), .A2(X[24]), .B1(n170), .B2(X[8]), .C1(X[0]), 
        .C2(n171), .X(n176) );
  SEN_OAI221_1 U460 ( .A1(n39), .A2(n173), .B1(n31), .B2(n174), .C(n178), .X(
        n177) );
  SEN_INV_S_1 U461 ( .A(X[12]), .X(n39) );
  SEN_OAI221_1 U462 ( .A1(n38), .A2(n173), .B1(n29), .B2(n174), .C(n182), .X(
        n181) );
  SEN_INV_S_1 U463 ( .A(X[13]), .X(n38) );
  SEN_OAI221_1 U464 ( .A1(n37), .A2(n173), .B1(n27), .B2(n174), .C(n175), .X(
        n172) );
  SEN_INV_S_1 U465 ( .A(X[14]), .X(n37) );
  SEN_INV_S_1 U466 ( .A(X[15]), .X(n36) );
  SEN_ND2_G_1 U467 ( .A1(S[0]), .A2(LEFT), .X(n191) );
  SEN_INV_S_1 U468 ( .A(X[16]), .X(n35) );
  SEN_INV_S_1 U469 ( .A(X[17]), .X(n34) );
  SEN_INV_S_1 U470 ( .A(X[18]), .X(n33) );
  SEN_INV_S_1 U471 ( .A(X[19]), .X(n32) );
  SEN_INV_S_1 U472 ( .A(X[29]), .X(n29) );
  SEN_INV_S_1 U473 ( .A(X[28]), .X(n31) );
  SEN_INV_S_1 U474 ( .A(X[30]), .X(n27) );
endmodule

