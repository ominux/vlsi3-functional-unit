
module Alu ( Z, A, B, INST, FLAGS, CLOCK );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [3:0] INST;
  output [3:0] FLAGS;
  input CLOCK;
  wire   \*Logic0* , n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774;
  wire   [31:0] A_qual;
  wire   [31:0] B_qual;
  wire   [3:0] INST_qual;
  assign FLAGS[3] = \*Logic0* ;

  SEN_FDPQ_4 \INST_qual_reg[3]  ( .D(INST[3]), .CK(CLOCK), .Q(INST_qual[3]) );
  SEN_FDPQ_4 \INST_qual_reg[2]  ( .D(INST[2]), .CK(CLOCK), .Q(INST_qual[2]) );
  SEN_FDPQ_4 \INST_qual_reg[1]  ( .D(INST[1]), .CK(CLOCK), .Q(INST_qual[1]) );
  SEN_FDPQ_4 \INST_qual_reg[0]  ( .D(INST[0]), .CK(CLOCK), .Q(INST_qual[0]) );
  SEN_FDPQ_D_1 \A_qual_reg[9]  ( .D(A[9]), .CK(CLOCK), .Q(A_qual[9]) );
  SEN_FDPQ_D_1 \A_qual_reg[8]  ( .D(A[8]), .CK(CLOCK), .Q(A_qual[8]) );
  SEN_FDPQ_D_1 \A_qual_reg[30]  ( .D(A[30]), .CK(CLOCK), .Q(A_qual[30]) );
  SEN_FDPQ_D_1 \A_qual_reg[29]  ( .D(A[29]), .CK(CLOCK), .Q(A_qual[29]) );
  SEN_FDPQ_D_1 \A_qual_reg[28]  ( .D(A[28]), .CK(CLOCK), .Q(A_qual[28]) );
  SEN_FDPQ_D_1 \A_qual_reg[27]  ( .D(A[27]), .CK(CLOCK), .Q(A_qual[27]) );
  SEN_FDPQ_D_1 \A_qual_reg[26]  ( .D(A[26]), .CK(CLOCK), .Q(A_qual[26]) );
  SEN_FDPQ_D_1 \A_qual_reg[25]  ( .D(A[25]), .CK(CLOCK), .Q(A_qual[25]) );
  SEN_FDPQ_D_1 \A_qual_reg[24]  ( .D(A[24]), .CK(CLOCK), .Q(A_qual[24]) );
  SEN_FDPQ_D_1 \A_qual_reg[23]  ( .D(A[23]), .CK(CLOCK), .Q(A_qual[23]) );
  SEN_FDPQ_D_1 \A_qual_reg[22]  ( .D(A[22]), .CK(CLOCK), .Q(A_qual[22]) );
  SEN_FDPQ_D_1 \A_qual_reg[21]  ( .D(A[21]), .CK(CLOCK), .Q(A_qual[21]) );
  SEN_FDPQ_D_1 \A_qual_reg[20]  ( .D(A[20]), .CK(CLOCK), .Q(A_qual[20]) );
  SEN_FDPQ_D_1 \A_qual_reg[19]  ( .D(A[19]), .CK(CLOCK), .Q(A_qual[19]) );
  SEN_FDPQ_D_1 \A_qual_reg[18]  ( .D(A[18]), .CK(CLOCK), .Q(A_qual[18]) );
  SEN_FDPQ_D_1 \A_qual_reg[17]  ( .D(A[17]), .CK(CLOCK), .Q(A_qual[17]) );
  SEN_FDPQ_D_1 \A_qual_reg[16]  ( .D(A[16]), .CK(CLOCK), .Q(A_qual[16]) );
  SEN_FDPQ_D_1 \A_qual_reg[14]  ( .D(A[14]), .CK(CLOCK), .Q(A_qual[14]) );
  SEN_FDPQ_D_1 \A_qual_reg[13]  ( .D(A[13]), .CK(CLOCK), .Q(A_qual[13]) );
  SEN_FDPQ_D_1 \A_qual_reg[12]  ( .D(A[12]), .CK(CLOCK), .Q(A_qual[12]) );
  SEN_FDPQ_D_1 \A_qual_reg[7]  ( .D(A[7]), .CK(CLOCK), .Q(A_qual[7]) );
  SEN_FDPQ_D_1 \A_qual_reg[5]  ( .D(A[5]), .CK(CLOCK), .Q(A_qual[5]) );
  SEN_FDPQ_D_1 \A_qual_reg[2]  ( .D(A[2]), .CK(CLOCK), .Q(A_qual[2]) );
  SEN_FDPQ_D_1 \A_qual_reg[1]  ( .D(A[1]), .CK(CLOCK), .Q(A_qual[1]) );
  SEN_FDPQ_D_1 \B_qual_reg[31]  ( .D(B[31]), .CK(CLOCK), .Q(B_qual[31]) );
  SEN_FDPQ_D_1 \B_qual_reg[30]  ( .D(B[30]), .CK(CLOCK), .Q(B_qual[30]) );
  SEN_FDPQ_D_1 \B_qual_reg[29]  ( .D(B[29]), .CK(CLOCK), .Q(B_qual[29]) );
  SEN_FDPQ_D_1 \B_qual_reg[28]  ( .D(B[28]), .CK(CLOCK), .Q(B_qual[28]) );
  SEN_FDPQ_D_1 \B_qual_reg[27]  ( .D(B[27]), .CK(CLOCK), .Q(B_qual[27]) );
  SEN_FDPQ_D_1 \B_qual_reg[26]  ( .D(B[26]), .CK(CLOCK), .Q(B_qual[26]) );
  SEN_FDPQ_D_1 \B_qual_reg[25]  ( .D(B[25]), .CK(CLOCK), .Q(B_qual[25]) );
  SEN_FDPQ_D_1 \B_qual_reg[24]  ( .D(B[24]), .CK(CLOCK), .Q(B_qual[24]) );
  SEN_FDPQ_D_1 \B_qual_reg[23]  ( .D(B[23]), .CK(CLOCK), .Q(B_qual[23]) );
  SEN_FDPQ_D_1 \B_qual_reg[22]  ( .D(B[22]), .CK(CLOCK), .Q(B_qual[22]) );
  SEN_FDPQ_D_1 \B_qual_reg[21]  ( .D(B[21]), .CK(CLOCK), .Q(B_qual[21]) );
  SEN_FDPQ_D_1 \B_qual_reg[20]  ( .D(B[20]), .CK(CLOCK), .Q(B_qual[20]) );
  SEN_FDPQ_D_1 \B_qual_reg[19]  ( .D(B[19]), .CK(CLOCK), .Q(B_qual[19]) );
  SEN_FDPQ_D_1 \B_qual_reg[18]  ( .D(B[18]), .CK(CLOCK), .Q(B_qual[18]) );
  SEN_FDPQ_D_1 \B_qual_reg[17]  ( .D(B[17]), .CK(CLOCK), .Q(B_qual[17]) );
  SEN_FDPQ_D_1 \B_qual_reg[16]  ( .D(B[16]), .CK(CLOCK), .Q(B_qual[16]) );
  SEN_FDPQ_D_1 \B_qual_reg[15]  ( .D(B[15]), .CK(CLOCK), .Q(B_qual[15]) );
  SEN_FDPQ_D_1 \B_qual_reg[14]  ( .D(B[14]), .CK(CLOCK), .Q(B_qual[14]) );
  SEN_FDPQ_D_1 \B_qual_reg[13]  ( .D(B[13]), .CK(CLOCK), .Q(B_qual[13]) );
  SEN_FDPQ_D_1 \B_qual_reg[12]  ( .D(B[12]), .CK(CLOCK), .Q(B_qual[12]) );
  SEN_FDPQ_D_1 \B_qual_reg[9]  ( .D(B[9]), .CK(CLOCK), .Q(B_qual[9]) );
  SEN_FDPQ_D_1 \B_qual_reg[7]  ( .D(B[7]), .CK(CLOCK), .Q(B_qual[7]) );
  SEN_FDPQ_D_1 \B_qual_reg[5]  ( .D(B[5]), .CK(CLOCK), .Q(B_qual[5]) );
  SEN_FDPQ_D_1 \B_qual_reg[2]  ( .D(B[2]), .CK(CLOCK), .Q(B_qual[2]) );
  SEN_FDPQ_D_1 \B_qual_reg[1]  ( .D(B[1]), .CK(CLOCK), .Q(B_qual[1]) );
  SEN_FDPQ_D_1 \B_qual_reg[6]  ( .D(B[6]), .CK(CLOCK), .Q(B_qual[6]) );
  SEN_FDPQ_D_1 \B_qual_reg[11]  ( .D(B[11]), .CK(CLOCK), .Q(B_qual[11]) );
  SEN_FDPQ_D_1 \B_qual_reg[4]  ( .D(B[4]), .CK(CLOCK), .Q(B_qual[4]) );
  SEN_FDPQ_D_1 \B_qual_reg[8]  ( .D(B[8]), .CK(CLOCK), .Q(B_qual[8]) );
  SEN_FDPQ_D_1 \B_qual_reg[3]  ( .D(B[3]), .CK(CLOCK), .Q(B_qual[3]) );
  SEN_FDPQ_D_1 \A_qual_reg[15]  ( .D(A[15]), .CK(CLOCK), .Q(A_qual[15]) );
  SEN_FDPQ_D_1 \B_qual_reg[10]  ( .D(B[10]), .CK(CLOCK), .Q(B_qual[10]) );
  SEN_FDPQ_D_1 \A_qual_reg[4]  ( .D(A[4]), .CK(CLOCK), .Q(A_qual[4]) );
  SEN_FDPQ_D_1 \A_qual_reg[0]  ( .D(A[0]), .CK(CLOCK), .Q(A_qual[0]) );
  SEN_FDPQ_D_1 \B_qual_reg[0]  ( .D(B[0]), .CK(CLOCK), .Q(B_qual[0]) );
  SEN_FDPQ_D_1 \A_qual_reg[11]  ( .D(A[11]), .CK(CLOCK), .Q(A_qual[11]) );
  SEN_FDPQ_D_1 \A_qual_reg[10]  ( .D(A[10]), .CK(CLOCK), .Q(A_qual[10]) );
  SEN_FDPQ_D_1 \A_qual_reg[6]  ( .D(A[6]), .CK(CLOCK), .Q(A_qual[6]) );
  SEN_FDPQ_D_1 \A_qual_reg[3]  ( .D(A[3]), .CK(CLOCK), .Q(A_qual[3]) );
  SEN_FDPQ_4 \A_qual_reg[31]  ( .D(A[31]), .CK(CLOCK), .Q(A_qual[31]) );
  SEN_ND2_T_1 U236 ( .A1(n756), .A2(n755), .X(n757) );
  SEN_ND2_T_3 U237 ( .A1(n272), .A2(n320), .X(n627) );
  SEN_BUF_1 U238 ( .A(n460), .X(n169) );
  SEN_MUXI2_S_2 U239 ( .D0(n259), .D1(n256), .S(B_qual[7]), .X(n305) );
  SEN_ND2_S_0P8 U240 ( .A1(n566), .A2(n565), .X(n572) );
  SEN_MUXI2_DG_4 U241 ( .D0(n227), .D1(n407), .S(A_qual[14]), .X(n320) );
  SEN_ND2_S_1P5 U242 ( .A1(n359), .A2(n485), .X(n222) );
  SEN_NR2_S_1 U243 ( .A1(n357), .A2(n486), .X(n359) );
  SEN_ND2_G_1 U244 ( .A1(n253), .A2(n509), .X(n528) );
  SEN_EN2_S_2 U245 ( .A1(n521), .A2(n523), .X(n253) );
  SEN_AOAI211_1 U246 ( .A1(n240), .A2(n501), .B(n500), .C(n553), .X(n502) );
  SEN_ND2_T_4 U247 ( .A1(n287), .A2(n288), .X(n402) );
  SEN_EO2_6 U248 ( .A1(n586), .A2(n302), .X(n589) );
  SEN_ND2_T_1 U249 ( .A1(n596), .A2(n598), .X(n328) );
  SEN_EN2_DG_1 U250 ( .A1(n254), .A2(n618), .X(n623) );
  SEN_MUXI2_S_1 U251 ( .D0(n227), .D1(n266), .S(A_qual[18]), .X(n313) );
  SEN_INV_2 U252 ( .A(n421), .X(n430) );
  SEN_INV_S_3 U253 ( .A(n447), .X(n634) );
  SEN_OA21_4 U254 ( .A1(n582), .A2(n589), .B(n592), .X(n191) );
  SEN_NR2_S_4 U255 ( .A1(n308), .A2(n307), .X(n312) );
  SEN_AN4B_2 U256 ( .B1(n580), .B2(n598), .B3(n596), .A(n472), .X(n308) );
  SEN_INV_0P8 U257 ( .A(n268), .X(n266) );
  SEN_EN2_0P5 U258 ( .A1(n245), .A2(n438), .X(n439) );
  SEN_AN2_4 U259 ( .A1(n546), .A2(n209), .X(n342) );
  SEN_AOI21B_4 U260 ( .A1(n339), .A2(n561), .B(n557), .X(n340) );
  SEN_INV_4 U261 ( .A(n625), .X(n362) );
  SEN_ND2_G_4 U262 ( .A1(n610), .A2(n606), .X(n632) );
  SEN_INV_0P65 U263 ( .A(n171), .X(n180) );
  SEN_OA21B_8 U264 ( .A1(n190), .A2(n677), .B(n172), .X(n171) );
  SEN_ND2_2 U265 ( .A1(n265), .A2(n298), .X(n600) );
  SEN_ND2_S_4 U266 ( .A1(n272), .A2(n299), .X(n599) );
  SEN_OAI21_G_4 U267 ( .A1(n312), .A2(n471), .B(n311), .X(n606) );
  SEN_OAI21_S_0P5 U268 ( .A1(n367), .A2(n366), .B(n430), .X(n170) );
  SEN_NR2_T_4 U269 ( .A1(n237), .A2(n644), .X(n367) );
  SEN_ND2_S_4 U270 ( .A1(n401), .A2(n350), .X(n290) );
  SEN_EO2_1 U271 ( .A1(n598), .A2(n597), .X(n602) );
  SEN_NR2_S_3 U272 ( .A1(Z[19]), .A2(Z[20]), .X(n766) );
  SEN_NR3_T_3 U273 ( .A1(n763), .A2(n762), .A3(Z[16]), .X(n764) );
  SEN_ND2_6 U274 ( .A1(n712), .A2(n247), .X(n726) );
  SEN_OAI21_S_8 U275 ( .A1(n396), .A2(n703), .B(n395), .X(n712) );
  SEN_ND2_S_3 U276 ( .A1(n207), .A2(n716), .X(Z[28]) );
  SEN_NR2_S_3 U277 ( .A1(n556), .A2(n558), .X(n358) );
  SEN_ND2_S_0P8 U278 ( .A1(n553), .A2(n487), .X(n556) );
  SEN_EN2_S_1 U279 ( .A1(n252), .A2(n464), .X(n465) );
  SEN_ND3_T_4 U280 ( .A1(n470), .A2(n469), .A3(n468), .X(Z[20]) );
  SEN_INV_4 U281 ( .A(n536), .X(n531) );
  SEN_NR2_2 U282 ( .A1(n529), .A2(n536), .X(n355) );
  SEN_OAI221_1 U283 ( .A1(n743), .A2(n536), .B1(n535), .B2(n212), .C(n534), 
        .X(Z[2]) );
  SEN_EN2_3 U284 ( .A1(n533), .A2(n532), .X(n536) );
  SEN_EN2_S_1 U285 ( .A1(n561), .A2(n502), .X(n508) );
  SEN_ND4_S_4 U286 ( .A1(n767), .A2(n766), .A3(n765), .A4(n764), .X(n768) );
  SEN_INV_32 U287 ( .A(n385), .X(n172) );
  SEN_AO21B_6 U288 ( .A1(n460), .A2(n461), .B(n252), .X(n371) );
  SEN_EO2_0P5 U289 ( .A1(n694), .A2(n697), .X(n696) );
  SEN_EN2_1 U290 ( .A1(n249), .A2(n489), .X(n494) );
  SEN_ND2_S_4 U291 ( .A1(n199), .A2(n249), .X(n554) );
  SEN_EO2_3 U292 ( .A1(n491), .A2(n490), .X(n249) );
  SEN_AO21B_8 U293 ( .A1(n663), .A2(n184), .B(n379), .X(n670) );
  SEN_ND3B_2 U294 ( .A(INST_qual[0]), .B1(A_qual[31]), .B2(INST_qual[2]), .X(
        n283) );
  SEN_INV_S_4 U295 ( .A(n512), .X(n423) );
  SEN_AN2_DG_1 U296 ( .A1(n572), .A2(n591), .X(n239) );
  SEN_ND2_2 U297 ( .A1(n616), .A2(n572), .X(n581) );
  SEN_NR3B_3 U298 ( .A(n580), .B1(n328), .B2(n327), .X(n343) );
  SEN_MUXI2_S_2 U299 ( .D0(n196), .D1(n407), .S(A_qual[3]), .X(n334) );
  SEN_BUF_6 U300 ( .A(n408), .X(n196) );
  SEN_ND2_S_4 U301 ( .A1(n271), .A2(n337), .X(n505) );
  SEN_MUXI2_S_1 U302 ( .D0(n259), .D1(n405), .S(B_qual[8]), .X(n295) );
  SEN_INV_5 U303 ( .A(n262), .X(n259) );
  SEN_INV_AS_10 U304 ( .A(n281), .X(n405) );
  SEN_EN2_DG_1 U305 ( .A1(n596), .A2(n584), .X(n588) );
  SEN_INV_2 U306 ( .A(n589), .X(n596) );
  SEN_OAI221_0P5 U307 ( .A1(n743), .A2(n589), .B1(n588), .B2(n212), .C(n587), 
        .X(Z[10]) );
  SEN_ND2_3 U308 ( .A1(n272), .A2(n334), .X(n540) );
  SEN_INV_S_3 U309 ( .A(n575), .X(n173) );
  SEN_INV_4 U310 ( .A(n173), .X(n174) );
  SEN_ND2_2 U311 ( .A1(n272), .A2(n296), .X(n575) );
  SEN_ND2_T_2 U312 ( .A1(n264), .A2(n336), .X(n338) );
  SEN_INV_5 U313 ( .A(n248), .X(n264) );
  SEN_MUXI2_S_2 U314 ( .D0(n260), .D1(n405), .S(B_qual[6]), .X(n336) );
  SEN_EO2_DG_2 U315 ( .A1(n441), .A2(n440), .X(n245) );
  SEN_AN2_1 U316 ( .A1(n263), .A2(n353), .X(n189) );
  SEN_ND2_3 U317 ( .A1(n272), .A2(n330), .X(n548) );
  SEN_AOI31_1 U318 ( .A1(n561), .A2(n560), .A3(n559), .B(n558), .X(n562) );
  SEN_ND2_3 U319 ( .A1(n364), .A2(n627), .X(n645) );
  SEN_EN2_S_2 U320 ( .A1(n566), .A2(n565), .X(n571) );
  SEN_ND2_S_2 U321 ( .A1(n272), .A2(n306), .X(n565) );
  SEN_ND2_S_1P5 U322 ( .A1(n272), .A2(n322), .X(n640) );
  SEN_ND2_S_1P5 U323 ( .A1(n272), .A2(n315), .X(n426) );
  SEN_MUXI2_DG_0P75 U324 ( .D0(n227), .D1(n226), .S(A_qual[17]), .X(n315) );
  SEN_ND2_6 U325 ( .A1(n272), .A2(n324), .X(n649) );
  SEN_ND2_2 U326 ( .A1(n264), .A2(n323), .X(n650) );
  SEN_ND2_T_1P5 U327 ( .A1(n407), .A2(A_qual[15]), .X(n219) );
  SEN_INV_2 U328 ( .A(n645), .X(n175) );
  SEN_INV_S_4 U329 ( .A(n175), .X(n176) );
  SEN_OAI31_3 U330 ( .A1(n554), .A2(n341), .A3(n342), .B(n340), .X(n570) );
  SEN_ND2_0P5 U331 ( .A1(n650), .A2(n649), .X(n202) );
  SEN_MUXI2_DG_0P75 U332 ( .D0(n227), .D1(n407), .S(A_qual[16]), .X(n322) );
  SEN_ND2_12 U333 ( .A1(n291), .A2(n290), .X(n407) );
  SEN_BUF_S_6 U334 ( .A(n408), .X(n227) );
  SEN_EO2_5 U335 ( .A1(n538), .A2(n540), .X(n546) );
  SEN_INV_2 U336 ( .A(n335), .X(n538) );
  SEN_ND2_S_0P5 U337 ( .A1(n445), .A2(n447), .X(n434) );
  SEN_ND3_1 U338 ( .A1(n447), .A2(n632), .A3(n241), .X(n418) );
  SEN_ND2_2 U339 ( .A1(n650), .A2(n649), .X(n447) );
  SEN_OAI21_2 U340 ( .A1(n191), .A2(n603), .B(n476), .X(n307) );
  SEN_NR2_S_2 U341 ( .A1(Z[17]), .A2(Z[18]), .X(n767) );
  SEN_ND3_1 U342 ( .A1(n444), .A2(n443), .A3(n442), .X(Z[18]) );
  SEN_NR3_T_0P5 U343 ( .A1(n591), .A2(n590), .A3(n589), .X(n594) );
  SEN_ND3_1 U344 ( .A1(n457), .A2(n456), .A3(n455), .X(Z[19]) );
  SEN_MUXI2_S_1 U345 ( .D0(n259), .D1(n405), .S(B_qual[10]), .X(n300) );
  SEN_ND2_2 U346 ( .A1(n264), .A2(n321), .X(n641) );
  SEN_MUXI2_DG_0P75 U347 ( .D0(n259), .D1(n256), .S(B_qual[16]), .X(n321) );
  SEN_ND2_S_0P5 U348 ( .A1(n176), .A2(n624), .X(n325) );
  SEN_NR2B_V1_1 U349 ( .A(n176), .B(n636), .X(n241) );
  SEN_OAI21_S_1P5 U350 ( .A1(n242), .A2(n646), .B(n176), .X(n647) );
  SEN_ND2_2 U351 ( .A1(n646), .A2(n176), .X(n417) );
  SEN_INV_6 U352 ( .A(n704), .X(n396) );
  SEN_ND2_T_5 U353 ( .A1(n726), .A2(n724), .X(n736) );
  SEN_OAI21B_4 U354 ( .A1(n747), .A2(n213), .B(n181), .X(Z[31]) );
  SEN_INV_2 U355 ( .A(n348), .X(n521) );
  SEN_OAI21_3 U356 ( .A1(n367), .A2(n366), .B(n430), .X(n435) );
  SEN_EN2_S_2 U357 ( .A1(n427), .A2(n426), .X(n421) );
  SEN_EN2_1 U358 ( .A1(n247), .A2(n712), .X(n718) );
  SEN_OAI21_S_1P5 U359 ( .A1(n239), .A2(n617), .B(n616), .X(n618) );
  SEN_ND2_6 U360 ( .A1(n617), .A2(n616), .X(n580) );
  SEN_ND2_2 U361 ( .A1(n297), .A2(n174), .X(n616) );
  SEN_INV_2 U362 ( .A(n188), .X(n262) );
  SEN_INV_4 U363 ( .A(n402), .X(n291) );
  SEN_BUF_S_1 U364 ( .A(n210), .X(n211) );
  SEN_EO2_2 U365 ( .A1(n620), .A2(n619), .X(n254) );
  SEN_EO2_1 U366 ( .A1(n454), .A2(n453), .X(n246) );
  SEN_INV_S_1 U367 ( .A(Z[10]), .X(n751) );
  SEN_ND2_T_1 U368 ( .A1(INST_qual[3]), .A2(INST_qual[0]), .X(n284) );
  SEN_ND2_S_3 U369 ( .A1(n338), .A2(n505), .X(n206) );
  SEN_INV_1 U370 ( .A(n505), .X(n204) );
  SEN_INV_2 U371 ( .A(n297), .X(n573) );
  SEN_ND2_T_1 U372 ( .A1(n272), .A2(n301), .X(n585) );
  SEN_ND2_G_1 U373 ( .A1(n254), .A2(n581), .X(n472) );
  SEN_ND2B_4 U374 ( .A(n475), .B(n361), .X(n625) );
  SEN_ND2_T_1P5 U375 ( .A1(n202), .A2(n203), .X(n416) );
  SEN_MUXI2_D_1 U376 ( .D0(n227), .D1(n407), .S(A_qual[7]), .X(n306) );
  SEN_ND2_2 U377 ( .A1(n264), .A2(n300), .X(n586) );
  SEN_INV_S_1 U378 ( .A(n211), .X(n212) );
  SEN_MUXI2_S_1 U379 ( .D0(n259), .D1(n405), .S(B_qual[11]), .X(n298) );
  SEN_EN2_3 U380 ( .A1(n600), .A2(n599), .X(n603) );
  SEN_OAI21_S_0P5 U381 ( .A1(n590), .A2(n583), .B(n582), .X(n595) );
  SEN_INV_3 U382 ( .A(n603), .X(n598) );
  SEN_ND2_2 U383 ( .A1(n233), .A2(n234), .X(n644) );
  SEN_ND2_G_1 U384 ( .A1(n641), .A2(n640), .X(n233) );
  SEN_ND2_G_1 U385 ( .A1(n231), .A2(n232), .X(n234) );
  SEN_INV_S_1 U386 ( .A(n641), .X(n231) );
  SEN_ND2_S_0P5 U387 ( .A1(n264), .A2(n318), .X(n454) );
  SEN_BUF_S_1 U388 ( .A(n695), .X(n210) );
  SEN_INV_S_1 U389 ( .A(n211), .X(n213) );
  SEN_ND2_G_1 U390 ( .A1(n264), .A2(n333), .X(n335) );
  SEN_MUXI2_S_1 U391 ( .D0(n260), .D1(n405), .S(B_qual[3]), .X(n333) );
  SEN_ND2_2 U392 ( .A1(n549), .A2(n548), .X(n487) );
  SEN_INV_S_1 U393 ( .A(n553), .X(n339) );
  SEN_ND2_T_1 U394 ( .A1(n564), .A2(n254), .X(n327) );
  SEN_ND2B_V1DG_2 U395 ( .A(n527), .B(n531), .X(n485) );
  SEN_INV_1 U396 ( .A(n364), .X(n214) );
  SEN_NR2_T_1P5 U397 ( .A1(n417), .A2(n634), .X(n365) );
  SEN_INV_2 U398 ( .A(n280), .X(n349) );
  SEN_MUXI2_S_1 U399 ( .D0(n260), .D1(n256), .S(B_qual[0]), .X(n353) );
  SEN_INV_S_1 U400 ( .A(n495), .X(n537) );
  SEN_INV_S_1 U401 ( .A(n545), .X(n486) );
  SEN_ND2_G_1 U402 ( .A1(n485), .A2(n484), .X(n495) );
  SEN_ND2_G_1 U403 ( .A1(n641), .A2(n640), .X(n445) );
  SEN_NR2_1 U404 ( .A1(n448), .A2(n636), .X(n458) );
  SEN_AO21B_4 U405 ( .A1(n435), .A2(n446), .B(n245), .X(n449) );
  SEN_EN2_0P5 U406 ( .A1(n656), .A2(n658), .X(n654) );
  SEN_ND2_G_1 U407 ( .A1(n224), .A2(n354), .X(n517) );
  SEN_MUXI2_S_1 U408 ( .D0(n196), .D1(n226), .S(A_qual[0]), .X(n354) );
  SEN_ND2_2 U409 ( .A1(n224), .A2(n347), .X(n532) );
  SEN_MUXI2_S_1 U410 ( .D0(n196), .D1(n407), .S(A_qual[2]), .X(n347) );
  SEN_ND2_G_1 U411 ( .A1(n263), .A2(n346), .X(n533) );
  SEN_EO2_2 U412 ( .A1(n189), .A2(n517), .X(n529) );
  SEN_OAI21_G_1 U413 ( .A1(n238), .A2(n546), .B(n221), .X(n547) );
  SEN_ND2_G_1 U414 ( .A1(n264), .A2(n331), .X(n491) );
  SEN_MUXI2_S_1 U415 ( .D0(n260), .D1(n405), .S(B_qual[5]), .X(n331) );
  SEN_INV_2 U416 ( .A(n341), .X(n561) );
  SEN_MUXI2_S_3 U417 ( .D0(n196), .D1(n267), .S(A_qual[6]), .X(n337) );
  SEN_NR2_T_2 U418 ( .A1(n235), .A2(n236), .X(n727) );
  SEN_OAI21_S_2 U419 ( .A1(n244), .A2(n414), .B(n413), .X(FLAGS[1]) );
  SEN_ND3_S_2 U420 ( .A1(n569), .A2(n568), .A3(n567), .X(Z[7]) );
  SEN_ND2_G_1 U421 ( .A1(n563), .A2(n210), .X(n569) );
  SEN_EO2_S_0P5 U422 ( .A1(n576), .A2(n239), .X(n579) );
  SEN_OAI211_1 U423 ( .A1(n213), .A2(n623), .B1(n622), .B2(n621), .X(Z[9]) );
  SEN_ND3_S_0P5 U424 ( .A1(n483), .A2(n482), .A3(n481), .X(Z[12]) );
  SEN_OAI211_1 U425 ( .A1(n213), .A2(n653), .B1(n652), .B2(n651), .X(Z[15]) );
  SEN_EO2_S_0P5 U426 ( .A1(n639), .A2(n638), .X(n643) );
  SEN_ND3_1 U427 ( .A1(n433), .A2(n432), .A3(n431), .X(Z[17]) );
  SEN_ND2_G_1 U428 ( .A1(n452), .A2(n210), .X(n457) );
  SEN_ND2_2 U429 ( .A1(n465), .A2(n210), .X(n470) );
  SEN_ND3_S_0P5 U430 ( .A1(n676), .A2(n675), .A3(n674), .X(Z[23]) );
  SEN_OAI21_G_1 U431 ( .A1(n711), .A2(n213), .B(n710), .X(Z[27]) );
  SEN_ND2_G_1 U432 ( .A1(n247), .A2(n274), .X(n716) );
  SEN_ND2_G_1 U433 ( .A1(n715), .A2(n714), .X(n717) );
  SEN_BUF_1 U434 ( .A(n663), .X(n177) );
  SEN_OAI21B_3 U435 ( .A1(n722), .A2(n213), .B(n178), .X(Z[29]) );
  SEN_AO31_1 U436 ( .A1(n276), .A2(n721), .A3(n720), .B(n719), .X(n178) );
  SEN_ND2_S_3 U437 ( .A1(n773), .A2(n772), .X(n774) );
  SEN_INV_S_0P5 U438 ( .A(n376), .X(n179) );
  SEN_INV_3 U439 ( .A(n268), .X(n226) );
  SEN_AN2_2 U440 ( .A1(n726), .A2(n725), .X(n235) );
  SEN_AO31_1 U441 ( .A1(n276), .A2(n746), .A3(n745), .B(n744), .X(n181) );
  SEN_BUF_3 U442 ( .A(n271), .X(n224) );
  SEN_INV_1 U443 ( .A(n273), .X(n271) );
  SEN_ND2_G_1 U444 ( .A1(n338), .A2(n505), .X(n557) );
  SEN_EO2_S_0P5 U445 ( .A1(n673), .A2(n672), .X(n182) );
  SEN_AN2_S_1 U446 ( .A1(n740), .A2(n735), .X(n183) );
  SEN_EO2_S_0P5 U447 ( .A1(n664), .A2(n666), .X(n184) );
  SEN_INV_1 U448 ( .A(n487), .X(n498) );
  SEN_INV_2 U449 ( .A(n268), .X(n225) );
  SEN_ND2_G_1 U450 ( .A1(n453), .A2(n454), .X(n461) );
  SEN_ND2_G_1 U451 ( .A1(n440), .A2(n441), .X(n459) );
  SEN_AN3_1 U452 ( .A1(n197), .A2(n545), .A3(n546), .X(n185) );
  SEN_OA31_1 U453 ( .A1(n554), .A2(n342), .A3(n341), .B(n340), .X(n186) );
  SEN_AOI21B_0P5 U454 ( .A1(n170), .A2(n446), .B(n245), .X(n187) );
  SEN_INV_2 U455 ( .A(n513), .X(n428) );
  SEN_ND2B_1 U456 ( .A(INST_qual[2]), .B(INST_qual[3]), .X(n513) );
  SEN_AN3_1 U457 ( .A1(INST_qual[1]), .A2(INST_qual[0]), .A3(n279), .X(n188)
         );
  SEN_INV_2 U458 ( .A(n546), .X(n541) );
  SEN_ND2_T_0P5 U459 ( .A1(n625), .A2(n624), .X(n636) );
  SEN_INV_1 U460 ( .A(n338), .X(n503) );
  SEN_INV_S_6 U461 ( .A(n655), .X(n376) );
  SEN_OAI21_S_1 U462 ( .A1(n499), .A2(n498), .B(n249), .X(n500) );
  SEN_ND3_S_1 U463 ( .A1(n243), .A2(n632), .A3(n458), .X(n450) );
  SEN_OAI21_T_4 U464 ( .A1(n376), .A2(n654), .B(n375), .X(n663) );
  SEN_INV_S_1 U465 ( .A(n194), .X(n257) );
  SEN_INV_S_0P5 U466 ( .A(n256), .X(n194) );
  SEN_AOI21B_8 U467 ( .A1(n670), .A2(n182), .B(n382), .X(n190) );
  SEN_NR3_T_3 U468 ( .A1(Z[24]), .A2(n768), .A3(Z[23]), .X(n769) );
  SEN_ND2_4 U469 ( .A1(n197), .A2(n198), .X(n199) );
  SEN_INV_2 U470 ( .A(n549), .X(n228) );
  SEN_EN2_S_2 U471 ( .A1(n480), .A2(n479), .X(n471) );
  SEN_ND2_G_3 U472 ( .A1(n356), .A2(n355), .X(n555) );
  SEN_ND2_T_2 U473 ( .A1(n335), .A2(n540), .X(n545) );
  SEN_ND2B_4 U474 ( .A(n607), .B(n605), .X(n475) );
  SEN_INV_2 U475 ( .A(n222), .X(n223) );
  SEN_ND2_T_2 U476 ( .A1(n204), .A2(n503), .X(n205) );
  SEN_ND2_T_2 U477 ( .A1(n264), .A2(n329), .X(n549) );
  SEN_ND2_3 U478 ( .A1(n265), .A2(n303), .X(n620) );
  SEN_BUF_1 U479 ( .A(n607), .X(n192) );
  SEN_ND2_0P65 U480 ( .A1(n348), .A2(n523), .X(n527) );
  SEN_ND2_S_1P5 U481 ( .A1(n271), .A2(n345), .X(n523) );
  SEN_MUXI2_DG_1 U482 ( .D0(n196), .D1(n407), .S(A_qual[1]), .X(n345) );
  SEN_ND2_T_1P5 U483 ( .A1(n272), .A2(n304), .X(n619) );
  SEN_MUXI2_DG_2 U484 ( .D0(n227), .D1(n407), .S(A_qual[9]), .X(n304) );
  SEN_EO2_1 U485 ( .A1(n467), .A2(n466), .X(n252) );
  SEN_INV_S_6 U486 ( .A(n262), .X(n260) );
  SEN_OAI21_S_1P5 U487 ( .A1(n244), .A2(n735), .B(n740), .X(n415) );
  SEN_INV_S_0P5 U488 ( .A(n190), .X(n193) );
  SEN_ND2_4 U489 ( .A1(n206), .A2(n205), .X(n341) );
  SEN_EO2_S_3 U490 ( .A1(n742), .A2(n741), .X(n747) );
  SEN_ND2_T_1P5 U491 ( .A1(n265), .A2(n295), .X(n297) );
  SEN_INV_2 U492 ( .A(n571), .X(n564) );
  SEN_ND2_3 U493 ( .A1(n570), .A2(n343), .X(n607) );
  SEN_MUXI2_DG_2 U494 ( .D0(n196), .D1(n407), .S(A_qual[4]), .X(n330) );
  SEN_AN2_DG_2 U495 ( .A1(n285), .A2(n423), .X(n248) );
  SEN_INV_S_4 U496 ( .A(n585), .X(n302) );
  SEN_INV_S_0P5 U497 ( .A(n228), .X(n195) );
  SEN_INV_10 U498 ( .A(n258), .X(n256) );
  SEN_INV_AS_10 U499 ( .A(n405), .X(n258) );
  SEN_OR3B_1 U500 ( .B1(n186), .B2(n571), .A(n605), .X(n591) );
  SEN_OR2_2 U501 ( .A1(n228), .A2(n548), .X(n229) );
  SEN_OAI211_1 U502 ( .A1(n692), .A2(n213), .B1(n691), .B2(n690), .X(Z[25]) );
  SEN_ND2_T_1 U503 ( .A1(n285), .A2(n284), .X(n288) );
  SEN_ND2_3 U504 ( .A1(n229), .A2(n230), .X(n251) );
  SEN_ND2_2 U505 ( .A1(n264), .A2(n305), .X(n566) );
  SEN_ND2_1P5 U506 ( .A1(n487), .A2(n545), .X(n208) );
  SEN_AOAI211_6 U507 ( .A1(n740), .A2(n739), .B(n183), .C(n738), .X(n741) );
  SEN_INV_2 U508 ( .A(Z[28]), .X(n773) );
  SEN_EO2_4 U509 ( .A1(n735), .A2(n727), .X(n734) );
  SEN_ND2_T_2 U510 ( .A1(n264), .A2(n319), .X(n364) );
  SEN_MUXI2_DG_3 U511 ( .D0(n259), .D1(n405), .S(B_qual[14]), .X(n319) );
  SEN_OR3B_4 U512 ( .B1(n737), .B2(n183), .A(n736), .X(n738) );
  SEN_AO21B_6 U513 ( .A1(n449), .A2(n459), .B(n246), .X(n460) );
  SEN_MUXI2_DG_2 U514 ( .D0(n196), .D1(n225), .S(A_qual[5]), .X(n332) );
  SEN_NR2_1 U515 ( .A1(INST_qual[0]), .A2(INST_qual[1]), .X(n286) );
  SEN_ND2_S_0P5 U516 ( .A1(n605), .A2(n604), .X(n608) );
  SEN_ND3_T_4 U517 ( .A1(n555), .A2(n358), .A3(n223), .X(n605) );
  SEN_MUXI2_DG_1 U518 ( .D0(n227), .D1(n407), .S(A_qual[8]), .X(n296) );
  SEN_MUXI2_DG_3 U519 ( .D0(n259), .D1(n256), .S(B_qual[15]), .X(n323) );
  SEN_ND2_T_1 U520 ( .A1(n227), .A2(n217), .X(n218) );
  SEN_INV_1 U521 ( .A(n649), .X(n201) );
  SEN_MUXI2_S_3 U522 ( .D0(n283), .D1(n512), .S(INST_qual[3]), .X(n408) );
  SEN_INV_S_0P5 U523 ( .A(n408), .X(n270) );
  SEN_ND2_G_3 U524 ( .A1(n214), .A2(n215), .X(n216) );
  SEN_EO2_5 U525 ( .A1(n573), .A2(n174), .X(n617) );
  SEN_INV_6 U526 ( .A(n407), .X(n268) );
  SEN_INV_0P65 U527 ( .A(INST_qual[0]), .X(n422) );
  SEN_ND2_G_1 U528 ( .A1(n586), .A2(n585), .X(n592) );
  SEN_INV_S_2 U529 ( .A(n627), .X(n215) );
  SEN_MUXI2_DG_3 U530 ( .D0(n260), .D1(n256), .S(B_qual[4]), .X(n329) );
  SEN_ND3B_1 U531 ( .A(n284), .B1(INST_qual[2]), .B2(INST_qual[1]), .X(n409)
         );
  SEN_ND2_T_2 U532 ( .A1(n218), .A2(n219), .X(n220) );
  SEN_ND2_2 U533 ( .A1(n200), .A2(n201), .X(n203) );
  SEN_ND2_3 U534 ( .A1(n645), .A2(n216), .X(n646) );
  SEN_INV_0P8 U535 ( .A(n650), .X(n200) );
  SEN_ND2_2 U536 ( .A1(n620), .A2(n619), .X(n582) );
  SEN_MUXI2_S_1 U537 ( .D0(n227), .D1(n407), .S(A_qual[11]), .X(n299) );
  SEN_INV_3 U538 ( .A(n248), .X(n265) );
  SEN_OAI21B_0P5 U539 ( .A1(n608), .A2(n192), .B(n606), .X(n609) );
  SEN_ND2_G_1 U540 ( .A1(n228), .A2(n548), .X(n230) );
  SEN_INV_2 U541 ( .A(n498), .X(n197) );
  SEN_INV_3 U542 ( .A(n251), .X(n198) );
  SEN_INV_1 U543 ( .A(n640), .X(n232) );
  SEN_NR3_T_3 U544 ( .A1(Z[27]), .A2(n771), .A3(Z[26]), .X(n772) );
  SEN_ND2_S_3 U545 ( .A1(n770), .A2(n769), .X(n771) );
  SEN_ND3_T_2 U546 ( .A1(n761), .A2(n760), .A3(n759), .X(n762) );
  SEN_NR3_T_2 U547 ( .A1(n758), .A2(n757), .A3(Z[12]), .X(n761) );
  SEN_ND2B_S_0P5 U548 ( .A(n248), .B(n377), .X(n664) );
  SEN_INV_1P25 U549 ( .A(n248), .X(n263) );
  SEN_ND4_S_0P5 U550 ( .A1(n243), .A2(n632), .A3(n459), .A4(n458), .X(n463) );
  SEN_NR3_T_2 U551 ( .A1(n326), .A2(n325), .A3(n434), .X(n363) );
  SEN_INV_1P5 U552 ( .A(n208), .X(n209) );
  SEN_MUXI2_DG_1 U553 ( .D0(n227), .D1(n407), .S(A_qual[10]), .X(n301) );
  SEN_ND2_2 U554 ( .A1(n491), .A2(n490), .X(n553) );
  SEN_AO21_2 U555 ( .A1(n416), .A2(n447), .B(n365), .X(n237) );
  SEN_OAI21_5 U556 ( .A1(n428), .A2(n349), .B(n422), .X(n281) );
  SEN_ND2B_V1DG_1 U557 ( .A(INST_qual[2]), .B(INST_qual[1]), .X(n280) );
  SEN_OA21_2 U558 ( .A1(n718), .A2(n213), .B(n717), .X(n207) );
  SEN_AOI21B_1 U559 ( .A1(n463), .A2(n462), .B(n461), .X(n464) );
  SEN_MUXI2_DG_3 U560 ( .D0(n423), .D1(n286), .S(INST_qual[3]), .X(n287) );
  SEN_MUXI2_DG_2 U561 ( .D0(n259), .D1(n256), .S(B_qual[9]), .X(n303) );
  SEN_EO2_G_2 U562 ( .A1(n737), .A2(n736), .X(n722) );
  SEN_OAI21_S_8 U563 ( .A1(n372), .A2(n371), .B(n370), .X(n655) );
  SEN_OAI221_1 U564 ( .A1(n743), .A2(n644), .B1(n643), .B2(n213), .C(n642), 
        .X(Z[16]) );
  SEN_NR4_3 U565 ( .A1(Z[31]), .A2(Z[30]), .A3(n774), .A4(Z[29]), .X(FLAGS[2])
         );
  SEN_ND2_T_1 U566 ( .A1(n272), .A2(n317), .X(n453) );
  SEN_INV_S_1P5 U567 ( .A(n445), .X(n366) );
  SEN_ND2_T_1 U568 ( .A1(n272), .A2(n313), .X(n440) );
  SEN_OAI21_S_8 U569 ( .A1(n392), .A2(n693), .B(n391), .X(n704) );
  SEN_INV_6 U570 ( .A(n694), .X(n392) );
  SEN_ND2_0P8 U571 ( .A1(n426), .A2(n427), .X(n446) );
  SEN_ND2_T_0P5 U572 ( .A1(n263), .A2(n373), .X(n656) );
  SEN_EN2_0P5 U573 ( .A1(n253), .A2(n250), .X(n526) );
  SEN_ND2_S_0P5 U574 ( .A1(n253), .A2(n275), .X(n524) );
  SEN_AOAI211_0P5 U575 ( .A1(n510), .A2(n529), .B(n250), .C(n210), .X(n520) );
  SEN_AN2_1 U576 ( .A1(n509), .A2(n511), .X(n250) );
  SEN_NR3_0P65 U577 ( .A1(n486), .A2(n495), .A3(n496), .X(n488) );
  SEN_ND2_G_1 U578 ( .A1(n272), .A2(n310), .X(n479) );
  SEN_OAI21_S_1 U579 ( .A1(n488), .A2(n497), .B(n197), .X(n489) );
  SEN_INV_1 U580 ( .A(n484), .X(n357) );
  SEN_ND2_G_1 U581 ( .A1(n533), .A2(n532), .X(n484) );
  SEN_OAI21_S_8 U582 ( .A1(n171), .A2(n685), .B(n388), .X(n694) );
  SEN_AOI21B_2 U583 ( .A1(n437), .A2(n436), .B(n446), .X(n438) );
  SEN_NR3_T_1 U584 ( .A1(Z[2]), .A2(Z[0]), .A3(Z[1]), .X(n752) );
  SEN_EO2_0P5 U585 ( .A1(n182), .A2(n670), .X(n671) );
  SEN_ND2_G_1 U586 ( .A1(n264), .A2(n316), .X(n427) );
  SEN_MUXI2_S_1 U587 ( .D0(n260), .D1(n405), .S(B_qual[1]), .X(n344) );
  SEN_INV_0P65 U588 ( .A(n557), .X(n558) );
  SEN_EN2_0P5 U589 ( .A1(n184), .A2(n177), .X(n669) );
  SEN_NR3_T_2 U590 ( .A1(Z[9]), .A2(Z[11]), .A3(Z[13]), .X(n760) );
  SEN_OAI21_T_4 U591 ( .A1(n734), .A2(n213), .B(n733), .X(Z[30]) );
  SEN_AOI211_G_1 U592 ( .A1(n596), .A2(n595), .B1(n594), .B2(n593), .X(n597)
         );
  SEN_EN2_DG_1 U593 ( .A1(n251), .A2(n547), .X(n552) );
  SEN_EN2_S_1 U594 ( .A1(n246), .A2(n451), .X(n452) );
  SEN_ND3_S_1 U595 ( .A1(n459), .A2(n446), .A3(n461), .X(n326) );
  SEN_NR3_T_2 U596 ( .A1(Z[7]), .A2(n754), .A3(Z[4]), .X(n755) );
  SEN_EN2_S_1 U597 ( .A1(n564), .A2(n562), .X(n563) );
  SEN_AOI21_S_0P5 U598 ( .A1(n447), .A2(n633), .B(n644), .X(n419) );
  SEN_ND2_G_1 U599 ( .A1(n254), .A2(n580), .X(n590) );
  SEN_ND2_G_1 U600 ( .A1(INST_qual[3]), .A2(INST_qual[2]), .X(n279) );
  SEN_ND2B_3 U601 ( .A(INST_qual[1]), .B(INST_qual[0]), .X(n512) );
  SEN_INV_2 U602 ( .A(n409), .X(n273) );
  SEN_INV_1P5 U603 ( .A(n268), .X(n267) );
  SEN_EN2_0P5 U604 ( .A1(n689), .A2(n180), .X(n692) );
  SEN_ND2_2 U605 ( .A1(n272), .A2(n332), .X(n490) );
  SEN_OR3B_1 U606 ( .B1(INST_qual[0]), .B2(A_qual[31]), .A(INST_qual[2]), .X(
        n289) );
  SEN_INV_S_1 U607 ( .A(A_qual[15]), .X(n217) );
  SEN_INV_3 U608 ( .A(n220), .X(n324) );
  SEN_INV_S_0P5 U609 ( .A(n486), .X(n221) );
  SEN_OA21_4 U610 ( .A1(n399), .A2(n737), .B(n739), .X(n244) );
  SEN_EO2_S_1 U611 ( .A1(FLAGS[1]), .A2(n415), .X(FLAGS[0]) );
  SEN_ND2_S_0P5 U612 ( .A1(n176), .A2(n632), .X(n637) );
  SEN_INV_S_1 U613 ( .A(n633), .X(n635) );
  SEN_ND2_S_0P5 U614 ( .A1(n251), .A2(n275), .X(n551) );
  SEN_ND2_G_1 U615 ( .A1(n648), .A2(n417), .X(n633) );
  SEN_EN2_S_1 U616 ( .A1(n648), .A2(n647), .X(n653) );
  SEN_ND2_S_0P5 U617 ( .A1(n689), .A2(n274), .X(n690) );
  SEN_INV_4 U618 ( .A(n273), .X(n272) );
  SEN_INV_S_0P5 U619 ( .A(n555), .X(n496) );
  SEN_NR2B_V1_1 U620 ( .A(n276), .B(n521), .X(n522) );
  SEN_NR2_S_0P5 U621 ( .A1(n743), .A2(n742), .X(n744) );
  SEN_NR2_S_0P5 U622 ( .A1(n743), .A2(n737), .X(n719) );
  SEN_NR2B_V1DG_1 U623 ( .A(n276), .B(n729), .X(n730) );
  SEN_NR2B_V1DG_1 U624 ( .A(n276), .B(n706), .X(n707) );
  SEN_INV_S_0P5 U625 ( .A(INST_qual[2]), .X(n285) );
  SEN_AN2_S_0P5 U626 ( .A1(n555), .A2(n537), .X(n238) );
  SEN_NR2_S_0P5 U627 ( .A1(n496), .A2(n498), .X(n501) );
  SEN_INV_S_1 U628 ( .A(n497), .X(n499) );
  SEN_INV_S_0P5 U629 ( .A(n360), .X(n610) );
  SEN_INV_1 U630 ( .A(n528), .X(n356) );
  SEN_INV_S_0P5 U631 ( .A(n416), .X(n648) );
  SEN_INV_S_0P5 U632 ( .A(n617), .X(n576) );
  SEN_INV_S_0P5 U633 ( .A(n644), .X(n639) );
  SEN_ND2_S_0P5 U634 ( .A1(n600), .A2(n599), .X(n476) );
  SEN_AN2_S_1 U635 ( .A1(n739), .A2(n737), .X(n236) );
  SEN_ND3B_V1DG_1 U636 ( .A(n556), .B1(n555), .B2(n240), .X(n559) );
  SEN_ND3B_0P5 U637 ( .A(n434), .B1(n632), .B2(n241), .X(n437) );
  SEN_OAOI211_1 U638 ( .A1(n637), .A2(n636), .B(n635), .C(n634), .X(n638) );
  SEN_INV_S_0P5 U639 ( .A(n581), .X(n583) );
  SEN_ND2_S_1 U640 ( .A1(n753), .A2(n752), .X(n754) );
  SEN_OAI21_S_0P5 U641 ( .A1(n541), .A2(n486), .B(n251), .X(n497) );
  SEN_ND2_S_1 U642 ( .A1(n749), .A2(n748), .X(n763) );
  SEN_ND2_S_0P5 U643 ( .A1(n176), .A2(n447), .X(n448) );
  SEN_INV_S_0P5 U644 ( .A(n471), .X(n604) );
  SEN_INV_S_0P5 U645 ( .A(n529), .X(n511) );
  SEN_AN3_0P5 U646 ( .A1(n624), .A2(n632), .A3(n625), .X(n242) );
  SEN_NR2B_V1DG_1 U647 ( .A(n276), .B(n538), .X(n539) );
  SEN_AN2_S_0P5 U648 ( .A1(n221), .A2(n537), .X(n240) );
  SEN_AN2_S_0P5 U649 ( .A1(n446), .A2(n445), .X(n243) );
  SEN_OAI21_S_0P5 U650 ( .A1(n423), .A2(n422), .B(n428), .X(n695) );
  SEN_ND2_S_0P5 U651 ( .A1(n610), .A2(n274), .X(n614) );
  SEN_ND2_S_0P5 U652 ( .A1(n648), .A2(n274), .X(n652) );
  SEN_ND2_S_0P5 U653 ( .A1(n666), .A2(n665), .X(n668) );
  SEN_ND2_S_0P5 U654 ( .A1(n254), .A2(n274), .X(n622) );
  SEN_ND2_S_0P5 U655 ( .A1(n576), .A2(n274), .X(n577) );
  SEN_ND2_S_0P5 U656 ( .A1(n249), .A2(n275), .X(n493) );
  SEN_ND2_S_0P5 U657 ( .A1(n658), .A2(n656), .X(n375) );
  SEN_INV_S_0P5 U658 ( .A(n425), .X(n277) );
  SEN_ND2_S_0P5 U659 ( .A1(n523), .A2(n522), .X(n525) );
  SEN_ND2_S_0P5 U660 ( .A1(n658), .A2(n657), .X(n661) );
  SEN_ND2_S_0P5 U661 ( .A1(n541), .A2(n275), .X(n542) );
  SEN_ND2_S_0P5 U662 ( .A1(n627), .A2(n626), .X(n630) );
  SEN_ND2_S_0P5 U663 ( .A1(n561), .A2(n275), .X(n506) );
  SEN_ND2_S_0P5 U664 ( .A1(n604), .A2(n275), .X(n482) );
  SEN_ND2_S_0P5 U665 ( .A1(n245), .A2(n275), .X(n443) );
  SEN_INV_S_0P5 U666 ( .A(n262), .X(n261) );
  SEN_ND2_S_0P5 U667 ( .A1(n480), .A2(n479), .X(n311) );
  SEN_EN2_S_1 U668 ( .A1(n612), .A2(n611), .X(n360) );
  SEN_INV_S_0P5 U669 ( .A(n270), .X(n269) );
  SEN_NR2B_V1_1 U670 ( .A(n276), .B(n189), .X(n516) );
  SEN_ND2_S_0P5 U671 ( .A1(n466), .A2(n467), .X(n370) );
  SEN_INV_S_0P5 U672 ( .A(n509), .X(n510) );
  SEN_AN2_S_0P5 U673 ( .A1(n276), .A2(n364), .X(n626) );
  SEN_AN2_S_0P5 U674 ( .A1(n276), .A2(n656), .X(n657) );
  SEN_AN2_S_0P5 U675 ( .A1(n276), .A2(n664), .X(n665) );
  SEN_AN2_S_0P5 U676 ( .A1(n276), .A2(n678), .X(n679) );
  SEN_AN2_S_0P5 U677 ( .A1(n276), .A2(n686), .X(n687) );
  SEN_AN2_S_0P5 U678 ( .A1(n276), .A2(n713), .X(n714) );
  SEN_ND2_S_0P5 U679 ( .A1(n672), .A2(n673), .X(n382) );
  SEN_INV_S_0P5 U680 ( .A(n425), .X(n278) );
  SEN_MUXI2_S_0P5 U681 ( .D0(n227), .D1(n266), .S(A_qual[19]), .X(n317) );
  SEN_MUXI2_S_0P5 U682 ( .D0(n227), .D1(n226), .S(A_qual[12]), .X(n310) );
  SEN_OR3B_0P5 U683 ( .B1(n429), .B2(INST_qual[0]), .A(n428), .X(n743) );
  SEN_INV_S_0P5 U684 ( .A(INST_qual[1]), .X(n429) );
  SEN_ND2_S_0P5 U685 ( .A1(n264), .A2(n314), .X(n441) );
  SEN_MUXI2_S_0P5 U686 ( .D0(n259), .D1(n405), .S(B_qual[18]), .X(n314) );
  SEN_ND3_S_0P5 U687 ( .A1(n265), .A2(n352), .A3(n351), .X(n509) );
  SEN_ND2_S_0P5 U688 ( .A1(n264), .A2(n406), .X(n728) );
  SEN_ND2_S_0P5 U689 ( .A1(n224), .A2(n398), .X(n720) );
  SEN_MUXI2_S_0P5 U690 ( .D0(n269), .D1(n266), .S(A_qual[29]), .X(n398) );
  SEN_ND2_S_0P5 U691 ( .A1(n224), .A2(n394), .X(n708) );
  SEN_MUXI2_S_0P5 U692 ( .D0(n269), .D1(n225), .S(A_qual[27]), .X(n394) );
  SEN_ND2_S_0P5 U693 ( .A1(n224), .A2(n404), .X(n745) );
  SEN_ND2_S_0P5 U694 ( .A1(n224), .A2(n374), .X(n658) );
  SEN_MUXI2_S_0P5 U695 ( .D0(n196), .D1(n226), .S(A_qual[21]), .X(n374) );
  SEN_ND2_S_0P5 U696 ( .A1(n224), .A2(n378), .X(n666) );
  SEN_MUXI2_S_0P5 U697 ( .D0(n196), .D1(n225), .S(A_qual[22]), .X(n378) );
  SEN_ND2_S_0P5 U698 ( .A1(n224), .A2(n384), .X(n680) );
  SEN_MUXI2_S_0P5 U699 ( .D0(n196), .D1(n266), .S(A_qual[24]), .X(n384) );
  SEN_ND2_S_0P5 U700 ( .A1(n224), .A2(n387), .X(n688) );
  SEN_MUXI2_S_0P5 U701 ( .D0(n196), .D1(n226), .S(A_qual[25]), .X(n387) );
  SEN_ND2_S_0P5 U702 ( .A1(n264), .A2(n309), .X(n480) );
  SEN_MUXI2_S_0P5 U703 ( .D0(n259), .D1(n405), .S(B_qual[12]), .X(n309) );
  SEN_MUXI2_S_0P5 U704 ( .D0(n259), .D1(n405), .S(B_qual[17]), .X(n316) );
  SEN_MUXI2_S_0P5 U705 ( .D0(n259), .D1(n405), .S(B_qual[19]), .X(n318) );
  SEN_ND2_S_0P5 U706 ( .A1(n263), .A2(n282), .X(n713) );
  SEN_MUXI2_S_0P5 U707 ( .D0(n259), .D1(n257), .S(B_qual[28]), .X(n282) );
  SEN_ND2_S_0P5 U708 ( .A1(n224), .A2(n369), .X(n466) );
  SEN_MUXI2_S_0P5 U709 ( .D0(n196), .D1(n226), .S(A_qual[20]), .X(n369) );
  SEN_ND2_S_0P5 U710 ( .A1(n263), .A2(n386), .X(n686) );
  SEN_MUXI2_S_0P5 U711 ( .D0(n260), .D1(n257), .S(B_qual[25]), .X(n386) );
  SEN_ND2_S_0P5 U712 ( .A1(n224), .A2(n381), .X(n672) );
  SEN_MUXI2_S_0P5 U713 ( .D0(n196), .D1(n266), .S(A_qual[23]), .X(n381) );
  SEN_ND2_S_0P5 U714 ( .A1(n224), .A2(n390), .X(n698) );
  SEN_MUXI2_S_0P5 U715 ( .D0(n196), .D1(n225), .S(A_qual[26]), .X(n390) );
  SEN_ND2_S_0P5 U716 ( .A1(n410), .A2(n224), .X(n731) );
  SEN_MUXI2_S_0P5 U717 ( .D0(n269), .D1(n266), .S(A_qual[30]), .X(n410) );
  SEN_ND2_S_0P5 U718 ( .A1(n263), .A2(n368), .X(n467) );
  SEN_MUXI2_S_0P5 U719 ( .D0(n260), .D1(n256), .S(B_qual[20]), .X(n368) );
  SEN_ND2_S_0P5 U720 ( .A1(n263), .A2(n393), .X(n705) );
  SEN_ND2_S_0P5 U721 ( .A1(n263), .A2(n400), .X(n746) );
  SEN_MUXI2_S_0P5 U722 ( .D0(n260), .D1(n257), .S(B_qual[21]), .X(n373) );
  SEN_MUXI2_S_0P5 U723 ( .D0(n260), .D1(n257), .S(B_qual[22]), .X(n377) );
  SEN_ND2_S_0P5 U724 ( .A1(n263), .A2(n383), .X(n678) );
  SEN_MUXI2_S_0P5 U725 ( .D0(n260), .D1(n257), .S(B_qual[24]), .X(n383) );
  SEN_ND2_S_0P5 U726 ( .A1(n263), .A2(n380), .X(n673) );
  SEN_MUXI2_S_0P5 U727 ( .D0(n260), .D1(n257), .S(B_qual[23]), .X(n380) );
  SEN_ND2_S_0P5 U728 ( .A1(n263), .A2(n389), .X(n699) );
  SEN_MUXI2_S_0P5 U729 ( .D0(n260), .D1(n257), .S(B_qual[26]), .X(n389) );
  SEN_ND2_S_0P5 U730 ( .A1(n263), .A2(n397), .X(n721) );
  SEN_ND2_S_0P5 U731 ( .A1(n271), .A2(n292), .X(n715) );
  SEN_MUXI2_S_0P5 U732 ( .D0(n227), .D1(n226), .S(A_qual[28]), .X(n292) );
  SEN_MUXI2_S_0P5 U733 ( .D0(n227), .D1(n226), .S(A_qual[13]), .X(n294) );
  SEN_MUXI2_S_0P5 U734 ( .D0(n259), .D1(n405), .S(B_qual[13]), .X(n293) );
  SEN_INV_S_0P5 U735 ( .A(INST_qual[3]), .X(n401) );
  SEN_INV_S_2 U736 ( .A(n289), .X(n350) );
  SEN_OR2_DG_1 U737 ( .A1(A_qual[0]), .A2(B_qual[0]), .X(n514) );
  SEN_OR3B_0P5 U738 ( .B1(INST_qual[1]), .B2(INST_qual[0]), .A(n428), .X(n425)
         );
  SEN_OAI21B_1 U739 ( .A1(n590), .A2(n591), .B(n595), .X(n584) );
  SEN_AOI21B_1 U740 ( .A1(n450), .A2(n187), .B(n459), .X(n451) );
  SEN_EN2_0P5 U741 ( .A1(n604), .A2(n477), .X(n478) );
  SEN_NR2B_1 U742 ( .A(n724), .B(n723), .X(n725) );
  SEN_INV_S_1 U743 ( .A(n739), .X(n723) );
  SEN_EO2_S_0P5 U744 ( .A1(n421), .A2(n420), .X(n424) );
  SEN_AOI21B_1 U745 ( .A1(n419), .A2(n418), .B(n445), .X(n420) );
  SEN_INV_S_1 U746 ( .A(n735), .X(n732) );
  SEN_INV_S_1 U747 ( .A(n685), .X(n689) );
  SEN_INV_S_1 U748 ( .A(n703), .X(n709) );
  SEN_INV_S_1 U749 ( .A(n654), .X(n659) );
  SEN_INV_S_1 U750 ( .A(n677), .X(n681) );
  SEN_INV_S_1 U751 ( .A(Z[21]), .X(n749) );
  SEN_INV_S_1 U752 ( .A(n742), .X(n411) );
  SEN_INV_S_1 U753 ( .A(Z[3]), .X(n753) );
  SEN_NR2B_V1_1 U754 ( .A(n276), .B(n503), .X(n504) );
  SEN_NR2B_1 U755 ( .A(n276), .B(n573), .X(n574) );
  SEN_INV_S_1 U756 ( .A(n693), .X(n697) );
  SEN_ND2_S_1 U757 ( .A1(n751), .A2(n750), .X(n758) );
  SEN_NR2_S_1 U758 ( .A1(Z[5]), .A2(Z[6]), .X(n756) );
  SEN_NR2_1 U759 ( .A1(n360), .A2(n471), .X(n361) );
  SEN_INV_S_1 U760 ( .A(Z[25]), .X(n770) );
  SEN_INV_S_1 U761 ( .A(Z[14]), .X(n759) );
  SEN_INV_S_1 U762 ( .A(Z[15]), .X(n748) );
  SEN_INV_S_1 U763 ( .A(Z[8]), .X(n750) );
  SEN_INV_S_1 U764 ( .A(Z[22]), .X(n765) );
  SEN_INV_S_1 U765 ( .A(n743), .X(n274) );
  SEN_INV_S_1 U766 ( .A(n743), .X(n275) );
  SEN_ND3_S_0P5 U767 ( .A1(n277), .A2(n600), .A3(n599), .X(n601) );
  SEN_ND2_G_1 U768 ( .A1(n680), .A2(n679), .X(n683) );
  SEN_ND2_G_1 U769 ( .A1(n681), .A2(n274), .X(n682) );
  SEN_EN2_0P5 U770 ( .A1(n681), .A2(n193), .X(n684) );
  SEN_EN2_0P5 U771 ( .A1(n728), .A2(n731), .X(n735) );
  SEN_EN2_0P5 U772 ( .A1(n746), .A2(n745), .X(n742) );
  SEN_EN2_0P5 U773 ( .A1(n721), .A2(n720), .X(n737) );
  SEN_ND3_S_0P5 U774 ( .A1(n277), .A2(n641), .A3(n640), .X(n642) );
  SEN_EN2_0P5 U775 ( .A1(n686), .A2(n688), .X(n685) );
  SEN_EN2_0P5 U776 ( .A1(n678), .A2(n680), .X(n677) );
  SEN_EN2_0P5 U777 ( .A1(n705), .A2(n708), .X(n703) );
  SEN_EN2_0P5 U778 ( .A1(n699), .A2(n698), .X(n693) );
  SEN_OAI211_1 U779 ( .A1(n212), .A2(n552), .B1(n551), .B2(n550), .X(Z[4]) );
  SEN_ND3_S_0P5 U780 ( .A1(n277), .A2(n195), .A3(n548), .X(n550) );
  SEN_OAI211_1 U781 ( .A1(n213), .A2(n615), .B1(n614), .B2(n613), .X(Z[13]) );
  SEN_ND3_S_0P5 U782 ( .A1(n277), .A2(n612), .A3(n611), .X(n613) );
  SEN_EN2_0P5 U783 ( .A1(n610), .A2(n609), .X(n615) );
  SEN_OAI211_1 U784 ( .A1(n526), .A2(n212), .B1(n525), .B2(n524), .X(Z[1]) );
  SEN_ND3_S_0P5 U785 ( .A1(n277), .A2(n533), .A3(n532), .X(n534) );
  SEN_EN2_0P5 U786 ( .A1(n531), .A2(n530), .X(n535) );
  SEN_OAI21_S_0P5 U787 ( .A1(n529), .A2(n528), .B(n527), .X(n530) );
  SEN_OAI211_1 U788 ( .A1(n508), .A2(n212), .B1(n507), .B2(n506), .X(Z[6]) );
  SEN_ND2_G_1 U789 ( .A1(n505), .A2(n504), .X(n507) );
  SEN_ND2_G_1 U790 ( .A1(n731), .A2(n728), .X(n740) );
  SEN_ND2_G_1 U791 ( .A1(n708), .A2(n705), .X(n395) );
  SEN_ND3_S_0P5 U792 ( .A1(n277), .A2(n620), .A3(n619), .X(n621) );
  SEN_OAI211_1 U793 ( .A1(n212), .A2(n494), .B1(n493), .B2(n492), .X(Z[5]) );
  SEN_ND3_S_0P5 U794 ( .A1(n277), .A2(n491), .A3(n490), .X(n492) );
  SEN_ND2_G_1 U795 ( .A1(n720), .A2(n721), .X(n739) );
  SEN_OAI211_1 U796 ( .A1(n544), .A2(n212), .B1(n543), .B2(n542), .X(Z[3]) );
  SEN_EO2_S_0P5 U797 ( .A1(n541), .A2(n238), .X(n544) );
  SEN_ND3_S_0P5 U798 ( .A1(n277), .A2(n650), .A3(n649), .X(n651) );
  SEN_OAI211_1 U799 ( .A1(n631), .A2(n213), .B1(n630), .B2(n629), .X(Z[14]) );
  SEN_ND2_G_1 U800 ( .A1(n628), .A2(n274), .X(n629) );
  SEN_EO2_S_0P5 U801 ( .A1(n628), .A2(n242), .X(n631) );
  SEN_ND2_G_1 U802 ( .A1(n698), .A2(n699), .X(n391) );
  SEN_OAI211_1 U803 ( .A1(n579), .A2(n212), .B1(n578), .B2(n577), .X(Z[8]) );
  SEN_ND2_G_1 U804 ( .A1(n174), .A2(n574), .X(n578) );
  SEN_OAI211_1 U805 ( .A1(n662), .A2(n213), .B1(n661), .B2(n660), .X(Z[21]) );
  SEN_ND2_G_1 U806 ( .A1(n659), .A2(n274), .X(n660) );
  SEN_EN2_0P5 U807 ( .A1(n659), .A2(n179), .X(n662) );
  SEN_OAI211_1 U808 ( .A1(n669), .A2(n213), .B1(n668), .B2(n667), .X(Z[22]) );
  SEN_ND2_G_1 U809 ( .A1(n184), .A2(n274), .X(n667) );
  SEN_ND2_G_1 U810 ( .A1(n688), .A2(n687), .X(n691) );
  SEN_ND2_G_1 U811 ( .A1(n680), .A2(n678), .X(n385) );
  SEN_EO2_S_0P5 U812 ( .A1(n713), .A2(n715), .X(n247) );
  SEN_ND3_S_0P5 U813 ( .A1(n520), .A2(n519), .A3(n518), .X(Z[0]) );
  SEN_AOI22_0P5 U814 ( .A1(n517), .A2(n516), .B1(n515), .B2(n514), .X(n518) );
  SEN_ND2_G_1 U815 ( .A1(n511), .A2(n275), .X(n519) );
  SEN_ND2_G_1 U816 ( .A1(n715), .A2(n713), .X(n724) );
  SEN_ND2_G_1 U817 ( .A1(n688), .A2(n686), .X(n388) );
  SEN_AOI21_S_1 U818 ( .A1(n746), .A2(n745), .B(n412), .X(n413) );
  SEN_ND2_G_1 U819 ( .A1(n411), .A2(n732), .X(n414) );
  SEN_NR2_1 U820 ( .A1(n742), .A2(n740), .X(n412) );
  SEN_ND3_S_0P5 U821 ( .A1(n277), .A2(n441), .A3(n440), .X(n442) );
  SEN_ND2_G_1 U822 ( .A1(n439), .A2(n210), .X(n444) );
  SEN_ND3_S_0P5 U823 ( .A1(n278), .A2(n467), .A3(n466), .X(n468) );
  SEN_ND2_G_1 U824 ( .A1(n252), .A2(n275), .X(n469) );
  SEN_ND3_S_1 U825 ( .A1(n702), .A2(n701), .A3(n700), .X(Z[26]) );
  SEN_ND3_S_0P5 U826 ( .A1(n277), .A2(n699), .A3(n698), .X(n700) );
  SEN_ND2_G_1 U827 ( .A1(n697), .A2(n274), .X(n701) );
  SEN_ND2_G_1 U828 ( .A1(n696), .A2(n210), .X(n702) );
  SEN_ND3_S_0P5 U829 ( .A1(n277), .A2(n673), .A3(n672), .X(n674) );
  SEN_ND2_G_1 U830 ( .A1(n182), .A2(n274), .X(n675) );
  SEN_ND2_G_1 U831 ( .A1(n671), .A2(n210), .X(n676) );
  SEN_ND3_S_0P5 U832 ( .A1(n277), .A2(n480), .A3(n479), .X(n481) );
  SEN_ND2_G_1 U833 ( .A1(n478), .A2(n210), .X(n483) );
  SEN_ND2_G_1 U834 ( .A1(n666), .A2(n664), .X(n379) );
  SEN_AOI22_1 U835 ( .A1(n709), .A2(n274), .B1(n708), .B2(n707), .X(n710) );
  SEN_EN2_0P5 U836 ( .A1(n704), .A2(n709), .X(n711) );
  SEN_ND3_S_0P5 U837 ( .A1(n277), .A2(n566), .A3(n565), .X(n567) );
  SEN_ND2_G_1 U838 ( .A1(n564), .A2(n275), .X(n568) );
  SEN_AOI22_1 U839 ( .A1(n732), .A2(n274), .B1(n731), .B2(n730), .X(n733) );
  SEN_ND3_S_0P5 U840 ( .A1(n278), .A2(n454), .A3(n453), .X(n455) );
  SEN_ND2_G_1 U841 ( .A1(n246), .A2(n275), .X(n456) );
  SEN_ND3_S_0P5 U842 ( .A1(n277), .A2(n427), .A3(n426), .X(n432) );
  SEN_ND2_G_1 U843 ( .A1(n430), .A2(n274), .X(n431) );
  SEN_ND2_G_1 U844 ( .A1(n424), .A2(n210), .X(n433) );
  SEN_ND2_G_1 U845 ( .A1(n612), .A2(n611), .X(n624) );
  SEN_INV_S_1 U846 ( .A(n705), .X(n706) );
  SEN_INV_S_1 U847 ( .A(n728), .X(n729) );
  SEN_INV_S_1 U848 ( .A(n425), .X(n276) );
  SEN_MUXI2_S_1 U849 ( .D0(n261), .D1(n257), .S(B_qual[27]), .X(n393) );
  SEN_ND2_S_0P5 U850 ( .A1(n422), .A2(n349), .X(n352) );
  SEN_MUXI2_S_1 U851 ( .D0(n261), .D1(n257), .S(B_qual[29]), .X(n397) );
  SEN_MUXI2_S_0P5 U852 ( .D0(n403), .D1(n402), .S(A_qual[31]), .X(n404) );
  SEN_MUXI2_S_1 U853 ( .D0(n261), .D1(n257), .S(B_qual[31]), .X(n400) );
  SEN_MUXI2_S_1 U854 ( .D0(n261), .D1(n257), .S(B_qual[30]), .X(n406) );
  SEN_ND2_G_1 U855 ( .A1(n224), .A2(n294), .X(n611) );
  SEN_ND2_G_1 U856 ( .A1(n265), .A2(n293), .X(n612) );
  SEN_MUXI2_S_1 U857 ( .D0(n260), .D1(n405), .S(B_qual[2]), .X(n346) );
  SEN_ND2_G_1 U858 ( .A1(n263), .A2(n344), .X(n348) );
  SEN_TIE0_1 U859 ( .X(\*Logic0* ) );
  SEN_OAI211_1 U860 ( .A1(n684), .A2(n213), .B1(n683), .B2(n682), .X(Z[24]) );
  SEN_INV_S_0P5 U861 ( .A(n302), .X(n255) );
  SEN_AN3B_0P5 U862 ( .B1(n475), .B2(n476), .A(n474), .X(n477) );
  SEN_ND2_S_0P5 U863 ( .A1(n580), .A2(n596), .X(n473) );
  SEN_OAI221_1 U864 ( .A1(n743), .A2(n603), .B1(n602), .B2(n213), .C(n601), 
        .X(Z[11]) );
  SEN_INV_S_1 U865 ( .A(n592), .X(n593) );
  SEN_ND3_S_0P5 U866 ( .A1(n277), .A2(n586), .A3(n255), .X(n587) );
  SEN_INV_S_0P5 U867 ( .A(n169), .X(n462) );
  SEN_INV_S_0P5 U868 ( .A(n646), .X(n628) );
  SEN_OAOI211_0P5 U869 ( .A1(n473), .A2(n472), .B(n191), .C(n603), .X(n474) );
  SEN_INV_S_3 U870 ( .A(n736), .X(n399) );
  SEN_OAI21_S_0P5 U871 ( .A1(n185), .A2(n554), .B(n553), .X(n560) );
  SEN_NR2_S_0P5 U872 ( .A1(n513), .A2(n512), .X(n515) );
  SEN_NR2_S_0P5 U873 ( .A1(n512), .A2(n401), .X(n403) );
  SEN_INV_S_0P5 U874 ( .A(n170), .X(n436) );
  SEN_NR2_S_0P5 U875 ( .A1(n350), .A2(INST_qual[3]), .X(n351) );
  SEN_ND2_S_0P5 U876 ( .A1(n540), .A2(n539), .X(n543) );
  SEN_AN3B_4 U877 ( .B1(n632), .B2(n363), .A(n362), .X(n372) );
endmodule

