
module Alu ( Z, A, B, DI, DO, CI, INST, FLAGS, FirstCyc );
  output [31:0] Z;
  input [31:0] A;
  input [31:0] B;
  input [31:0] DI;
  output [31:0] DO;
  input [3:0] INST;
  output [3:0] FLAGS;
  input CI, FirstCyc;
  wire   \*Logic0* , \Z_SUM_[32] , N68, n218, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317;
  assign FLAGS[3] = \*Logic0* ;
  assign DO[31] = DI[30];
  assign DO[30] = DI[29];
  assign DO[29] = DI[28];
  assign DO[28] = DI[27];
  assign DO[27] = DI[26];
  assign DO[26] = DI[25];
  assign DO[25] = DI[24];
  assign DO[24] = DI[23];
  assign DO[23] = DI[22];
  assign DO[22] = DI[21];
  assign DO[21] = DI[20];
  assign DO[20] = DI[19];
  assign DO[19] = DI[18];
  assign DO[18] = DI[17];
  assign DO[17] = DI[16];
  assign DO[16] = DI[15];
  assign DO[15] = DI[14];
  assign DO[14] = DI[13];
  assign DO[13] = DI[12];
  assign DO[12] = DI[11];
  assign DO[11] = DI[10];
  assign DO[10] = DI[9];
  assign DO[9] = DI[8];
  assign DO[8] = DI[7];
  assign DO[7] = DI[6];
  assign DO[6] = DI[5];
  assign DO[5] = DI[4];
  assign DO[4] = DI[3];
  assign DO[3] = DI[2];
  assign DO[2] = DI[1];
  assign DO[1] = DI[0];
  assign DO[0] = \Z_SUM_[32] ;
  assign FLAGS[1] = \Z_SUM_[32] ;
  assign N68 = INST[0];

  SEN_INV_AS_5 U408 ( .A(n852), .X(n685) );
  SEN_OR2_1P5 U409 ( .A1(n479), .A2(n957), .X(n480) );
  SEN_ND2_2 U410 ( .A1(n479), .A2(n957), .X(n481) );
  SEN_EN2_S_1 U411 ( .A1(A[15]), .A2(n330), .X(n629) );
  SEN_NR2_T_3 U412 ( .A1(n469), .A2(n350), .X(n957) );
  SEN_INV_2 U413 ( .A(n669), .X(n666) );
  SEN_ND2_2 U414 ( .A1(n663), .A2(n327), .X(n669) );
  SEN_ND2_G_3 U415 ( .A1(n465), .A2(n466), .X(n1285) );
  SEN_EN2_DG_4 U416 ( .A1(n934), .A2(n933), .X(n1295) );
  SEN_ND2B_V1_6 U417 ( .A(n888), .B(n887), .X(n892) );
  SEN_ND2_G_3 U418 ( .A1(n695), .A2(n694), .X(n887) );
  SEN_OAI21_6 U419 ( .A1(n893), .A2(n412), .B(n866), .X(n904) );
  SEN_MUXI2_S_2 U420 ( .D0(n1242), .D1(n1241), .S(INST[3]), .X(FLAGS[2]) );
  SEN_INV_S_3 U421 ( .A(n394), .X(n694) );
  SEN_INV_S_4 U422 ( .A(n390), .X(n585) );
  SEN_NR2_2 U423 ( .A1(n875), .A2(n874), .X(n877) );
  SEN_ND2_T_2 U424 ( .A1(n402), .A2(A[9]), .X(n477) );
  SEN_INV_AS_5 U425 ( .A(n836), .X(n1000) );
  SEN_OAI221_4 U426 ( .A1(n658), .A2(n498), .B1(n657), .B2(n656), .C(n655), 
        .X(n861) );
  SEN_INV_4 U427 ( .A(n658), .X(n657) );
  SEN_INV_4 U428 ( .A(n796), .X(n521) );
  SEN_INV_3 U429 ( .A(n769), .X(n770) );
  SEN_ND2_6 U430 ( .A1(n411), .A2(n1034), .X(n785) );
  SEN_ND2_T_2 U431 ( .A1(n327), .A2(n620), .X(n625) );
  SEN_AN2_4 U432 ( .A1(n861), .A2(n971), .X(n492) );
  SEN_ND2_2 U433 ( .A1(n415), .A2(n416), .X(n417) );
  SEN_AO21B_4 U434 ( .A1(n973), .A2(n972), .B(n971), .X(n490) );
  SEN_ND2_G_4 U435 ( .A1(n496), .A2(n699), .X(n702) );
  SEN_ND2_T_2 U436 ( .A1(n690), .A2(n689), .X(n699) );
  SEN_ND2_G_6 U437 ( .A1(n879), .A2(n872), .X(n874) );
  SEN_INV_2P5 U438 ( .A(n521), .X(n520) );
  SEN_AOI22_T_1P5 U439 ( .A1(n1041), .A2(n1014), .B1(n1013), .B2(n1012), .X(
        n1015) );
  SEN_EO2_3 U440 ( .A1(n1016), .A2(n1015), .X(n1313) );
  SEN_NR2_S_8 U441 ( .A1(n913), .A2(n1268), .X(n428) );
  SEN_ND2_S_4 U442 ( .A1(n487), .A2(n1265), .X(n913) );
  SEN_AOI31_T_4 U443 ( .A1(n776), .A2(n328), .A3(n779), .B(n775), .X(n777) );
  SEN_AN2_6 U444 ( .A1(n1012), .A2(n334), .X(n1001) );
  SEN_ND2_S_3 U445 ( .A1(n328), .A2(n587), .X(n919) );
  SEN_AOAI211_4 U446 ( .A1(n327), .A2(n497), .B(n513), .C(n593), .X(n958) );
  SEN_MUXI2_DG_0P75 U447 ( .D0(n797), .D1(n796), .S(B[20]), .X(n583) );
  SEN_ND2_4 U448 ( .A1(n497), .A2(n594), .X(n592) );
  SEN_INV_6 U449 ( .A(n521), .X(n404) );
  SEN_INV_3 U450 ( .A(n946), .X(n683) );
  SEN_INV_4 U451 ( .A(n945), .X(n464) );
  SEN_ND2_S_1 U452 ( .A1(n1012), .A2(n377), .X(n806) );
  SEN_INV_1 U453 ( .A(n806), .X(n457) );
  SEN_INV_6 U454 ( .A(n874), .X(n691) );
  SEN_INV_S_0P5 U455 ( .A(n735), .X(n343) );
  SEN_ND2_S_4 U456 ( .A1(n453), .A2(n452), .X(n735) );
  SEN_ND2_T_2 U457 ( .A1(n852), .A2(n923), .X(n936) );
  SEN_INV_5 U458 ( .A(n923), .X(n854) );
  SEN_NR2_T_6 U459 ( .A1(n685), .A2(n684), .X(n756) );
  SEN_INV_2 U460 ( .A(n737), .X(n745) );
  SEN_INV_1 U461 ( .A(n854), .X(n450) );
  SEN_EO2_3 U462 ( .A1(n925), .A2(n924), .X(n926) );
  SEN_ND2_S_4 U463 ( .A1(n488), .A2(n459), .X(n462) );
  SEN_AO21B_8 U464 ( .A1(n897), .A2(n898), .B(n870), .X(n488) );
  SEN_NR2_T_8 U465 ( .A1(n552), .A2(n551), .X(n555) );
  SEN_INV_6 U466 ( .A(n607), .X(n832) );
  SEN_INV_1P5 U467 ( .A(n890), .X(n703) );
  SEN_ND2_3 U468 ( .A1(n660), .A2(n661), .X(n662) );
  SEN_ND2_T_6 U469 ( .A1(n756), .A2(n923), .X(n836) );
  SEN_EN2_DG_2 U470 ( .A1(n892), .A2(n891), .X(n1247) );
  SEN_ND2_S_0P5 U471 ( .A1(n890), .A2(n889), .X(n891) );
  SEN_ND2_2 U472 ( .A1(n648), .A2(n527), .X(n661) );
  SEN_EN2_3 U473 ( .A1(A[10]), .A2(n330), .X(n648) );
  SEN_ND2_6 U474 ( .A1(n696), .A2(n697), .X(n706) );
  SEN_INV_S_4 U475 ( .A(n488), .X(n460) );
  SEN_INV_S_2 U476 ( .A(n364), .X(n709) );
  SEN_INV_5 U477 ( .A(n910), .X(n754) );
  SEN_ND2_T_4 U478 ( .A1(n716), .A2(n979), .X(n910) );
  SEN_INV_S_1 U479 ( .A(n856), .X(n857) );
  SEN_INV_12 U480 ( .A(n808), .X(n402) );
  SEN_ND2_0P65 U481 ( .A1(n808), .A2(A[2]), .X(n419) );
  SEN_AO21B_16 U482 ( .A1(n546), .A2(n547), .B(INST[2]), .X(n808) );
  SEN_ND2_T_2 U483 ( .A1(n476), .A2(n477), .X(n651) );
  SEN_INV_5 U484 ( .A(n552), .X(n693) );
  SEN_ND2_6 U485 ( .A1(n544), .A2(INST[1]), .X(n552) );
  SEN_INV_S_0P5 U486 ( .A(n878), .X(n886) );
  SEN_ND2_T_1 U487 ( .A1(n665), .A2(n664), .X(n667) );
  SEN_ND2_T_4 U488 ( .A1(n966), .A2(n670), .X(n967) );
  SEN_ND2_T_2 U489 ( .A1(n669), .A2(n668), .X(n670) );
  SEN_NR2_2 U490 ( .A1(n918), .A2(n958), .X(n921) );
  SEN_ND2_T_2 U491 ( .A1(n751), .A2(n899), .X(n978) );
  SEN_ND2_2 U492 ( .A1(n379), .A2(n380), .X(n498) );
  SEN_ND2_2 U493 ( .A1(n511), .A2(B[9]), .X(n380) );
  SEN_ND2_2 U494 ( .A1(n652), .A2(n498), .X(n656) );
  SEN_ND2_G_0P65 U495 ( .A1(B[8]), .A2(n483), .X(n652) );
  SEN_ND2B_V1DG_4 U496 ( .A(n763), .B(n761), .X(n1034) );
  SEN_ND2_S_2 U497 ( .A1(n574), .A2(n573), .X(n761) );
  SEN_EN2_S_1 U498 ( .A1(A[23]), .A2(n329), .X(n559) );
  SEN_EN2_S_2 U499 ( .A1(A[8]), .A2(n329), .X(n711) );
  SEN_EN2_3 U500 ( .A1(A[1]), .A2(n329), .X(n698) );
  SEN_EN2_S_2 U501 ( .A1(A[13]), .A2(n329), .X(n617) );
  SEN_ND2_T_1 U502 ( .A1(n904), .A2(n872), .X(n885) );
  SEN_ND2_T_6 U503 ( .A1(n634), .A2(n939), .X(n954) );
  SEN_INV_3 U504 ( .A(n997), .X(n998) );
  SEN_ND2_4 U505 ( .A1(n644), .A2(n828), .X(n997) );
  SEN_INV_S_3 U506 ( .A(n720), .X(n721) );
  SEN_ND2_S_3 U507 ( .A1(n719), .A2(n718), .X(n720) );
  SEN_ND2_2 U508 ( .A1(n736), .A2(n368), .X(n731) );
  SEN_ND2_G_3 U509 ( .A1(n327), .A2(n548), .X(n767) );
  SEN_ND2B_4 U510 ( .A(n767), .B(n765), .X(n839) );
  SEN_ND2_T_4 U511 ( .A1(n407), .A2(n979), .X(n972) );
  SEN_ND2_S_0P65 U512 ( .A1(n980), .A2(n979), .X(n985) );
  SEN_ND2_0P5 U513 ( .A1(n971), .A2(n979), .X(n856) );
  SEN_ND2_4 U514 ( .A1(n715), .A2(n714), .X(n979) );
  SEN_OAI21_G_6 U515 ( .A1(INST[2]), .A2(n553), .B(n351), .X(n554) );
  SEN_INV_10 U516 ( .A(INST[1]), .X(n351) );
  SEN_EN2_1 U517 ( .A1(A[5]), .A2(n808), .X(n724) );
  SEN_ND2_S_3 U518 ( .A1(B[13]), .A2(n483), .X(n682) );
  SEN_ND3_T_4 U519 ( .A1(n642), .A2(n326), .A3(n940), .X(n643) );
  SEN_NR3_T_8 U520 ( .A1(n1274), .A2(n912), .A3(n429), .X(n930) );
  SEN_INV_6 U521 ( .A(N68), .X(n547) );
  SEN_INV_S_1 U522 ( .A(n808), .X(n403) );
  SEN_ND2_S_1P5 U523 ( .A1(B[10]), .A2(n483), .X(n665) );
  SEN_MUXI2_S_2 U524 ( .D0(n522), .D1(n796), .S(B[11]), .X(n664) );
  SEN_INV_10 U525 ( .A(A[31]), .X(n470) );
  SEN_ND2_T_3 U526 ( .A1(n641), .A2(n640), .X(n642) );
  SEN_ND2_T_4 U527 ( .A1(n335), .A2(n848), .X(n828) );
  SEN_ND2_T_2 U528 ( .A1(n328), .A2(n617), .X(n678) );
  SEN_MUXI2_D_1 U529 ( .D0(n522), .D1(n796), .S(B[7]), .X(n718) );
  SEN_INV_S_0P5 U530 ( .A(n977), .X(n964) );
  SEN_NR2_S_0P65 U531 ( .A1(n433), .A2(n962), .X(n963) );
  SEN_ND2_3 U532 ( .A1(n650), .A2(n649), .X(n659) );
  SEN_INV_S_2 U533 ( .A(n417), .X(n649) );
  SEN_INV_1P5 U534 ( .A(n659), .X(n660) );
  SEN_AN2_4 U535 ( .A1(n863), .A2(n870), .X(n491) );
  SEN_ND2_T_3 U536 ( .A1(n517), .A2(n731), .X(n870) );
  SEN_ND2_0P5 U537 ( .A1(n434), .A2(n952), .X(n437) );
  SEN_AO21B_4 U538 ( .A1(n953), .A2(n952), .B(n951), .X(n485) );
  SEN_OAOI211_3 U539 ( .A1(n986), .A2(n985), .B(n984), .C(n983), .X(n987) );
  SEN_EO2_2 U540 ( .A1(n988), .A2(n987), .X(n1273) );
  SEN_BUF_2 U541 ( .A(n961), .X(n341) );
  SEN_INV_6 U542 ( .A(n931), .X(n1041) );
  SEN_NR2_S_1 U543 ( .A1(n932), .A2(n931), .X(n933) );
  SEN_ND2_T_4 U544 ( .A1(n836), .A2(n997), .X(n931) );
  SEN_EN2_DG_4 U545 ( .A1(n895), .A2(n894), .X(n1250) );
  SEN_ND2_T_16 U546 ( .A1(n472), .A2(n473), .X(n546) );
  SEN_ND2_T_16 U547 ( .A1(n471), .A2(n470), .X(n473) );
  SEN_ND2_16 U548 ( .A1(A[31]), .A2(n338), .X(n472) );
  SEN_ND2_T_4 U549 ( .A1(n639), .A2(n328), .X(n637) );
  SEN_ND2_S_4 U550 ( .A1(n643), .A2(n683), .X(n848) );
  SEN_INV_4 U551 ( .A(n915), .X(n956) );
  SEN_ND2_2 U552 ( .A1(n830), .A2(n852), .X(n914) );
  SEN_EN2_S_1 U553 ( .A1(A[11]), .A2(n329), .X(n663) );
  SEN_ND3_T_1 U554 ( .A1(n341), .A2(n971), .A3(n966), .X(n977) );
  SEN_AN4B_4 U555 ( .B1(n982), .B2(n966), .B3(n341), .A(n856), .X(n755) );
  SEN_ND2_6 U556 ( .A1(n667), .A2(n666), .X(n966) );
  SEN_AO21_1 U557 ( .A1(n905), .A2(n904), .B(n903), .X(n401) );
  SEN_INV_S_4 U558 ( .A(n904), .X(n875) );
  SEN_OAI21B_2 U559 ( .A1(n1022), .A2(n1024), .B(n837), .X(n821) );
  SEN_INV_S_2 U560 ( .A(n839), .X(n837) );
  SEN_INV_0P5 U561 ( .A(n981), .X(n984) );
  SEN_ND2_G_3 U562 ( .A1(n604), .A2(n591), .X(n916) );
  SEN_ND2_2 U563 ( .A1(n589), .A2(n588), .X(n604) );
  SEN_INV_1P5 U564 ( .A(n605), .X(n591) );
  SEN_ND2_S_4 U565 ( .A1(n1026), .A2(n1023), .X(n932) );
  SEN_AN3B_2 U566 ( .B1(n908), .B2(n907), .A(n906), .X(n909) );
  SEN_ND2_2 U567 ( .A1(n584), .A2(n583), .X(n595) );
  SEN_INV_S_2 U568 ( .A(n595), .X(n596) );
  SEN_NR2_T_4 U569 ( .A1(n458), .A2(n805), .X(n950) );
  SEN_NR3_T_4 U570 ( .A1(n456), .A2(n457), .A3(n325), .X(n458) );
  SEN_ND2B_6 U571 ( .A(n702), .B(n328), .X(n872) );
  SEN_MUXI2_S_0P5 U572 ( .D0(n1317), .D1(n1316), .S(INST[3]), .X(Z[31]) );
  SEN_NR3_T_6 U573 ( .A1(n1277), .A2(n989), .A3(n1288), .X(n1006) );
  SEN_ND2_G_3 U574 ( .A1(n444), .A2(n445), .X(n1277) );
  SEN_EN2_S_4 U575 ( .A1(n494), .A2(n950), .X(n1317) );
  SEN_MUXI2_S_3 U576 ( .D0(n522), .D1(n520), .S(B[12]), .X(n646) );
  SEN_INV_2 U577 ( .A(n970), .X(n340) );
  SEN_NR2B_V1_2 U578 ( .A(n937), .B(n936), .X(n943) );
  SEN_NR3_T_2 U579 ( .A1(n936), .A2(n845), .A3(n927), .X(n846) );
  SEN_NR2_T_1P5 U580 ( .A1(n936), .A2(n927), .X(n928) );
  SEN_ND2_S_4 U581 ( .A1(n1295), .A2(n1285), .X(n947) );
  SEN_AOI31_3 U582 ( .A1(n858), .A2(n859), .A3(n514), .B(n959), .X(n860) );
  SEN_INV_4 U583 ( .A(n428), .X(n429) );
  SEN_EN2_1 U584 ( .A1(A[17]), .A2(n329), .X(n609) );
  SEN_ND2_2 U585 ( .A1(n327), .A2(n609), .X(n615) );
  SEN_ND2_4 U586 ( .A1(n486), .A2(n966), .X(n339) );
  SEN_NR3_G_4 U587 ( .A1(n1000), .A2(n999), .A3(n998), .X(n1003) );
  SEN_ND2_T_4 U588 ( .A1(n342), .A2(n899), .X(n433) );
  SEN_INV_8 U589 ( .A(n402), .X(n524) );
  SEN_OR4B_4 U590 ( .B1(n837), .B2(n990), .B3(n600), .A(n1017), .X(n999) );
  SEN_EO2_S_3 U591 ( .A1(n1043), .A2(n1042), .X(n1297) );
  SEN_ND2_T_4 U592 ( .A1(n1306), .A2(n1297), .X(n1044) );
  SEN_AOI211_3 U593 ( .A1(n879), .A2(n336), .B1(n877), .B2(n876), .X(n882) );
  SEN_ND2_T_2 U594 ( .A1(n359), .A2(n360), .X(n1255) );
  SEN_ND2_T_1P5 U595 ( .A1(n402), .A2(A[14]), .X(n423) );
  SEN_INV_S_6 U596 ( .A(n681), .X(n639) );
  SEN_ND2_3 U597 ( .A1(n996), .A2(n382), .X(n383) );
  SEN_INV_3 U598 ( .A(n699), .X(n700) );
  SEN_INV_S_6 U599 ( .A(n926), .X(n1291) );
  SEN_NR2_S_4 U600 ( .A1(n882), .A2(n881), .X(n883) );
  SEN_NR2_T_3 U601 ( .A1(n956), .A2(n917), .X(n918) );
  SEN_OAI21B_6 U602 ( .A1(n859), .A2(n959), .B(n967), .X(n671) );
  SEN_INV_S_6 U603 ( .A(n974), .X(n859) );
  SEN_ND2B_V1DG_4 U604 ( .A(n478), .B(n654), .X(n658) );
  SEN_INV_4 U605 ( .A(n651), .X(n654) );
  SEN_NR2_G_2 U606 ( .A1(n401), .A2(n902), .X(n906) );
  SEN_ND2_S_6 U607 ( .A1(n339), .A2(n340), .X(n981) );
  SEN_ND2B_V1_2 U608 ( .A(n975), .B(n852), .X(n855) );
  SEN_INV_1 U609 ( .A(n952), .X(n435) );
  SEN_OAI21_S_8 U610 ( .A1(n855), .A2(n854), .B(n853), .X(n952) );
  SEN_ND2_S_4 U611 ( .A1(n386), .A2(n519), .X(n912) );
  SEN_ND2_T_2 U612 ( .A1(n746), .A2(n741), .X(n742) );
  SEN_MUX2_DG_1 U613 ( .D0(n1286), .D1(n1287), .S(INST[3]), .X(Z[18]) );
  SEN_EO2_2 U614 ( .A1(n850), .A2(n849), .X(n1286) );
  SEN_ND2_T_6 U615 ( .A1(n981), .A2(n982), .X(n852) );
  SEN_ND2_T_2 U616 ( .A1(n327), .A2(n577), .X(n580) );
  SEN_ND2_S_0P8 U617 ( .A1(B[4]), .A2(n483), .X(n726) );
  SEN_BUF_20 U618 ( .A(n812), .X(n483) );
  SEN_INV_3 U619 ( .A(n713), .X(n714) );
  SEN_ND2_2 U620 ( .A1(n712), .A2(n713), .X(n716) );
  SEN_ND2_3 U621 ( .A1(n328), .A2(n711), .X(n713) );
  SEN_AOAI211_G_3 U622 ( .A1(n328), .A2(n779), .B(n778), .C(n777), .X(n934) );
  SEN_EN2_S_2 U623 ( .A1(A[4]), .A2(n329), .X(n686) );
  SEN_OA2BB2_2 U624 ( .A1(n1034), .A2(n1033), .B1(n1032), .B2(n1031), .X(n1035) );
  SEN_ND2_3 U625 ( .A1(n422), .A2(n423), .X(n681) );
  SEN_OR3B_2 U626 ( .B1(n651), .B2(n478), .A(n656), .X(n971) );
  SEN_ND2_4 U627 ( .A1(n961), .A2(n662), .X(n974) );
  SEN_ND3_T_4 U628 ( .A1(n1048), .A2(n1317), .A3(n1047), .X(n1242) );
  SEN_ND2_S_6 U629 ( .A1(n1313), .A2(n1300), .X(n1045) );
  SEN_MUXI2_S_0P5 U630 ( .D0(n1313), .D1(n1312), .S(INST[3]), .X(Z[29]) );
  SEN_NR3_T_4 U631 ( .A1(n949), .A2(n948), .A3(n947), .X(n1048) );
  SEN_NR2_T_2 U632 ( .A1(n346), .A2(n347), .X(\Z_SUM_[32] ) );
  SEN_NR2_T_1P5 U633 ( .A1(n458), .A2(n348), .X(n346) );
  SEN_EO2_2 U634 ( .A1(n876), .A2(n873), .X(n1253) );
  SEN_ND2B_V1_2 U635 ( .A(n661), .B(n659), .X(n961) );
  SEN_INV_2 U636 ( .A(n914), .X(n922) );
  SEN_OAI211_3 U637 ( .A1(n736), .A2(n344), .B1(n752), .B2(n734), .X(n863) );
  SEN_INV_S_2 U638 ( .A(n343), .X(n344) );
  SEN_ND3_S_4 U639 ( .A1(n1271), .A2(n489), .A3(n1273), .X(n989) );
  SEN_EO2_G_2 U640 ( .A1(n974), .A2(n490), .X(n489) );
  SEN_AO21B_16 U641 ( .A1(n546), .A2(n547), .B(INST[2]), .X(n330) );
  SEN_MUXI2_D_1 U642 ( .D0(n1295), .D1(n1294), .S(INST[3]), .X(Z[22]) );
  SEN_ND2_6 U643 ( .A1(n698), .A2(n328), .X(n704) );
  SEN_EO2_1 U644 ( .A1(n886), .A2(n885), .X(n1251) );
  SEN_INV_2P5 U645 ( .A(n478), .X(n327) );
  SEN_EN2_0P5 U646 ( .A1(A[29]), .A2(n523), .X(n601) );
  SEN_ND2B_V1_3 U647 ( .A(n678), .B(n676), .X(n853) );
  SEN_INV_S_3 U648 ( .A(n835), .X(n608) );
  SEN_EN2_S_3 U649 ( .A1(A[21]), .A2(n524), .X(n577) );
  SEN_ND2_T_2 U650 ( .A1(n576), .A2(n575), .X(n579) );
  SEN_MUXI2_DG_2 U651 ( .D0(n522), .D1(n520), .S(B[21]), .X(n575) );
  SEN_ND2B_V1_3 U652 ( .A(n788), .B(n786), .X(n991) );
  SEN_INV_3 U653 ( .A(n932), .X(n1017) );
  SEN_ND2_S_6 U654 ( .A1(n633), .A2(n632), .X(n939) );
  SEN_INV_S_3 U655 ( .A(n631), .X(n632) );
  SEN_ND2_T_2 U656 ( .A1(n606), .A2(n916), .X(n850) );
  SEN_INV_3 U657 ( .A(n773), .X(n779) );
  SEN_INV_0P65 U658 ( .A(\Z_SUM_[32] ), .X(n439) );
  SEN_ND2B_V1DG_4 U659 ( .A(n478), .B(n518), .X(n746) );
  SEN_ND2_2 U660 ( .A1(n403), .A2(A[6]), .X(n453) );
  SEN_ND2_2 U661 ( .A1(n329), .A2(n451), .X(n452) );
  SEN_ND2_G_1 U662 ( .A1(n796), .A2(B[10]), .X(n416) );
  SEN_ND2_2 U663 ( .A1(n797), .A2(n414), .X(n415) );
  SEN_ND2_S_3 U664 ( .A1(n388), .A2(n389), .X(n390) );
  SEN_ND2_G_1 U665 ( .A1(n431), .A2(n432), .X(n717) );
  SEN_ND2_T_1 U666 ( .A1(n430), .A2(n402), .X(n432) );
  SEN_ND2_2 U667 ( .A1(n612), .A2(n613), .X(n847) );
  SEN_ND2_2 U668 ( .A1(n774), .A2(n562), .X(n778) );
  SEN_ND2_2 U669 ( .A1(n528), .A2(n559), .X(n771) );
  SEN_AOAI211_6 U670 ( .A1(n790), .A2(n992), .B(n827), .C(n991), .X(n993) );
  SEN_NR2_1 U671 ( .A1(n1244), .A2(n1245), .X(n1091) );
  SEN_ND2_S_3 U672 ( .A1(n392), .A2(n393), .X(n394) );
  SEN_ND2B_3 U673 ( .A(n706), .B(n704), .X(n890) );
  SEN_INV_S_2 U674 ( .A(n704), .X(n705) );
  SEN_ND2_3 U675 ( .A1(n579), .A2(n578), .X(n1026) );
  SEN_ND2_G_1 U676 ( .A1(n1013), .A2(n760), .X(n996) );
  SEN_INV_S_0P5 U677 ( .A(n992), .X(n1007) );
  SEN_ND2B_S_2 U678 ( .A(n990), .B(n1017), .X(n1009) );
  SEN_INV_S_1 U679 ( .A(n791), .X(n792) );
  SEN_ND2B_1 U680 ( .A(n793), .B(n791), .X(n1002) );
  SEN_ND3_S_4 U681 ( .A1(n1293), .A2(n1309), .A3(n1303), .X(n949) );
  SEN_ND2_G_1 U682 ( .A1(n440), .A2(n441), .X(FLAGS[0]) );
  SEN_ND2_G_1 U683 ( .A1(n438), .A2(n439), .X(n441) );
  SEN_INV_10 U684 ( .A(n545), .X(n471) );
  SEN_ND2_G_1 U685 ( .A1(n330), .A2(n421), .X(n422) );
  SEN_ND2_G_1 U686 ( .A1(n797), .A2(n446), .X(n447) );
  SEN_INV_S_1 U687 ( .A(n652), .X(n653) );
  SEN_INV_2 U688 ( .A(n402), .X(n523) );
  SEN_INV_4 U689 ( .A(INST[3]), .X(n544) );
  SEN_ND2_2 U690 ( .A1(n796), .A2(B[0]), .X(n393) );
  SEN_ND2_G_1 U691 ( .A1(n797), .A2(n397), .X(n398) );
  SEN_INV_S_1 U692 ( .A(B[1]), .X(n397) );
  SEN_ND2_2 U693 ( .A1(n420), .A2(n419), .X(n496) );
  SEN_INV_S_1 U694 ( .A(A[2]), .X(n418) );
  SEN_ND2_T_1 U695 ( .A1(B[1]), .A2(n483), .X(n690) );
  SEN_INV_3 U696 ( .A(n895), .X(n866) );
  SEN_ND2_T_1 U697 ( .A1(n619), .A2(n618), .X(n676) );
  SEN_MUXI2_D_1 U698 ( .D0(n522), .D1(n796), .S(B[13]), .X(n618) );
  SEN_ND2_2 U699 ( .A1(n328), .A2(n629), .X(n631) );
  SEN_AN2_3 U700 ( .A1(n951), .A2(n853), .X(n493) );
  SEN_MUXI2_S_1 U701 ( .D0(n522), .D1(n404), .S(B[18]), .X(n588) );
  SEN_ND2_G_1 U702 ( .A1(n680), .A2(n951), .X(n640) );
  SEN_ND2_G_1 U703 ( .A1(B[21]), .A2(n525), .X(n774) );
  SEN_INV_2 U704 ( .A(n1039), .X(n838) );
  SEN_ND2_2 U705 ( .A1(n1025), .A2(n934), .X(n1039) );
  SEN_INV_1 U706 ( .A(n1030), .X(n1033) );
  SEN_ND2_T_1 U707 ( .A1(n565), .A2(n564), .X(n786) );
  SEN_ND2_G_1 U708 ( .A1(n327), .A2(n563), .X(n788) );
  SEN_MUXI2_D_1 U709 ( .D0(n522), .D1(n404), .S(B[25]), .X(n573) );
  SEN_INV_S_2 U710 ( .A(n961), .X(n959) );
  SEN_ND2_G_4 U711 ( .A1(n831), .A2(n598), .X(n925) );
  SEN_ND2_G_1 U712 ( .A1(n597), .A2(n596), .X(n598) );
  SEN_ND2_G_4 U713 ( .A1(n581), .A2(n1026), .X(n835) );
  SEN_ND2_S_6 U714 ( .A1(n1024), .A2(n772), .X(n1043) );
  SEN_ND2_2 U715 ( .A1(n771), .A2(n770), .X(n772) );
  SEN_ND2_2 U716 ( .A1(n992), .A2(n783), .X(n1037) );
  SEN_INV_S_1 U717 ( .A(n780), .X(n781) );
  SEN_MUXI2_S_1 U718 ( .D0(n406), .D1(n1088), .S(A[1]), .X(n1089) );
  SEN_EO2_2 U719 ( .A1(n754), .A2(n909), .X(n519) );
  SEN_INV_S_4 U720 ( .A(n862), .X(n1265) );
  SEN_ND2_S_2 U721 ( .A1(n436), .A2(n437), .X(n1274) );
  SEN_ND2_G_1 U722 ( .A1(n953), .A2(n435), .X(n436) );
  SEN_ND2_G_1 U723 ( .A1(n954), .A2(n485), .X(n444) );
  SEN_AN3B_1 U724 ( .B1(n848), .B2(n335), .A(n846), .X(n849) );
  SEN_MUX2_DG_1 U725 ( .D0(n323), .D1(n1269), .S(INST[3]), .X(Z[11]) );
  SEN_MUXI2_S_1 U726 ( .D0(n1282), .D1(n1281), .S(INST[3]), .X(Z[16]) );
  SEN_MUXI2_S_1 U727 ( .D0(n1300), .D1(n1299), .S(INST[3]), .X(Z[24]) );
  SEN_ND2_3 U728 ( .A1(n371), .A2(n372), .X(n1306) );
  SEN_ND2_S_3 U729 ( .A1(n911), .A2(n484), .X(n385) );
  SEN_ND2_G_4 U730 ( .A1(n461), .A2(n462), .X(n487) );
  SEN_MUX2_DG_1 U731 ( .D0(n1255), .D1(n1256), .S(INST[3]), .X(Z[5]) );
  SEN_ND2_T_1P5 U732 ( .A1(n753), .A2(n752), .X(n426) );
  SEN_ND2B_V1_1 U733 ( .A(n491), .B(n899), .X(n903) );
  SEN_NR2_S_0P65 U734 ( .A1(n893), .A2(n412), .X(n894) );
  SEN_INV_2 U735 ( .A(n517), .X(n732) );
  SEN_ND2_T_2 U736 ( .A1(n369), .A2(n370), .X(n372) );
  SEN_INV_2 U737 ( .A(n636), .X(n322) );
  SEN_INV_3 U738 ( .A(n635), .X(n636) );
  SEN_ND2B_2 U739 ( .A(n638), .B(n682), .X(n635) );
  SEN_ND3_S_8 U740 ( .A1(n408), .A2(n409), .A3(n410), .X(n411) );
  SEN_INV_S_6 U741 ( .A(n820), .X(n409) );
  SEN_INV_2 U742 ( .A(n869), .X(n424) );
  SEN_ND2_G_3 U743 ( .A1(n796), .A2(B[1]), .X(n399) );
  SEN_ND2_G_4 U744 ( .A1(n880), .A2(n750), .X(n876) );
  SEN_EO2_G_4 U745 ( .A1(n970), .A2(n969), .X(n1271) );
  SEN_INV_2 U746 ( .A(n1037), .X(n784) );
  SEN_ND2_G_1 U747 ( .A1(n982), .A2(n675), .X(n970) );
  SEN_ND2_G_1 U748 ( .A1(n674), .A2(n673), .X(n675) );
  SEN_ND2_3 U749 ( .A1(n767), .A2(n766), .X(n768) );
  SEN_ND2_T_4 U750 ( .A1(n561), .A2(n560), .X(n769) );
  SEN_MUXI2_DG_5 U751 ( .D0(n797), .D1(n404), .S(B[23]), .X(n560) );
  SEN_INV_S_1 U752 ( .A(n1274), .X(n1276) );
  SEN_AN3B_4 U753 ( .B1(n829), .B2(n608), .A(n832), .X(n644) );
  SEN_AOAI211_6 U754 ( .A1(n919), .A2(n958), .B(n925), .C(n831), .X(n607) );
  SEN_ND2_3 U755 ( .A1(n607), .A2(n468), .X(n1023) );
  SEN_INV_3 U756 ( .A(n867), .X(n905) );
  SEN_ND2_T_6 U757 ( .A1(n691), .A2(n880), .X(n867) );
  SEN_INV_2 U758 ( .A(n765), .X(n766) );
  SEN_INV_8 U759 ( .A(n871), .X(n901) );
  SEN_OAI21_S_2 U760 ( .A1(n838), .A2(n1043), .B(n1024), .X(n1019) );
  SEN_ND2B_3 U761 ( .A(n625), .B(n623), .X(n940) );
  SEN_ND2_S_4 U762 ( .A1(n1034), .A2(n764), .X(n844) );
  SEN_ND2_2 U763 ( .A1(n763), .A2(n762), .X(n764) );
  SEN_INV_S_16 U764 ( .A(n738), .X(n796) );
  SEN_BUF_1 U765 ( .A(n1268), .X(n323) );
  SEN_AN4B_2 U766 ( .B1(n992), .B2(n1011), .B3(n991), .A(n1009), .X(n994) );
  SEN_INV_S_6 U767 ( .A(n865), .X(n893) );
  SEN_OAI21_4 U768 ( .A1(n702), .A2(n478), .B(n701), .X(n895) );
  SEN_EN2_S_3 U769 ( .A1(A[18]), .A2(n523), .X(n590) );
  SEN_BUF_1 U770 ( .A(n1315), .X(n324) );
  SEN_ND2_T_4 U771 ( .A1(n480), .A2(n481), .X(n1288) );
  SEN_MUXI2_DG_1 U772 ( .D0(n797), .D1(n796), .S(B[4]), .X(n687) );
  SEN_OAI21_G_12 U773 ( .A1(n550), .A2(INST[1]), .B(N68), .X(n810) );
  SEN_INV_S_1 U774 ( .A(n478), .X(n527) );
  SEN_INV_3 U775 ( .A(n478), .X(n328) );
  SEN_INV_4 U776 ( .A(n810), .X(n797) );
  SEN_INV_S_1 U777 ( .A(n900), .X(n357) );
  SEN_AO21_1 U778 ( .A1(n1016), .A2(n1002), .B(n1005), .X(n325) );
  SEN_INV_S_1 U779 ( .A(n218), .X(n540) );
  SEN_ND2_G_3 U780 ( .A1(n940), .A2(n626), .X(n935) );
  SEN_ND2B_V1_4 U781 ( .A(n771), .B(n769), .X(n1024) );
  SEN_OR2_1 U782 ( .A1(n935), .A2(n939), .X(n326) );
  SEN_ND2_2 U783 ( .A1(n692), .A2(n327), .X(n888) );
  SEN_INV_2 U784 ( .A(n810), .X(n522) );
  SEN_INV_S_1 U785 ( .A(n368), .X(n733) );
  SEN_AO21B_8 U786 ( .A1(n546), .A2(n547), .B(INST[2]), .X(n329) );
  SEN_INV_1P25 U787 ( .A(n747), .X(n748) );
  SEN_ND3_2 U788 ( .A1(n831), .A2(n919), .A3(n916), .X(n599) );
  SEN_INV_3 U789 ( .A(n844), .X(n408) );
  SEN_ND2_2 U790 ( .A1(n357), .A2(n358), .X(n360) );
  SEN_ND2_G_1 U791 ( .A1(n678), .A2(n677), .X(n679) );
  SEN_ND2B_3 U792 ( .A(n592), .B(n327), .X(n593) );
  SEN_EN2_1 U793 ( .A1(n898), .A2(n897), .X(n484) );
  SEN_ND2_T_1 U794 ( .A1(n330), .A2(n475), .X(n476) );
  SEN_EN2_1 U795 ( .A1(A[16]), .A2(n330), .X(n620) );
  SEN_EN2_S_1 U796 ( .A1(n345), .A2(n402), .X(n582) );
  SEN_ND2B_3 U797 ( .A(n729), .B(n727), .X(n868) );
  SEN_INV_S_1 U798 ( .A(n838), .X(n331) );
  SEN_INV_S_0P5 U799 ( .A(n639), .X(n332) );
  SEN_INV_S_6 U800 ( .A(n976), .X(n962) );
  SEN_ND2_T_1 U801 ( .A1(n796), .A2(B[8]), .X(n363) );
  SEN_ND2_S_0P8 U802 ( .A1(B[6]), .A2(n483), .X(n719) );
  SEN_ND2_2 U803 ( .A1(n630), .A2(n631), .X(n634) );
  SEN_EO2_3 U804 ( .A1(n844), .A2(n843), .X(n1303) );
  SEN_ND2_0P5 U805 ( .A1(B[14]), .A2(n483), .X(n628) );
  SEN_ND2B_V1_6 U806 ( .A(n996), .B(n993), .X(n1012) );
  SEN_ND2_3 U807 ( .A1(n828), .A2(n829), .X(n915) );
  SEN_BUF_1 U808 ( .A(n887), .X(n333) );
  SEN_ND2_G_1 U809 ( .A1(n1002), .A2(n794), .X(n1016) );
  SEN_ND2_G_1 U810 ( .A1(n793), .A2(n792), .X(n794) );
  SEN_ND2_G_1 U811 ( .A1(n529), .A2(n601), .X(n793) );
  SEN_INV_S_0P5 U812 ( .A(n1024), .X(n1018) );
  SEN_ND2B_S_4 U813 ( .A(n749), .B(n747), .X(n880) );
  SEN_ND2_2 U814 ( .A1(n647), .A2(n646), .X(n672) );
  SEN_ND2_0P5 U815 ( .A1(n586), .A2(n585), .X(n513) );
  SEN_INV_S_4 U816 ( .A(n892), .X(n864) );
  SEN_INV_0P8 U817 ( .A(n919), .X(n920) );
  SEN_ND2_3 U818 ( .A1(n868), .A2(n730), .X(n884) );
  SEN_INV_0P8 U819 ( .A(n1023), .X(n1029) );
  SEN_INV_S_6 U820 ( .A(n884), .X(n900) );
  SEN_AN2_6 U821 ( .A1(n706), .A2(n705), .X(n412) );
  SEN_ND2_T_4 U822 ( .A1(n383), .A2(n384), .X(n1311) );
  SEN_ND2_2 U823 ( .A1(n868), .A2(n870), .X(n753) );
  SEN_ND2_T_8 U824 ( .A1(n482), .A2(n755), .X(n923) );
  SEN_AN2_S_1 U825 ( .A1(n1002), .A2(n1013), .X(n334) );
  SEN_ND2B_S_2 U826 ( .A(n759), .B(n757), .X(n1013) );
  SEN_ND2_2 U827 ( .A1(n900), .A2(n883), .X(n359) );
  SEN_AO21B_4 U828 ( .A1(n496), .A2(n528), .B(n700), .X(n701) );
  SEN_ND2_T_2 U829 ( .A1(n625), .A2(n624), .X(n626) );
  SEN_INV_S_4 U830 ( .A(n623), .X(n624) );
  SEN_ND2_2 U831 ( .A1(n599), .A2(n608), .X(n467) );
  SEN_ND2B_3 U832 ( .A(n674), .B(n672), .X(n982) );
  SEN_ND2_2 U833 ( .A1(n724), .A2(n328), .X(n729) );
  SEN_ND2_0P8 U834 ( .A1(B[9]), .A2(n483), .X(n650) );
  SEN_ND2B_1 U835 ( .A(n604), .B(n605), .X(n606) );
  SEN_NR2_4 U836 ( .A1(n978), .A2(n962), .X(n395) );
  SEN_ND2_S_2 U837 ( .A1(n946), .A2(n945), .X(n465) );
  SEN_ND2_G_4 U838 ( .A1(n864), .A2(n890), .X(n865) );
  SEN_EN2_0P5 U839 ( .A1(n888), .A2(n333), .X(n1243) );
  SEN_ND2_T_8 U840 ( .A1(n1050), .A2(n693), .X(n549) );
  SEN_INV_S_4 U841 ( .A(n400), .X(n696) );
  SEN_NR2_T_16 U842 ( .A1(n351), .A2(B[31]), .X(n338) );
  SEN_INV_3 U843 ( .A(n551), .X(n1050) );
  SEN_INV_S_16 U844 ( .A(n549), .X(n812) );
  SEN_ND2_S_0P65 U845 ( .A1(B[3]), .A2(n483), .X(n688) );
  SEN_BUF_1 U846 ( .A(n847), .X(n335) );
  SEN_ND2_G_1 U847 ( .A1(n529), .A2(n795), .X(n802) );
  SEN_ND2_S_4 U848 ( .A1(n398), .A2(n399), .X(n400) );
  SEN_INV_2 U849 ( .A(n467), .X(n468) );
  SEN_BUF_S_2 U850 ( .A(n878), .X(n336) );
  SEN_ND2B_6 U851 ( .A(n337), .B(n322), .X(n951) );
  SEN_ND2_T_2 U852 ( .A1(n639), .A2(n327), .X(n337) );
  SEN_OR3B_8 U853 ( .B1(n835), .B2(n832), .A(n830), .X(n684) );
  SEN_ND2_4 U854 ( .A1(n424), .A2(n900), .X(n425) );
  SEN_ND3_T_6 U855 ( .A1(n905), .A2(n708), .A3(n707), .X(n976) );
  SEN_ND2B_2 U856 ( .A(n579), .B(n580), .X(n581) );
  SEN_MUXI2_DG_3 U857 ( .D0(n797), .D1(n796), .S(B[2]), .X(n689) );
  SEN_ND2_T_1P5 U858 ( .A1(n749), .A2(n748), .X(n750) );
  SEN_ND2_T_1 U859 ( .A1(n796), .A2(B[16]), .X(n448) );
  SEN_INV_S_3 U860 ( .A(n449), .X(n621) );
  SEN_INV_S_2 U861 ( .A(n935), .X(n942) );
  SEN_ND2_T_4 U862 ( .A1(n425), .A2(n868), .X(n897) );
  SEN_ND2_T_2 U863 ( .A1(n726), .A2(n725), .X(n727) );
  SEN_MUXI2_DG_2 U864 ( .D0(n522), .D1(n796), .S(B[5]), .X(n725) );
  SEN_INV_2 U865 ( .A(n727), .X(n728) );
  SEN_ND2_G_1 U866 ( .A1(n939), .A2(n938), .X(n941) );
  SEN_NR3_T_3 U867 ( .A1(n493), .A2(n935), .A3(n954), .X(n641) );
  SEN_ND2_T_1 U868 ( .A1(n402), .A2(n418), .X(n420) );
  SEN_OR3B_2 U869 ( .B1(n892), .B2(n703), .A(n866), .X(n708) );
  SEN_INV_S_4 U870 ( .A(n838), .X(n410) );
  SEN_ND2_S_0P5 U871 ( .A1(n950), .A2(\Z_SUM_[32] ), .X(n440) );
  SEN_ND2_2 U872 ( .A1(n442), .A2(n443), .X(n445) );
  SEN_NR3_T_12 U873 ( .A1(n927), .A2(n845), .A3(n850), .X(n830) );
  SEN_OAOI211_3 U874 ( .A1(n968), .A2(n352), .B(n966), .C(n965), .X(n969) );
  SEN_ND2_S_4 U875 ( .A1(n586), .A2(n585), .X(n594) );
  SEN_ND2B_V1_3 U876 ( .A(n597), .B(n595), .X(n831) );
  SEN_INV_S_2 U877 ( .A(n807), .X(n456) );
  SEN_MUXI2_S_0P5 U878 ( .D0(n1271), .D1(n1270), .S(INST[3]), .X(Z[12]) );
  SEN_INV_S_1P5 U879 ( .A(n995), .X(n382) );
  SEN_ND2_S_2 U880 ( .A1(n995), .A2(n381), .X(n384) );
  SEN_ND2_6 U881 ( .A1(n851), .A2(n951), .X(n937) );
  SEN_INV_1P5 U882 ( .A(n633), .X(n630) );
  SEN_ND2_3 U883 ( .A1(n327), .A2(n590), .X(n605) );
  SEN_AN3_8 U884 ( .A1(INST[2]), .A2(INST[1]), .A3(N68), .X(n478) );
  SEN_AN2_24 U885 ( .A1(N68), .A2(INST[1]), .X(n556) );
  SEN_NR2_T_2 U886 ( .A1(n833), .A2(n515), .X(n834) );
  SEN_AOAI211_0P75 U887 ( .A1(n409), .A2(n331), .B(n821), .C(n1032), .X(n823)
         );
  SEN_ND2_S_0P5 U888 ( .A1(n1024), .A2(n1025), .X(n990) );
  SEN_INV_S_3 U889 ( .A(n385), .X(n386) );
  SEN_ND2_3 U890 ( .A1(n1022), .A2(n374), .X(n375) );
  SEN_MUXI2_S_2 U891 ( .D0(n810), .D1(n738), .S(B[3]), .X(n737) );
  SEN_INV_8 U892 ( .A(n743), .X(n518) );
  SEN_ND2_T_2 U893 ( .A1(n328), .A2(n572), .X(n763) );
  SEN_ND2_S_4 U894 ( .A1(n460), .A2(n871), .X(n461) );
  SEN_EO2_S_3 U895 ( .A1(n835), .A2(n834), .X(n1293) );
  SEN_ND2_4 U896 ( .A1(n558), .A2(n557), .X(n765) );
  SEN_AOI31_0P5 U897 ( .A1(n1034), .A2(n823), .A3(n992), .B(n822), .X(n824) );
  SEN_ND2_G_4 U898 ( .A1(n622), .A2(n621), .X(n623) );
  SEN_ND2_S_1P5 U899 ( .A1(B[15]), .A2(n483), .X(n622) );
  SEN_ND3B_V1DG_2 U900 ( .A(n999), .B1(n1002), .B2(n1041), .X(n807) );
  SEN_OR3B_8 U901 ( .B1(n975), .B2(n954), .A(n937), .X(n927) );
  SEN_ND2_T_6 U902 ( .A1(n907), .A2(n723), .X(n871) );
  SEN_ND2B_4 U903 ( .A(n722), .B(n720), .X(n907) );
  SEN_ND2_3 U904 ( .A1(n722), .A2(n721), .X(n723) );
  SEN_NR2_T_4 U905 ( .A1(n395), .A2(n396), .X(n482) );
  SEN_EN2_S_2 U906 ( .A1(n330), .A2(A[19]), .X(n497) );
  SEN_ND2_T_1 U907 ( .A1(n853), .A2(n679), .X(n975) );
  SEN_OAI211_4 U908 ( .A1(n737), .A2(n739), .B1(n518), .B2(n328), .X(n879) );
  SEN_ND2_2 U909 ( .A1(n645), .A2(n327), .X(n674) );
  SEN_AN4B_4 U910 ( .B1(n754), .B2(n901), .B3(n900), .A(n491), .X(n342) );
  SEN_ND2_4 U911 ( .A1(n901), .A2(n427), .X(n908) );
  SEN_ND2_S_4 U912 ( .A1(n463), .A2(n464), .X(n466) );
  SEN_AN4B_4 U913 ( .B1(n754), .B2(n901), .B3(n900), .A(n491), .X(n751) );
  SEN_ND2_S_0P5 U914 ( .A1(n901), .A2(n900), .X(n902) );
  SEN_MUXI2_DG_2 U915 ( .D0(n797), .D1(n404), .S(B[17]), .X(n610) );
  SEN_EO2_4 U916 ( .A1(n330), .A2(A[22]), .X(n773) );
  SEN_AOI21B_2 U917 ( .A1(n842), .A2(n841), .B(n1030), .X(n843) );
  SEN_OAI211_2 U918 ( .A1(n433), .A2(n962), .B1(n980), .B2(n857), .X(n858) );
  SEN_OA21_2 U919 ( .A1(n433), .A2(n962), .B(n980), .X(n407) );
  SEN_INV_2P5 U920 ( .A(n980), .X(n396) );
  SEN_AOAI211_6 U921 ( .A1(n1032), .A2(n821), .B(n785), .C(n784), .X(n790) );
  SEN_NR2_T_2 U922 ( .A1(n773), .A2(n774), .X(n775) );
  SEN_AOAI211_6 U923 ( .A1(n878), .A2(n879), .B(n876), .C(n880), .X(n899) );
  SEN_INV_32 U924 ( .A(A[20]), .X(n345) );
  SEN_ND2_T_1P5 U925 ( .A1(n611), .A2(n610), .X(n613) );
  SEN_INV_0P8 U926 ( .A(n613), .X(n614) );
  SEN_INV_S_2 U927 ( .A(n592), .X(n587) );
  SEN_AN2_S_1 U928 ( .A1(n817), .A2(n494), .X(n347) );
  SEN_OR2_1 U929 ( .A1(n805), .A2(n349), .X(n348) );
  SEN_INV_S_1 U930 ( .A(n817), .X(n349) );
  SEN_ND2_T_2 U931 ( .A1(n943), .A2(n944), .X(n454) );
  SEN_OAI21B_4 U932 ( .A1(n682), .A2(n332), .B(n680), .X(n851) );
  SEN_ND2_3 U933 ( .A1(n683), .A2(n942), .X(n845) );
  SEN_AN3B_2 U934 ( .B1(n939), .B2(n938), .A(n928), .X(n929) );
  SEN_ND2_T_4 U935 ( .A1(n839), .A2(n768), .X(n1022) );
  SEN_MUXI2_S_0P5 U936 ( .D0(n1273), .D1(n1272), .S(INST[3]), .X(Z[13]) );
  SEN_ND2_2 U937 ( .A1(n1025), .A2(n1017), .X(n1038) );
  SEN_ND2_2 U938 ( .A1(n327), .A2(n582), .X(n597) );
  SEN_ND2_G_3 U939 ( .A1(n571), .A2(n570), .X(n780) );
  SEN_MUXI2_DG_2 U940 ( .D0(n522), .D1(n520), .S(B[26]), .X(n570) );
  SEN_MUXI2_S_0P5 U941 ( .D0(n487), .D1(n1260), .S(INST[3]), .X(Z[7]) );
  SEN_ND2_3 U942 ( .A1(n717), .A2(n327), .X(n722) );
  SEN_NR2_3 U943 ( .A1(n914), .A2(n854), .X(n469) );
  SEN_ND2B_2 U944 ( .A(n469), .B(n916), .X(n955) );
  SEN_AO32_4 U945 ( .A1(n638), .A2(n639), .A3(n328), .B1(n637), .B2(n636), .X(
        n680) );
  SEN_OR2_5 U946 ( .A1(n1022), .A2(n1043), .X(n820) );
  SEN_EO2_S_3 U947 ( .A1(n1005), .A2(n1004), .X(n1315) );
  SEN_EN2_1 U948 ( .A1(A[28]), .A2(n524), .X(n566) );
  SEN_OR2_2 U949 ( .A1(n956), .A2(n917), .X(n350) );
  SEN_ND2_S_4 U950 ( .A1(n847), .A2(n616), .X(n946) );
  SEN_ND2_T_1 U951 ( .A1(n1037), .A2(n516), .X(n371) );
  SEN_EO2_3 U952 ( .A1(n352), .A2(n860), .X(n1268) );
  SEN_NR2B_V1_4 U953 ( .A(n328), .B(n735), .X(n517) );
  SEN_EN2_8 U954 ( .A1(n402), .A2(A[3]), .X(n743) );
  SEN_EO2_G_4 U955 ( .A1(n942), .A2(n929), .X(n1282) );
  SEN_ND2_2 U956 ( .A1(n528), .A2(n686), .X(n749) );
  SEN_ND2_0P5 U957 ( .A1(B[12]), .A2(n483), .X(n619) );
  SEN_BUF_1 U958 ( .A(n967), .X(n352) );
  SEN_EN2_1 U959 ( .A1(A[24]), .A2(n329), .X(n548) );
  SEN_ND2_2 U960 ( .A1(n628), .A2(n627), .X(n633) );
  SEN_INV_S_2 U961 ( .A(n761), .X(n762) );
  SEN_AOI21B_2 U962 ( .A1(n1041), .A2(n825), .B(n824), .X(n826) );
  SEN_MUXI2_S_0P5 U963 ( .D0(n519), .D1(n1262), .S(INST[3]), .X(Z[8]) );
  SEN_OR3B_2 U964 ( .B1(n556), .B2(n555), .A(n554), .X(n511) );
  SEN_INV_2 U965 ( .A(n850), .X(n829) );
  SEN_ND2_3 U966 ( .A1(n354), .A2(n355), .X(n356) );
  SEN_ND2_2 U967 ( .A1(n796), .A2(B[15]), .X(n355) );
  SEN_INV_S_0P5 U968 ( .A(n863), .X(n898) );
  SEN_MUXI2_DG_5 U969 ( .D0(n522), .D1(n404), .S(B[24]), .X(n557) );
  SEN_INV_S_0P5 U970 ( .A(n851), .X(n953) );
  SEN_INV_2 U971 ( .A(n1021), .X(n374) );
  SEN_NR3_T_6 U972 ( .A1(n1046), .A2(n1045), .A3(n1044), .X(n1047) );
  SEN_ND2_2 U973 ( .A1(B[0]), .A2(n483), .X(n697) );
  SEN_ND3B_V1DG_4 U974 ( .A(n1243), .B1(n1247), .B2(n1250), .X(n896) );
  SEN_AOI21B_2 U975 ( .A1(n886), .A2(n885), .B(n879), .X(n873) );
  SEN_OR3B_12 U976 ( .B1(n555), .B2(n556), .A(n554), .X(n738) );
  SEN_ND2_T_1 U977 ( .A1(n738), .A2(B[6]), .X(n367) );
  SEN_MUXI2_S_3 U978 ( .D0(n810), .D1(n511), .S(B[22]), .X(n776) );
  SEN_MUXI2_DG_1 U979 ( .D0(n810), .D1(n511), .S(B[3]), .X(n740) );
  SEN_AOI21B_3 U980 ( .A1(n1041), .A2(n1040), .B(n331), .X(n1042) );
  SEN_ND3_T_4 U981 ( .A1(n1006), .A2(n1311), .A3(n1315), .X(n1046) );
  SEN_NR3_0P5 U982 ( .A1(n935), .A2(n975), .A3(n954), .X(n944) );
  SEN_INV_S_1 U983 ( .A(n975), .X(n988) );
  SEN_ND2_G_1 U984 ( .A1(n665), .A2(n664), .X(n512) );
  SEN_ND2_4 U985 ( .A1(n375), .A2(n376), .X(n1300) );
  SEN_AO21B_4 U986 ( .A1(n1041), .A2(n1036), .B(n1035), .X(n516) );
  SEN_INV_S_2 U987 ( .A(n844), .X(n1032) );
  SEN_OAI21_S_2 U988 ( .A1(n840), .A2(n1022), .B(n839), .X(n1030) );
  SEN_INV_5 U989 ( .A(N68), .X(n553) );
  SEN_INV_2 U990 ( .A(n676), .X(n677) );
  SEN_INV_0P8 U991 ( .A(n715), .X(n712) );
  SEN_INV_4 U992 ( .A(n812), .X(n526) );
  SEN_ND2_2 U993 ( .A1(B[5]), .A2(n525), .X(n736) );
  SEN_INV_4 U994 ( .A(n526), .X(n525) );
  SEN_NR2_T_16 U995 ( .A1(n474), .A2(B[31]), .X(n545) );
  SEN_INV_32 U996 ( .A(INST[1]), .X(n474) );
  SEN_EN2_S_1 U997 ( .A1(A[27]), .A2(n524), .X(n563) );
  SEN_ND2_2 U998 ( .A1(n413), .A2(n899), .X(n869) );
  SEN_AOI311_4 U999 ( .A1(n450), .A2(n922), .A3(n479), .B1(n921), .B2(n920), 
        .X(n924) );
  SEN_ND2_2 U1000 ( .A1(n654), .A2(n653), .X(n655) );
  SEN_AOI21B_3 U1001 ( .A1(n1041), .A2(n1020), .B(n1019), .X(n1021) );
  SEN_NR2_T_1 U1002 ( .A1(n1038), .A2(n1018), .X(n1020) );
  SEN_AO21_4 U1003 ( .A1(n492), .A2(n341), .B(n671), .X(n486) );
  SEN_ND3B_V1DG_4 U1004 ( .A(n733), .B1(n732), .B2(n736), .X(n752) );
  SEN_ND2_3 U1005 ( .A1(B[2]), .A2(n483), .X(n744) );
  SEN_INV_3 U1006 ( .A(n744), .X(n739) );
  SEN_ND2_2 U1007 ( .A1(n866), .A2(n412), .X(n707) );
  SEN_AN4B_1 U1008 ( .B1(n831), .B2(n915), .B3(n919), .A(n955), .X(n833) );
  SEN_INV_S_1 U1009 ( .A(n672), .X(n673) );
  SEN_ND2_T_2 U1010 ( .A1(n796), .A2(B[19]), .X(n389) );
  SEN_OAI221_4 U1011 ( .A1(n746), .A2(n745), .B1(n743), .B2(n744), .C(n742), 
        .X(n878) );
  SEN_ND4B_2 U1012 ( .A(n1008), .B1(n1013), .B2(n992), .B3(n1034), .X(n600) );
  SEN_AN4B_1 U1013 ( .B1(n980), .B2(n979), .B3(n964), .A(n963), .X(n965) );
  SEN_MUXI2_S_3 U1014 ( .D0(n810), .D1(n738), .S(B[14]), .X(n638) );
  SEN_AN3_2 U1015 ( .A1(n454), .A2(n455), .A3(n940), .X(n945) );
  SEN_ND2B_16 U1016 ( .A(N68), .B(INST[2]), .X(n551) );
  SEN_OAI21B_1 U1017 ( .A1(n433), .A2(n962), .B(n977), .X(n986) );
  SEN_MUXI2_S_0P5 U1018 ( .D0(n489), .D1(n1267), .S(INST[3]), .X(Z[10]) );
  SEN_INV_1 U1019 ( .A(n883), .X(n358) );
  SEN_EO2_2 U1020 ( .A1(n827), .A2(n826), .X(n1309) );
  SEN_ND4B_8 U1021 ( .A(n1286), .B1(n930), .B2(n1291), .B3(n1282), .X(n948) );
  SEN_ND2_S_3 U1022 ( .A1(n447), .A2(n448), .X(n449) );
  SEN_AO21B_6 U1023 ( .A1(n908), .A2(n907), .B(n754), .X(n980) );
  SEN_ND2_S_3 U1024 ( .A1(n688), .A2(n687), .X(n747) );
  SEN_ND2_G_0P65 U1025 ( .A1(n797), .A2(n353), .X(n354) );
  SEN_INV_S_1 U1026 ( .A(B[15]), .X(n353) );
  SEN_INV_S_3 U1027 ( .A(n356), .X(n627) );
  SEN_ND2_T_0P5 U1028 ( .A1(n797), .A2(n361), .X(n362) );
  SEN_ND2_2 U1029 ( .A1(n362), .A2(n363), .X(n364) );
  SEN_INV_S_1 U1030 ( .A(B[8]), .X(n361) );
  SEN_ND2_T_2 U1031 ( .A1(n710), .A2(n709), .X(n715) );
  SEN_ND2_G_0P65 U1032 ( .A1(n810), .A2(n365), .X(n366) );
  SEN_ND2_2 U1033 ( .A1(n366), .A2(n367), .X(n368) );
  SEN_INV_1 U1034 ( .A(B[6]), .X(n365) );
  SEN_ND2_G_1 U1035 ( .A1(n517), .A2(n733), .X(n734) );
  SEN_INV_S_1 U1036 ( .A(n1037), .X(n369) );
  SEN_INV_S_3 U1037 ( .A(n516), .X(n370) );
  SEN_ND2_S_3 U1038 ( .A1(n373), .A2(n1021), .X(n376) );
  SEN_INV_S_0P5 U1039 ( .A(n1022), .X(n373) );
  SEN_AN2_S_0P5 U1040 ( .A1(n1002), .A2(n1013), .X(n377) );
  SEN_ND2_S_0P5 U1041 ( .A1(n810), .A2(n378), .X(n379) );
  SEN_INV_S_1 U1042 ( .A(B[9]), .X(n378) );
  SEN_INV_S_0P5 U1043 ( .A(n996), .X(n381) );
  SEN_AOI21B_2 U1044 ( .A1(n1041), .A2(n994), .B(n993), .X(n995) );
  SEN_MUXI2_S_1 U1045 ( .D0(n1311), .D1(n1310), .S(INST[3]), .X(Z[28]) );
  SEN_NR4_6 U1046 ( .A1(n1255), .A2(n896), .A3(n1251), .A4(n1253), .X(n911) );
  SEN_ND2_G_1 U1047 ( .A1(n797), .A2(n387), .X(n388) );
  SEN_INV_1 U1048 ( .A(B[19]), .X(n387) );
  SEN_ND2_G_1 U1049 ( .A1(n797), .A2(n391), .X(n392) );
  SEN_INV_S_1 U1050 ( .A(B[0]), .X(n391) );
  SEN_EO2_2 U1051 ( .A1(n973), .A2(n972), .X(n862) );
  SEN_OAOI211_4 U1052 ( .A1(n1003), .A2(n1016), .B(n1002), .C(n1001), .X(n1004) );
  SEN_AN4B_1 U1053 ( .B1(n1024), .B2(n819), .B3(n992), .A(n932), .X(n825) );
  SEN_ND2B_V1_3 U1054 ( .A(n782), .B(n780), .X(n992) );
  SEN_EN2_S_2 U1055 ( .A1(A[0]), .A2(n330), .X(n692) );
  SEN_INV_2 U1056 ( .A(n615), .X(n612) );
  SEN_ND2_2 U1057 ( .A1(n615), .A2(n614), .X(n616) );
  SEN_OR3B_2 U1058 ( .B1(n773), .B2(n478), .A(n778), .X(n1025) );
  SEN_MUXI2_S_1 U1059 ( .D0(n1303), .D1(n1302), .S(INST[3]), .X(Z[25]) );
  SEN_MUXI2_S_1 U1060 ( .D0(n1306), .D1(n1305), .S(INST[3]), .X(Z[26]) );
  SEN_ND2_G_1 U1061 ( .A1(n729), .A2(n728), .X(n730) );
  SEN_AN4B_1 U1062 ( .B1(n997), .B2(n1023), .B3(n1026), .A(n1000), .X(n842) );
  SEN_MUXI2_S_1 U1063 ( .D0(n1297), .D1(n1296), .S(INST[3]), .X(Z[23]) );
  SEN_INV_0P8 U1064 ( .A(n871), .X(n459) );
  SEN_INV_S_0P5 U1065 ( .A(n1225), .X(n405) );
  SEN_INV_1 U1066 ( .A(n1225), .X(n1203) );
  SEN_INV_0P5 U1067 ( .A(n1227), .X(n406) );
  SEN_OR2_2 U1068 ( .A1(n875), .A2(n867), .X(n413) );
  SEN_INV_1 U1069 ( .A(B[10]), .X(n414) );
  SEN_INV_1 U1070 ( .A(A[14]), .X(n421) );
  SEN_INV_S_3 U1071 ( .A(n426), .X(n427) );
  SEN_ND2_0P5 U1072 ( .A1(A[7]), .A2(n330), .X(n431) );
  SEN_INV_S_1 U1073 ( .A(A[7]), .X(n430) );
  SEN_INV_S_0P5 U1074 ( .A(n953), .X(n434) );
  SEN_INV_S_0P5 U1075 ( .A(n950), .X(n438) );
  SEN_INV_S_0P5 U1076 ( .A(n954), .X(n442) );
  SEN_INV_S_2 U1077 ( .A(n485), .X(n443) );
  SEN_INV_1 U1078 ( .A(n1277), .X(n1279) );
  SEN_INV_S_0P5 U1079 ( .A(n958), .X(n479) );
  SEN_ND2_S_0P5 U1080 ( .A1(n706), .A2(n705), .X(n889) );
  SEN_ND2_S_0P65 U1081 ( .A1(n1203), .A2(n1202), .X(n1204) );
  SEN_ND2_S_1 U1082 ( .A1(n1203), .A2(n1080), .X(n1081) );
  SEN_INV_S_1 U1083 ( .A(B[16]), .X(n446) );
  SEN_INV_S_32 U1084 ( .A(INST[2]), .X(n550) );
  SEN_ND2B_1 U1085 ( .A(n816), .B(n815), .X(n817) );
  SEN_EO2_S_0P5 U1086 ( .A1(n816), .A2(n815), .X(n494) );
  SEN_INV_1 U1087 ( .A(A[6]), .X(n451) );
  SEN_INV_S_0P5 U1088 ( .A(n804), .X(n805) );
  SEN_ND2_S_0P5 U1089 ( .A1(n942), .A2(n941), .X(n455) );
  SEN_INV_1 U1090 ( .A(A[9]), .X(n475) );
  SEN_INV_1 U1091 ( .A(n1038), .X(n1040) );
  SEN_MUXI2_S_0P5 U1092 ( .D0(n1285), .D1(n1284), .S(INST[3]), .X(Z[17]) );
  SEN_ND2_S_0P5 U1093 ( .A1(n1203), .A2(n1156), .X(n1157) );
  SEN_INV_S_0P5 U1094 ( .A(n946), .X(n463) );
  SEN_ND2_S_1 U1095 ( .A1(n991), .A2(n789), .X(n827) );
  SEN_NR2_S_1 U1096 ( .A1(n1261), .A2(n1263), .X(n1115) );
  SEN_NR2_S_1 U1097 ( .A1(n1266), .A2(n1269), .X(n1116) );
  SEN_INV_S_2 U1098 ( .A(n580), .X(n578) );
  SEN_NR3_1 U1099 ( .A1(n1184), .A2(n1183), .A3(n1182), .X(n1238) );
  SEN_ND2_S_1 U1100 ( .A1(n1161), .A2(n1160), .X(n1184) );
  SEN_NR3_1 U1101 ( .A1(n1236), .A2(n1235), .A3(n1234), .X(n1237) );
  SEN_ND2_S_1 U1102 ( .A1(n1209), .A2(n1208), .X(n1236) );
  SEN_ND2_S_1 U1103 ( .A1(n1159), .A2(n1158), .X(n1301) );
  SEN_ND2_S_1 U1104 ( .A1(n1207), .A2(n1206), .X(n1283) );
  SEN_ND2_S_1 U1105 ( .A1(n1144), .A2(n1143), .X(n1304) );
  SEN_ND2_S_1 U1106 ( .A1(n1154), .A2(n1153), .X(n1298) );
  SEN_ND2_S_1 U1107 ( .A1(n1189), .A2(n1188), .X(n1287) );
  SEN_ND2_S_1 U1108 ( .A1(n1149), .A2(n1148), .X(n1307) );
  SEN_NR2_1 U1109 ( .A1(n1027), .A2(n818), .X(n819) );
  SEN_ND4B_1 U1110 ( .A(n1240), .B1(n1239), .B2(n1238), .B3(n1237), .X(n1241)
         );
  SEN_NR3_G_1 U1111 ( .A1(n1139), .A2(n1138), .A3(n1137), .X(n1239) );
  SEN_INV_S_0P5 U1112 ( .A(n861), .X(n973) );
  SEN_NR2_1 U1113 ( .A1(n1257), .A2(n1259), .X(n1094) );
  SEN_NR2_1 U1114 ( .A1(n1254), .A2(n1256), .X(n1093) );
  SEN_NR2_1 U1115 ( .A1(n1248), .A2(n1252), .X(n1092) );
  SEN_INV_S_0P5 U1116 ( .A(n800), .X(n801) );
  SEN_INV_1 U1117 ( .A(n786), .X(n787) );
  SEN_NR2_1 U1118 ( .A1(n1280), .A2(n1283), .X(n1208) );
  SEN_NR2_1 U1119 ( .A1(n1298), .A2(n1301), .X(n1160) );
  SEN_NR2_1 U1120 ( .A1(n1304), .A2(n1307), .X(n1161) );
  SEN_NR2_1 U1121 ( .A1(n1287), .A2(n1289), .X(n1209) );
  SEN_ND2_S_0P5 U1122 ( .A1(n1203), .A2(n1191), .X(n1192) );
  SEN_ND2_S_0P5 U1123 ( .A1(n1203), .A2(n1151), .X(n1152) );
  SEN_ND2_S_0P5 U1124 ( .A1(n1203), .A2(n1141), .X(n1142) );
  SEN_ND2_S_0P5 U1125 ( .A1(n1203), .A2(n1111), .X(n1112) );
  SEN_INV_1 U1126 ( .A(n1027), .X(n1011) );
  SEN_INV_0P8 U1127 ( .A(n478), .X(n528) );
  SEN_INV_S_0P5 U1128 ( .A(n478), .X(n529) );
  SEN_NR2_S_0P5 U1129 ( .A1(n960), .A2(n959), .X(n968) );
  SEN_INV_S_0P5 U1130 ( .A(n982), .X(n983) );
  SEN_INV_S_0P5 U1131 ( .A(n916), .X(n917) );
  SEN_ND2_S_0P5 U1132 ( .A1(n1034), .A2(n839), .X(n1027) );
  SEN_INV_S_0P5 U1133 ( .A(n1025), .X(n818) );
  SEN_ND3_S_0P5 U1134 ( .A1(n1026), .A2(n1025), .A3(n1024), .X(n1028) );
  SEN_NR2_S_0P5 U1135 ( .A1(n492), .A2(n974), .X(n960) );
  SEN_NR2B_V1DG_1 U1136 ( .A(n1037), .B(n1007), .X(n822) );
  SEN_INV_S_0P5 U1137 ( .A(n1034), .X(n1031) );
  SEN_INV_S_0P5 U1138 ( .A(n540), .X(n538) );
  SEN_ND2_S_1 U1139 ( .A1(n804), .A2(n803), .X(n1005) );
  SEN_MUXI2_S_0P5 U1140 ( .D0(n1293), .D1(n1292), .S(INST[3]), .X(Z[21]) );
  SEN_ND4_S_1 U1141 ( .A1(n1094), .A2(n1093), .A3(n1092), .A4(n1091), .X(n1240) );
  SEN_ND2_S_1 U1142 ( .A1(n782), .A2(n781), .X(n783) );
  SEN_MUXI2_S_0P5 U1143 ( .D0(n1247), .D1(n1246), .S(INST[3]), .X(Z[1]) );
  SEN_INV_S_0P5 U1144 ( .A(n1245), .X(n1246) );
  SEN_INV_S_0P5 U1145 ( .A(n540), .X(n539) );
  SEN_ND2B_S_0P5 U1146 ( .A(n802), .B(n800), .X(n804) );
  SEN_INV_S_0P5 U1147 ( .A(n757), .X(n758) );
  SEN_ND2_S_1 U1148 ( .A1(n1116), .A2(n1115), .X(n1139) );
  SEN_MUX2_DG_1 U1149 ( .D0(n1288), .D1(n1289), .S(INST[3]), .X(Z[19]) );
  SEN_ND2_S_0P5 U1150 ( .A1(B[30]), .A2(n525), .X(n813) );
  SEN_ND2_S_0P5 U1151 ( .A1(n809), .A2(n529), .X(n816) );
  SEN_NR2_S_1 U1152 ( .A1(n1233), .A2(n1232), .X(n1294) );
  SEN_MUXI2_D_1 U1153 ( .D0(n1227), .D1(n1226), .S(A[22]), .X(n1233) );
  SEN_NR2_S_0P5 U1154 ( .A1(n1229), .A2(n539), .X(n1230) );
  SEN_NR2_S_1 U1155 ( .A1(n1131), .A2(n1130), .X(n1278) );
  SEN_NR2_S_0P5 U1156 ( .A1(n1128), .A2(n539), .X(n1129) );
  SEN_NR2_S_0P5 U1157 ( .A1(n1211), .A2(n539), .X(n1212) );
  SEN_NR2_S_0P5 U1158 ( .A1(n1123), .A2(n539), .X(n1124) );
  SEN_NR2_S_0P5 U1159 ( .A1(n1216), .A2(n539), .X(n1217) );
  SEN_NR2_S_1 U1160 ( .A1(n1171), .A2(n1170), .X(n1310) );
  SEN_NR2_S_0P5 U1161 ( .A1(n1168), .A2(n539), .X(n1169) );
  SEN_NR2_S_1 U1162 ( .A1(n1181), .A2(n1180), .X(n1314) );
  SEN_MUXI2_D_1 U1163 ( .D0(n1227), .D1(n1177), .S(A[30]), .X(n1181) );
  SEN_NR2_S_0P5 U1164 ( .A1(n1178), .A2(n539), .X(n1179) );
  SEN_ND2_G_1 U1165 ( .A1(B[18]), .A2(n812), .X(n586) );
  SEN_NR2_S_0P5 U1166 ( .A1(n1118), .A2(n539), .X(n1119) );
  SEN_NR2_S_0P5 U1167 ( .A1(n1221), .A2(n539), .X(n1222) );
  SEN_NR2_S_0P5 U1168 ( .A1(n1163), .A2(n539), .X(n1164) );
  SEN_NR2_S_1 U1169 ( .A1(n1176), .A2(n1175), .X(n1316) );
  SEN_NR2_S_0P5 U1170 ( .A1(n1173), .A2(n218), .X(n1174) );
  SEN_ND2_S_0P5 U1171 ( .A1(n1203), .A2(n1101), .X(n1102) );
  SEN_ND2_S_0P5 U1172 ( .A1(n1203), .A2(n1096), .X(n1097) );
  SEN_ND2_S_0P5 U1173 ( .A1(n1203), .A2(n1106), .X(n1107) );
  SEN_ND2_S_0P5 U1174 ( .A1(n1203), .A2(n1146), .X(n1147) );
  SEN_ND2_S_0P5 U1175 ( .A1(n1203), .A2(n1076), .X(n1077) );
  SEN_ND2_S_0P5 U1176 ( .A1(n405), .A2(n1071), .X(n1072) );
  SEN_ND2_S_0P5 U1177 ( .A1(n405), .A2(n1061), .X(n1062) );
  SEN_ND2_S_0P5 U1178 ( .A1(n405), .A2(n1056), .X(n1057) );
  SEN_ND2_S_0P5 U1179 ( .A1(n405), .A2(n1066), .X(n1067) );
  SEN_ND2_S_0P5 U1180 ( .A1(n405), .A2(n1051), .X(n1052) );
  SEN_ND2_S_0P5 U1181 ( .A1(n1203), .A2(n1186), .X(n1187) );
  SEN_ND2_S_0P5 U1182 ( .A1(n405), .A2(n1087), .X(n1088) );
  SEN_ND2_S_0P5 U1183 ( .A1(n1203), .A2(n1196), .X(n1197) );
  SEN_ND2_S_0P5 U1184 ( .A1(B[24]), .A2(n812), .X(n574) );
  SEN_NR2_S_0P5 U1185 ( .A1(n499), .A2(n1225), .X(n1122) );
  SEN_NR2_S_0P5 U1186 ( .A1(n502), .A2(n1225), .X(n1117) );
  SEN_NR2_S_0P5 U1187 ( .A1(n500), .A2(n1225), .X(n1132) );
  SEN_NR2_S_0P5 U1188 ( .A1(n501), .A2(n1225), .X(n1127) );
  SEN_NR2_S_0P5 U1189 ( .A1(n503), .A2(n1225), .X(n1167) );
  SEN_NR2_S_0P5 U1190 ( .A1(n504), .A2(n1225), .X(n1162) );
  SEN_NR2_S_0P5 U1191 ( .A1(n505), .A2(n1225), .X(n1177) );
  SEN_NR2_S_0P5 U1192 ( .A1(n506), .A2(n1225), .X(n1172) );
  SEN_NR2_S_0P5 U1193 ( .A1(n507), .A2(n1225), .X(n1210) );
  SEN_NR2_S_0P5 U1194 ( .A1(n509), .A2(n1225), .X(n1220) );
  SEN_NR2_S_0P5 U1195 ( .A1(n510), .A2(n1225), .X(n1215) );
  SEN_NR2_S_0P5 U1196 ( .A1(n508), .A2(n1225), .X(n1226) );
  SEN_NR2_G_1 U1197 ( .A1(n740), .A2(n739), .X(n741) );
  SEN_ND2_S_0P5 U1198 ( .A1(B[7]), .A2(n483), .X(n710) );
  SEN_ND2_S_0P5 U1199 ( .A1(B[22]), .A2(n812), .X(n561) );
  SEN_AN4B_1 U1200 ( .B1(n1011), .B2(n1010), .B3(n1013), .A(n1009), .X(n1014)
         );
  SEN_NR2_1 U1201 ( .A1(n1008), .A2(n1007), .X(n1010) );
  SEN_NR3_1 U1202 ( .A1(n1029), .A2(n1028), .A3(n1027), .X(n1036) );
  SEN_NR2_G_1 U1203 ( .A1(n837), .A2(n990), .X(n841) );
  SEN_INV_1 U1204 ( .A(n1019), .X(n840) );
  SEN_INV_2 U1205 ( .A(n991), .X(n1008) );
  SEN_INV_S_1 U1206 ( .A(n533), .X(n531) );
  SEN_INV_S_1 U1207 ( .A(n534), .X(n530) );
  SEN_INV_S_1 U1208 ( .A(n1231), .X(n1201) );
  SEN_INV_S_1 U1209 ( .A(n1227), .X(n1205) );
  SEN_INV_S_1 U1210 ( .A(n1231), .X(n1083) );
  SEN_AO21_DG_1 U1211 ( .A1(n351), .A2(n1050), .B(n218), .X(n1225) );
  SEN_INV_S_1 U1212 ( .A(n1248), .X(n1249) );
  SEN_INV_S_1 U1213 ( .A(n1304), .X(n1305) );
  SEN_INV_S_1 U1214 ( .A(n1298), .X(n1299) );
  SEN_INV_S_1 U1215 ( .A(n1259), .X(n1260) );
  SEN_INV_S_1 U1216 ( .A(n1261), .X(n1262) );
  SEN_INV_1 U1217 ( .A(n512), .X(n668) );
  SEN_ND2_G_1 U1218 ( .A1(n788), .A2(n787), .X(n789) );
  SEN_MUX2_DG_1 U1219 ( .D0(n1243), .D1(n1244), .S(INST[3]), .X(Z[0]) );
  SEN_MUX2_DG_1 U1220 ( .D0(n1251), .D1(n1252), .S(INST[3]), .X(Z[3]) );
  SEN_INV_S_1 U1221 ( .A(n1301), .X(n1302) );
  SEN_MUXI2_S_0P5 U1222 ( .D0(n1309), .D1(n1308), .S(INST[3]), .X(Z[27]) );
  SEN_INV_S_1 U1223 ( .A(n1307), .X(n1308) );
  SEN_MUXI2_S_0P5 U1224 ( .D0(n484), .D1(n1258), .S(INST[3]), .X(Z[6]) );
  SEN_INV_S_1 U1225 ( .A(n1257), .X(n1258) );
  SEN_MUXI2_S_0P5 U1226 ( .D0(n1265), .D1(n1264), .S(INST[3]), .X(Z[9]) );
  SEN_INV_S_1 U1227 ( .A(n1263), .X(n1264) );
  SEN_INV_S_1 U1228 ( .A(n1266), .X(n1267) );
  SEN_MUXI2_S_1 U1229 ( .D0(n1276), .D1(n1275), .S(INST[3]), .X(Z[14]) );
  SEN_INV_S_1 U1230 ( .A(n1280), .X(n1281) );
  SEN_INV_S_1 U1231 ( .A(n1283), .X(n1284) );
  SEN_MUX2_DG_1 U1232 ( .D0(n1253), .D1(n1254), .S(INST[3]), .X(Z[4]) );
  SEN_MUXI2_S_1 U1233 ( .D0(n1279), .D1(n1278), .S(INST[3]), .X(Z[15]) );
  SEN_INV_S_1 U1234 ( .A(n495), .X(n541) );
  SEN_INV_S_1 U1235 ( .A(n495), .X(n542) );
  SEN_ND2_G_1 U1236 ( .A1(n759), .A2(n758), .X(n760) );
  SEN_ND2_G_1 U1237 ( .A1(n802), .A2(n801), .X(n803) );
  SEN_INV_1 U1238 ( .A(n776), .X(n562) );
  SEN_ND2_G_1 U1239 ( .A1(n1292), .A2(n1290), .X(n1235) );
  SEN_ND2_G_1 U1240 ( .A1(n1296), .A2(n1294), .X(n1234) );
  SEN_ND2_G_1 U1241 ( .A1(n1316), .A2(n1314), .X(n1182) );
  SEN_ND2_G_1 U1242 ( .A1(n1312), .A2(n1310), .X(n1183) );
  SEN_BUF_S_1 U1243 ( .A(n537), .X(n533) );
  SEN_BUF_S_1 U1244 ( .A(n537), .X(n532) );
  SEN_BUF_S_1 U1245 ( .A(n537), .X(n534) );
  SEN_ND2_G_1 U1246 ( .A1(n1278), .A2(n1275), .X(n1137) );
  SEN_ND2_G_1 U1247 ( .A1(n1272), .A2(n1270), .X(n1138) );
  SEN_INV_S_1 U1248 ( .A(n495), .X(n543) );
  SEN_BUF_S_1 U1249 ( .A(n537), .X(n536) );
  SEN_BUF_S_1 U1250 ( .A(n537), .X(n535) );
  SEN_ND3B_1 U1251 ( .A(INST[2]), .B1(INST[1]), .B2(N68), .X(n1231) );
  SEN_ND3B_1 U1252 ( .A(INST[1]), .B1(N68), .B2(INST[2]), .X(n1227) );
  SEN_EN2_0P5 U1253 ( .A1(n811), .A2(n810), .X(n814) );
  SEN_INV_S_1 U1254 ( .A(n1228), .X(n537) );
  SEN_OR2_1 U1255 ( .A1(INST[1]), .A2(INST[2]), .X(n495) );
  SEN_NR3B_1 U1256 ( .A(N68), .B1(INST[1]), .B2(INST[2]), .X(n218) );
  SEN_ND2_G_1 U1257 ( .A1(n527), .A2(n566), .X(n759) );
  SEN_EN2_0P5 U1258 ( .A1(A[12]), .A2(n330), .X(n645) );
  SEN_EN2_0P5 U1259 ( .A1(A[31]), .A2(n523), .X(n809) );
  SEN_ND2_G_1 U1260 ( .A1(n799), .A2(n798), .X(n800) );
  SEN_ND2_G_1 U1261 ( .A1(B[29]), .A2(n525), .X(n799) );
  SEN_MUXI2_S_0P5 U1262 ( .D0(n797), .D1(n520), .S(B[30]), .X(n798) );
  SEN_NR2_1 U1263 ( .A1(n1136), .A2(n1135), .X(n1275) );
  SEN_MUXI2_S_1 U1264 ( .D0(n1231), .D1(n1134), .S(B[14]), .X(n1135) );
  SEN_MUXI2_S_1 U1265 ( .D0(n1227), .D1(n1132), .S(A[14]), .X(n1136) );
  SEN_NR2_1 U1266 ( .A1(n1133), .A2(n218), .X(n1134) );
  SEN_NR2_1 U1267 ( .A1(n1126), .A2(n1125), .X(n1270) );
  SEN_MUXI2_S_1 U1268 ( .D0(n1231), .D1(n1124), .S(B[12]), .X(n1125) );
  SEN_MUXI2_S_1 U1269 ( .D0(n1227), .D1(n1122), .S(A[12]), .X(n1126) );
  SEN_MUXI2_S_1 U1270 ( .D0(n1231), .D1(n1230), .S(B[22]), .X(n1232) );
  SEN_MUXI2_S_1 U1271 ( .D0(n1231), .D1(n1169), .S(B[28]), .X(n1170) );
  SEN_MUXI2_S_1 U1272 ( .D0(n1227), .D1(n1167), .S(A[28]), .X(n1171) );
  SEN_NR2_1 U1273 ( .A1(n1121), .A2(n1120), .X(n1272) );
  SEN_MUXI2_S_1 U1274 ( .D0(n1231), .D1(n1119), .S(B[13]), .X(n1120) );
  SEN_MUXI2_S_1 U1275 ( .D0(n1227), .D1(n1117), .S(A[13]), .X(n1121) );
  SEN_NR2_1 U1276 ( .A1(n1224), .A2(n1223), .X(n1296) );
  SEN_MUXI2_S_1 U1277 ( .D0(n1231), .D1(n1222), .S(B[23]), .X(n1223) );
  SEN_MUXI2_S_1 U1278 ( .D0(n1227), .D1(n1220), .S(A[23]), .X(n1224) );
  SEN_NR2_1 U1279 ( .A1(n1214), .A2(n1213), .X(n1292) );
  SEN_MUXI2_S_1 U1280 ( .D0(n1231), .D1(n1212), .S(B[21]), .X(n1213) );
  SEN_MUXI2_S_1 U1281 ( .D0(n1227), .D1(n1210), .S(A[21]), .X(n1214) );
  SEN_NR2_1 U1282 ( .A1(n1166), .A2(n1165), .X(n1312) );
  SEN_MUXI2_S_1 U1283 ( .D0(n1231), .D1(n1164), .S(B[29]), .X(n1165) );
  SEN_MUXI2_S_1 U1284 ( .D0(n1227), .D1(n1162), .S(A[29]), .X(n1166) );
  SEN_MUXI2_S_1 U1285 ( .D0(n1231), .D1(n1129), .S(B[15]), .X(n1130) );
  SEN_MUXI2_S_1 U1286 ( .D0(n1227), .D1(n1127), .S(A[15]), .X(n1131) );
  SEN_NR2_1 U1287 ( .A1(n1219), .A2(n1218), .X(n1290) );
  SEN_MUXI2_S_1 U1288 ( .D0(n1231), .D1(n1217), .S(B[20]), .X(n1218) );
  SEN_MUXI2_S_1 U1289 ( .D0(n1227), .D1(n1215), .S(A[20]), .X(n1219) );
  SEN_MUXI2_S_1 U1290 ( .D0(n1231), .D1(n1179), .S(B[30]), .X(n1180) );
  SEN_MUXI2_S_1 U1291 ( .D0(n1231), .D1(n1174), .S(B[31]), .X(n1175) );
  SEN_MUXI2_S_1 U1292 ( .D0(n1227), .D1(n1172), .S(A[31]), .X(n1176) );
  SEN_ND2_G_1 U1293 ( .A1(n1114), .A2(n1113), .X(n1263) );
  SEN_MUXI2_S_1 U1294 ( .D0(n1201), .D1(n1110), .S(B[9]), .X(n1114) );
  SEN_MUXI2_S_1 U1295 ( .D0(n1205), .D1(n1112), .S(A[9]), .X(n1113) );
  SEN_OAI21B_1 U1296 ( .A1(n530), .A2(A[9]), .B(n538), .X(n1110) );
  SEN_ND2_G_1 U1297 ( .A1(n1104), .A2(n1103), .X(n1269) );
  SEN_MUXI2_S_1 U1298 ( .D0(n1201), .D1(n1100), .S(B[11]), .X(n1104) );
  SEN_MUXI2_S_1 U1299 ( .D0(n1205), .D1(n1102), .S(A[11]), .X(n1103) );
  SEN_OAI21B_1 U1300 ( .A1(n530), .A2(A[11]), .B(n538), .X(n1100) );
  SEN_ND2_G_1 U1301 ( .A1(n1079), .A2(n1078), .X(n1252) );
  SEN_MUXI2_S_1 U1302 ( .D0(n1083), .D1(n1075), .S(B[3]), .X(n1079) );
  SEN_MUXI2_S_1 U1303 ( .D0(n406), .D1(n1077), .S(A[3]), .X(n1078) );
  SEN_OAI21B_1 U1304 ( .A1(n530), .A2(A[3]), .B(n539), .X(n1075) );
  SEN_ND2_G_1 U1305 ( .A1(n1069), .A2(n1068), .X(n1256) );
  SEN_MUXI2_S_1 U1306 ( .D0(n1083), .D1(n1065), .S(B[5]), .X(n1069) );
  SEN_MUXI2_S_1 U1307 ( .D0(n406), .D1(n1067), .S(A[5]), .X(n1068) );
  SEN_OAI21B_1 U1308 ( .A1(n531), .A2(A[5]), .B(n539), .X(n1065) );
  SEN_ND2_G_1 U1309 ( .A1(n1059), .A2(n1058), .X(n1259) );
  SEN_MUXI2_S_1 U1310 ( .D0(n1083), .D1(n1055), .S(B[7]), .X(n1059) );
  SEN_MUXI2_S_1 U1311 ( .D0(n406), .D1(n1057), .S(A[7]), .X(n1058) );
  SEN_OAI21B_1 U1312 ( .A1(n531), .A2(A[7]), .B(n538), .X(n1055) );
  SEN_MUXI2_S_1 U1313 ( .D0(n1083), .D1(n1200), .S(B[17]), .X(n1207) );
  SEN_MUXI2_S_1 U1314 ( .D0(n1205), .D1(n1204), .S(A[17]), .X(n1206) );
  SEN_OAI21B_1 U1315 ( .A1(n530), .A2(A[17]), .B(n538), .X(n1200) );
  SEN_ND2_G_1 U1316 ( .A1(n1194), .A2(n1193), .X(n1289) );
  SEN_MUXI2_S_1 U1317 ( .D0(n1201), .D1(n1190), .S(B[19]), .X(n1194) );
  SEN_MUXI2_S_1 U1318 ( .D0(n1205), .D1(n1192), .S(A[19]), .X(n1193) );
  SEN_OAI21B_1 U1319 ( .A1(n530), .A2(A[19]), .B(n538), .X(n1190) );
  SEN_MUXI2_S_1 U1320 ( .D0(n1083), .D1(n1155), .S(B[25]), .X(n1159) );
  SEN_MUXI2_S_1 U1321 ( .D0(n1205), .D1(n1157), .S(A[25]), .X(n1158) );
  SEN_OAI21B_1 U1322 ( .A1(n530), .A2(A[25]), .B(n538), .X(n1155) );
  SEN_MUXI2_S_1 U1323 ( .D0(n1201), .D1(n1145), .S(B[27]), .X(n1149) );
  SEN_MUXI2_S_1 U1324 ( .D0(n1205), .D1(n1147), .S(A[27]), .X(n1148) );
  SEN_OAI21B_1 U1325 ( .A1(n530), .A2(A[27]), .B(n538), .X(n1145) );
  SEN_ND2_G_1 U1326 ( .A1(n1090), .A2(n1089), .X(n1245) );
  SEN_MUXI2_S_1 U1327 ( .D0(n1083), .D1(n1086), .S(B[1]), .X(n1090) );
  SEN_OAI21B_1 U1328 ( .A1(n531), .A2(A[1]), .B(n538), .X(n1086) );
  SEN_ND3_S_0P5 U1329 ( .A1(n1085), .A2(n1084), .A3(n529), .X(n1244) );
  SEN_MUXI2_S_1 U1330 ( .D0(n1201), .D1(n1082), .S(B[0]), .X(n1084) );
  SEN_MUXI2_S_1 U1331 ( .D0(n1205), .D1(n1081), .S(A[0]), .X(n1085) );
  SEN_OAI21B_1 U1332 ( .A1(n531), .A2(A[0]), .B(n538), .X(n1082) );
  SEN_ND2_G_1 U1333 ( .A1(n1109), .A2(n1108), .X(n1261) );
  SEN_MUXI2_S_1 U1334 ( .D0(n1083), .D1(n1105), .S(B[8]), .X(n1109) );
  SEN_MUXI2_S_1 U1335 ( .D0(n1205), .D1(n1107), .S(A[8]), .X(n1108) );
  SEN_OAI21B_1 U1336 ( .A1(n530), .A2(A[8]), .B(n538), .X(n1105) );
  SEN_ND2_G_1 U1337 ( .A1(n1099), .A2(n1098), .X(n1266) );
  SEN_MUXI2_S_1 U1338 ( .D0(n1201), .D1(n1095), .S(B[10]), .X(n1099) );
  SEN_MUXI2_S_1 U1339 ( .D0(n406), .D1(n1097), .S(A[10]), .X(n1098) );
  SEN_OAI21B_1 U1340 ( .A1(n530), .A2(A[10]), .B(n538), .X(n1095) );
  SEN_ND2_G_1 U1341 ( .A1(n1074), .A2(n1073), .X(n1248) );
  SEN_MUXI2_S_1 U1342 ( .D0(n1201), .D1(n1070), .S(B[2]), .X(n1074) );
  SEN_MUXI2_S_1 U1343 ( .D0(n406), .D1(n1072), .S(A[2]), .X(n1073) );
  SEN_OAI21B_1 U1344 ( .A1(n531), .A2(A[2]), .B(n539), .X(n1070) );
  SEN_ND2_G_1 U1345 ( .A1(n1064), .A2(n1063), .X(n1254) );
  SEN_MUXI2_S_1 U1346 ( .D0(n1201), .D1(n1060), .S(B[4]), .X(n1064) );
  SEN_MUXI2_S_1 U1347 ( .D0(n406), .D1(n1062), .S(A[4]), .X(n1063) );
  SEN_OAI21B_1 U1348 ( .A1(n531), .A2(A[4]), .B(n539), .X(n1060) );
  SEN_ND2_G_1 U1349 ( .A1(n1054), .A2(n1053), .X(n1257) );
  SEN_MUXI2_S_1 U1350 ( .D0(n1201), .D1(n1049), .S(B[6]), .X(n1054) );
  SEN_MUXI2_S_1 U1351 ( .D0(n406), .D1(n1052), .S(A[6]), .X(n1053) );
  SEN_OAI21B_1 U1352 ( .A1(n530), .A2(A[6]), .B(n538), .X(n1049) );
  SEN_ND2_G_1 U1353 ( .A1(n1199), .A2(n1198), .X(n1280) );
  SEN_MUXI2_S_1 U1354 ( .D0(n1083), .D1(n1195), .S(B[16]), .X(n1199) );
  SEN_MUXI2_S_1 U1355 ( .D0(n1205), .D1(n1197), .S(A[16]), .X(n1198) );
  SEN_OAI21B_1 U1356 ( .A1(n530), .A2(A[16]), .B(n539), .X(n1195) );
  SEN_MUXI2_S_1 U1357 ( .D0(n1083), .D1(n1185), .S(B[18]), .X(n1189) );
  SEN_MUXI2_S_1 U1358 ( .D0(n406), .D1(n1187), .S(A[18]), .X(n1188) );
  SEN_OAI21B_1 U1359 ( .A1(n530), .A2(A[18]), .B(n538), .X(n1185) );
  SEN_MUXI2_S_1 U1360 ( .D0(n1083), .D1(n1150), .S(B[24]), .X(n1154) );
  SEN_MUXI2_S_1 U1361 ( .D0(n406), .D1(n1152), .S(A[24]), .X(n1153) );
  SEN_OAI21B_1 U1362 ( .A1(n530), .A2(A[24]), .B(n538), .X(n1150) );
  SEN_MUXI2_S_1 U1363 ( .D0(n1201), .D1(n1140), .S(B[26]), .X(n1144) );
  SEN_MUXI2_S_1 U1364 ( .D0(n406), .D1(n1142), .S(A[26]), .X(n1143) );
  SEN_OAI21B_1 U1365 ( .A1(n530), .A2(A[26]), .B(n538), .X(n1140) );
  SEN_MUX2_DG_1 U1366 ( .D0(n535), .D1(n541), .S(B[12]), .X(n499) );
  SEN_MUX2_DG_1 U1367 ( .D0(n535), .D1(n542), .S(B[14]), .X(n500) );
  SEN_MUX2_DG_1 U1368 ( .D0(n535), .D1(n542), .S(B[15]), .X(n501) );
  SEN_MUX2_DG_1 U1369 ( .D0(n535), .D1(n541), .S(B[13]), .X(n502) );
  SEN_MUX2_DG_1 U1370 ( .D0(n535), .D1(n542), .S(B[28]), .X(n503) );
  SEN_MUX2_DG_1 U1371 ( .D0(n535), .D1(n542), .S(B[29]), .X(n504) );
  SEN_MUX2_DG_1 U1372 ( .D0(n535), .D1(n542), .S(B[30]), .X(n505) );
  SEN_MUX2_DG_1 U1373 ( .D0(n535), .D1(n542), .S(B[31]), .X(n506) );
  SEN_MUX2_DG_1 U1374 ( .D0(n536), .D1(n543), .S(B[21]), .X(n507) );
  SEN_MUX2_DG_1 U1375 ( .D0(n536), .D1(n543), .S(B[22]), .X(n508) );
  SEN_MUX2_DG_1 U1376 ( .D0(n536), .D1(n543), .S(B[23]), .X(n509) );
  SEN_MUX2_DG_1 U1377 ( .D0(n536), .D1(n543), .S(B[20]), .X(n510) );
  SEN_ND3_S_0P5 U1378 ( .A1(DI[31]), .A2(n1050), .A3(n693), .X(n695) );
  SEN_ND2_G_1 U1379 ( .A1(n529), .A2(n569), .X(n782) );
  SEN_EN2_0P5 U1380 ( .A1(A[26]), .A2(n329), .X(n569) );
  SEN_EN2_0P5 U1381 ( .A1(A[30]), .A2(n524), .X(n795) );
  SEN_ND2_G_1 U1382 ( .A1(n603), .A2(n602), .X(n791) );
  SEN_ND2_S_0P5 U1383 ( .A1(B[28]), .A2(n812), .X(n603) );
  SEN_MUXI2_S_0P5 U1384 ( .D0(n522), .D1(n404), .S(B[29]), .X(n602) );
  SEN_ND2_S_0P5 U1385 ( .A1(B[16]), .A2(n525), .X(n611) );
  SEN_ND2_G_1 U1386 ( .A1(n568), .A2(n567), .X(n757) );
  SEN_ND2_S_0P5 U1387 ( .A1(B[27]), .A2(n812), .X(n568) );
  SEN_MUXI2_S_0P5 U1388 ( .D0(n797), .D1(n520), .S(B[28]), .X(n567) );
  SEN_ND2_S_0P5 U1389 ( .A1(B[26]), .A2(n812), .X(n565) );
  SEN_MUXI2_S_0P5 U1390 ( .D0(n522), .D1(n404), .S(B[27]), .X(n564) );
  SEN_ND2_S_0P5 U1391 ( .A1(B[19]), .A2(n525), .X(n584) );
  SEN_ND2_S_0P5 U1392 ( .A1(B[11]), .A2(n483), .X(n647) );
  SEN_ND2_S_0P5 U1393 ( .A1(B[25]), .A2(n812), .X(n571) );
  SEN_ND2_S_0P5 U1394 ( .A1(B[17]), .A2(n812), .X(n589) );
  SEN_ND2_S_0P5 U1395 ( .A1(B[20]), .A2(n812), .X(n576) );
  SEN_ND2_S_0P5 U1396 ( .A1(B[23]), .A2(n812), .X(n558) );
  SEN_MUXI2_S_1 U1397 ( .D0(n534), .D1(n541), .S(B[9]), .X(n1111) );
  SEN_MUXI2_S_1 U1398 ( .D0(n534), .D1(n541), .S(B[8]), .X(n1106) );
  SEN_MUXI2_S_1 U1399 ( .D0(n534), .D1(n541), .S(B[11]), .X(n1101) );
  SEN_MUXI2_S_1 U1400 ( .D0(n534), .D1(n541), .S(B[10]), .X(n1096) );
  SEN_MUXI2_S_1 U1401 ( .D0(n535), .D1(n542), .S(B[27]), .X(n1146) );
  SEN_MUXI2_S_1 U1402 ( .D0(n533), .D1(n541), .S(B[3]), .X(n1076) );
  SEN_MUXI2_S_1 U1403 ( .D0(n533), .D1(n541), .S(B[2]), .X(n1071) );
  SEN_MUXI2_S_1 U1404 ( .D0(n532), .D1(n541), .S(B[5]), .X(n1066) );
  SEN_MUXI2_S_1 U1405 ( .D0(n532), .D1(n541), .S(B[4]), .X(n1061) );
  SEN_MUXI2_S_1 U1406 ( .D0(n532), .D1(n541), .S(B[7]), .X(n1056) );
  SEN_MUXI2_S_1 U1407 ( .D0(n532), .D1(n541), .S(B[6]), .X(n1051) );
  SEN_MUXI2_S_1 U1408 ( .D0(n536), .D1(n542), .S(B[18]), .X(n1186) );
  SEN_MUXI2_S_1 U1409 ( .D0(n535), .D1(n542), .S(B[26]), .X(n1141) );
  SEN_MUXI2_S_1 U1410 ( .D0(n536), .D1(n542), .S(B[17]), .X(n1202) );
  SEN_MUXI2_S_1 U1411 ( .D0(n536), .D1(n542), .S(B[19]), .X(n1191) );
  SEN_MUXI2_S_1 U1412 ( .D0(n535), .D1(n542), .S(B[25]), .X(n1156) );
  SEN_MUXI2_S_1 U1413 ( .D0(n535), .D1(n542), .S(B[24]), .X(n1151) );
  SEN_MUXI2_S_1 U1414 ( .D0(n533), .D1(n541), .S(B[1]), .X(n1087) );
  SEN_MUXI2_S_1 U1415 ( .D0(n533), .D1(n541), .S(B[0]), .X(n1080) );
  SEN_MUXI2_S_1 U1416 ( .D0(n536), .D1(n542), .S(B[16]), .X(n1196) );
  SEN_NR2_1 U1417 ( .A1(n531), .A2(A[21]), .X(n1211) );
  SEN_NR2_1 U1418 ( .A1(n531), .A2(A[28]), .X(n1168) );
  SEN_NR2_1 U1419 ( .A1(n531), .A2(A[29]), .X(n1163) );
  SEN_NR2_1 U1420 ( .A1(n531), .A2(A[30]), .X(n1178) );
  SEN_NR2_1 U1421 ( .A1(n531), .A2(A[31]), .X(n1173) );
  SEN_NR2_1 U1422 ( .A1(n531), .A2(A[14]), .X(n1133) );
  SEN_NR2_1 U1423 ( .A1(n531), .A2(A[15]), .X(n1128) );
  SEN_NR2_1 U1424 ( .A1(n531), .A2(A[12]), .X(n1123) );
  SEN_NR2_1 U1425 ( .A1(n531), .A2(A[13]), .X(n1118) );
  SEN_NR2_1 U1426 ( .A1(n1228), .A2(A[22]), .X(n1229) );
  SEN_NR2_1 U1427 ( .A1(n530), .A2(A[23]), .X(n1221) );
  SEN_NR2_1 U1428 ( .A1(n1228), .A2(A[20]), .X(n1216) );
  SEN_TIE0_1 U1429 ( .X(\*Logic0* ) );
  SEN_OR3B_1 U1430 ( .B1(N68), .B2(INST[2]), .A(INST[1]), .X(n1228) );
  SEN_ND2_G_1 U1431 ( .A1(INST[1]), .A2(B[31]), .X(n811) );
  SEN_INV_S_1 U1432 ( .A(n880), .X(n881) );
  SEN_MUXI2_S_0P5 U1433 ( .D0(n1250), .D1(n1249), .S(INST[3]), .X(Z[2]) );
  SEN_MUXI2_S_0P5 U1434 ( .D0(n1291), .D1(n1290), .S(INST[3]), .X(Z[20]) );
  SEN_INV_S_0P5 U1435 ( .A(n492), .X(n514) );
  SEN_BUF_1 U1436 ( .A(n832), .X(n515) );
  SEN_MUXI2_S_0P5 U1437 ( .D0(n324), .D1(n1314), .S(INST[3]), .X(Z[30]) );
  SEN_AOAI211_G_0P5 U1438 ( .A1(n544), .A2(n1050), .B(n814), .C(n813), .X(n815) );
  SEN_OR3B_0P5 U1439 ( .B1(n493), .B2(n954), .A(n937), .X(n938) );
  SEN_EN2_5 U1440 ( .A1(A[25]), .A2(n524), .X(n572) );
endmodule

